* Extracted by KLayout with SG13G2 LVS runset on : 07/04/2025 12:09

.SUBCKT Mixer5GHz GND ICC OSCN VCC OSCP IDC IFP RFN LOP LON VDC IFN RFP
M$1 GND ICC \$93896 GND sg13_lv_nmos L=0.13u W=120u AS=23.7p AD=23.7p PS=133.9u
+ PD=133.9u
M$21 GND ICC ICC GND sg13_lv_nmos L=0.13u W=120u AS=23.7p AD=23.7p PS=133.9u
+ PD=133.9u
M$41 \$93896 OSCP OSCN GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p PS=102u
+ PD=102u
M$56 \$93896 OSCN OSCP GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p PS=102u
+ PD=102u
M$71 GND IDC \$478393 GND sg13_lv_nmos L=0.13u W=120u AS=23.7p AD=23.7p
+ PS=133.9u PD=133.9u
M$91 GND IDC IDC GND sg13_lv_nmos L=0.13u W=240u AS=47.4p AD=47.4p PS=267.8u
+ PD=267.8u
M$131 GND IDC \$478394 GND sg13_lv_nmos L=0.13u W=120u AS=23.7p AD=23.7p
+ PS=133.9u PD=133.9u
M$151 \$478393 LON LOP GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p PS=102u
+ PD=102u
M$166 \$478393 LOP LON GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p PS=102u
+ PD=102u
M$181 \$478394 IFP \$486703 GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p
+ PS=102u PD=102u
M$196 \$478394 IFN \$486704 GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p
+ PS=102u PD=102u
M$211 \$486703 LOP RFP GND sg13_lv_nmos L=0.13u W=60u AS=12.3p AD=12.3p
+ PS=70.1u PD=70.1u
M$221 \$486703 LON RFN GND sg13_lv_nmos L=0.13u W=60u AS=12.3p AD=12.3p
+ PS=70.1u PD=70.1u
M$231 \$486704 LON RFP GND sg13_lv_nmos L=0.13u W=60u AS=12.3p AD=12.3p
+ PS=70.1u PD=70.1u
M$241 \$486704 LOP RFN GND sg13_lv_nmos L=0.13u W=60u AS=12.3p AD=12.3p
+ PS=70.1u PD=70.1u
R$251 OSCP VCC rppd w=4.35u l=1.5u ps=0 b=0 m=1
R$252 OSCN VCC rppd w=4.35u l=1.5u ps=0 b=0 m=1
R$253 RFP VDC rppd w=4.5u l=3.2u ps=0 b=0 m=1
R$254 RFN VDC rppd w=4.5u l=3.2u ps=0 b=0 m=1
R$255 LON VDC rppd w=4.4u l=1.5u ps=0 b=0 m=1
R$256 LOP VDC rppd w=4.4u l=1.5u ps=0 b=0 m=1
C$257 VCC OSCN cap_cmim w=19.1u l=10.7u A=204.37p P=59.6u m=1
C$258 VCC OSCP cap_cmim w=19.1u l=10.7u A=204.37p P=59.6u m=1
C$259 VDC LOP cap_cmim w=11.745u l=9.445u A=110.931525p P=42.38u m=1
C$260 VDC LON cap_cmim w=11.745u l=9.445u A=110.931525p P=42.38u m=1
.ENDS Mixer5GHz
