* Extracted by KLayout with SG13G2 LVS runset on : 05/04/2025 02:52

.SUBCKT lna_full_base_lvs
C$1 \$I6 \$8 \$1 rfcmim w=60u l=55u A=3300p P=230u m=1 wfeed=5u
M$2 \$I28 \$I28 \$1 \$1 rfnmos L=0.36u W=10u AS=2.055p AD=2.055p PS=15.11u
+ PD=15.11u
Q$12 \$5 \$2 \$I17 \$1 npn13G2 AE=0.063p PE=1.94u AB=63.456p PB=45.22u
+ AC=63.429884p PC=45.21u NE=60 m=60
Q$22 \$I17 \$8 \$1 \$1 npn13G2 AE=0.063p PE=1.94u AB=63.456p PB=45.22u
+ AC=63.429884p PC=45.21u NE=60 m=60
R$132 \$4 \$I6 rsil w=0.5u l=2.4u ps=0 b=0 m=1
R$133 \$I28 \$2 rppd w=0.5u l=1.8u ps=0 b=0 m=1
R$134 \$8 \$I28 rppd w=0.5u l=3.6u ps=0 b=0 m=1
.ENDS lna_full_base_lvs
