** sch_path: /home/noritsuna/LNA/202504/submit/lvs/parts/vbias_inp_lvs.sch
.subckt vbias_inp_lvs VDD IN VSS VBIAS_OUT
*.PININFO VDD:B IN:I VSS:B VBIAS_OUT:B
R2 VBIAS_OUT net1 rppd w=0.5e-6 l=3.6e-6 m=1 b=0
R1 net1 VDD rppd w=0.5e-6 l=1.8e-6 m=1 b=0
R3 net2 IN rsil w=0.5e-6 l=2.4e-6 m=1 b=0
C1 net2 VBIAS_OUT VSS rfcmim w=60.0e-6 l=55.0e-6 wfeed=5.0e-6
M3 net1 net1 VSS VSS rfnmos l=0.36u w=10.0u ng=5
.ends
.end
