*Modified Qucs-s netlist for KLAYOUT LVS check

.SUBCKT TOP

Rbulk VSS VSS ptap1 A=3.6504p P=18.72u

Rq2 OUTPUT VDD2V1 rppd w=11.5u l=2u ps=0 b=0 m=1

Rq1 VDD2V \connection rppd w=15u l=4u ps=0 b=0 m=1

Rrf INPUT \connection rppd w=30u l=6u ps=0 b=0 m=1

Qq1 \connection INPUT VSS VSS npn13G2 AE=0.063p PE=1.94u AB=31.9135p PB=26.72u
+ AC=31.896634p PC=26.71u NE=5 m=5

Qq2 OUTPUT \connection VSS VSS npn13G2 AE=0.063p PE=1.94u AB=25.605p PB=23.02u
+ AC=25.589984p PC=23.01u NE=4 m=4

C19 VDD2V VSS cap_cmim w=30u l=30u A=900p P=120u m=1

C20 VDD2V1 VSS cap_cmim w=30u l=30u A=900p P=120u m=1
.ENDS TOP
