.SUBCKT TOP GND|TLA|TLB TLA|TLB|VCC2 RFIN|RFIN1|TLA|TLB RFIN2|RFOUT1
+ RFIN3|RFOUT2|TLA|TLB RFOUT|RFOUT3|TLA|TLB TLA|TLB|VCC1|VCC3
+ TLA|TLB|VCC1|VCC31
Q1 RFIN2|RFOUT1 RFIN|RFIN1|TLA|TLB GND|TLA|TLB GND|TLA|TLB npn13G2 AE=0.063p
+ PE=1.94u AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=10 m=10
Q11 RFOUT|RFOUT3|TLA|TLB RFIN3|RFOUT2|TLA|TLB GND|TLA|TLB GND|TLA|TLB npn13G2
+ AE=0.063p PE=1.94u AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=10 m=10
Q21 TLA|TLB|VCC2 RFIN2|RFOUT1 RFIN3|RFOUT2|TLA|TLB GND|TLA|TLB npn13G2
+ AE=0.063p PE=1.94u AB=31.9135p PB=26.72u AC=31.896634p PC=26.71u NE=5 m=5
R26 GND|TLA|TLB GND|TLA|TLB rsil w=4u l=3u ps=0 b=0 m=1
R27 RFOUT|RFOUT3|TLA|TLB TLA|TLB|VCC1|VCC3 rsil w=4u l=14.5u ps=0 b=0 m=1
R28 GND|TLA|TLB RFIN3|RFOUT2|TLA|TLB rppd w=3u l=6u ps=0 b=0 m=1
R29 RFIN|RFIN1|TLA|TLB RFIN3|RFOUT2|TLA|TLB rppd w=2u l=6.5u ps=0 b=0 m=1
R30 RFIN2|RFOUT1 TLA|TLB|VCC1|VCC31 rppd w=8u l=4.5u ps=0 b=0 m=1
C31 TLA|TLB|VCC2 GND|TLA|TLB cap_cmim w=30u l=60u A=1800p P=180u m=2
C32 TLA|TLB|VCC1|VCC31 GND|TLA|TLB cap_cmim w=30u l=60u A=1800p P=180u m=2
C34 TLA|TLB|VCC1|VCC3 GND|TLA|TLB cap_cmim w=30u l=60u A=1800p P=180u m=2
.ENDS TOP
