* Qucs 25.1.0  C:/Users/rupok_nsl/QucsWorkspace/Final_prj/new_design_netlist.sch

.SUBCKT FMD_QNC_01_LIN_TIA


CDC3 \VCC1 \GND cap_cmim w=20u l=100u A=2000p P=240u m=1
CDC1 \VCC1 \GND cap_cmim w=60u l=60u A=3600p P=240u m=2
CDC24 \VCC2 \GND cap_cmim w=60u l=60u A=3600p P=240u m=2

RRC1 \VCC1 \NET12 rppd w=8.5U l=2U m=1
RRE2 \NET23 \GND rhigh w=8U l=8.2U m=1
RRE3 \NET34 \GND rppd w=4U l=2.9U m=1
RRC4 \VCC2 \RFOUT rppd w=20.6U l=2.1U m=1
QQ11 \NET1 \RFIN \GND \GND npn13G2 AE=0.063p PE=1.94u AB=63.456p PB=45.22u
+ AC=63.429884p PC=45.21u NE=10 m=10
QQ12 \NET12 \VB1 \NET1 \GND npn13G2 AE=0.063p PE=1.94u AB=12.988p PB=15.62u
+ AC=12.976684p PC=15.61u NE=2 m=2
QQ21 \VCC2 \NET12 \NET23 \GND npn13G2 AE=0.063p PE=1.94u AB=31.9135p PB=26.72u
+ AC=31.896634p PC=26.71u NE=5 m=5
QQ31 \NET3 \NET23 \NET34 \GND npn13G2 AE=0.063p PE=1.94u AB=31.9135p PB=26.72u
+ AC=31.896634p PC=26.71u NE=5 m=5
QQ32 \VCC1 \VCC1 \NET3 \GND npn13G2 AE=0.063p PE=1.94u AB=12.988p PB=15.62u
+ AC=12.976684p PC=15.61u NE=2 m=2
QQ41 \NET4 \NET34 \_net0 \GND npn13G2 AE=0.063p PE=1.94u AB=63.456p PB=45.22u
+ AC=63.429884p PC=45.21u NE=10 m=10

CCB1 \VB1 \GND cap_cmim w=30u l=30u A=900p P=120u m=1
CCB2 \VB2 \GND cap_cmim w=30u l=30u A=900p P=120u m=1

QQB11 \VB1 \_net1 \_net2 \GND npn13G2 AE=0.063p PE=1.94u AB=6.6795p PB=11.92u
+ AC=6.670034p PC=11.91u NE=1 m=1
QQB12 \_net3 \_net4 \GND \GND npn13G2 AE=0.063p PE=1.94u AB=6.6795p PB=11.92u
+ AC=6.670034p PC=11.91u NE=1 m=1
QQB21 \VB2 \_net5 \_net6 \GND npn13G2 AE=0.063p PE=1.94u AB=6.6795p PB=11.92u
+ AC=6.670034p PC=11.91u NE=1 m=1
QQB22 \_net7 \_net8 \GND \GND npn13G2 AE=0.063p PE=1.94u AB=6.6795p PB=11.92u
+ AC=6.670034p PC=11.91u NE=1 m=1
RRB1_RB1 \_net1 \VB1 rhigh w=3U l=2U m=1
RRB1_RC1 \VCC1 \VB1 rhigh w=3U l=2.94U m=1
RRB1_RC2 \_net2 \_net3 rhigh w=3U l=2U m=1
RRB1_RB2 \_net4 \_net3 rhigh w=3U l=2U m=1
RRB2_RC1 \VCC2 VB2 rhigh w=3U l=1.94U m=1
RRB2_RB1 \_net5 \VB2 rhigh w=3U l=2U m=1
RRB2_RC2 \_net7 \_net6 rhigh w=3U l=2U m=1
RRB2_RB2 \_net8 \_net7 rhigh w=3U l=2U m=1
QQF \NET23 \NET23 \NETF \GND npn13G2 AE=0.063p PE=1.94u AB=6.6795p PB=11.92u
+ AC=6.670034p PC=11.91u NE=1 m=1
RRF1 \RFIN \NETF rppd w=4U l=13.3U m=1
RRF2 \GND \RFIN rhigh w=4U l=9.9U m=1


RRE4 \_net0 \GND rsil w=18U l=30U m=1
QQ42 \RFOUT \VB2 \NET4 \GND npn13G2 AE=0.063p PE=1.94u AB=25.605p PB=23.02u
+ AC=25.589984p PC=23.01u NE=4 m=4
.END
