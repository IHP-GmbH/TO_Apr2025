.SUBCKT TOP

Cc1 \vcc1 \gnd cap_cmim w=30u l=60u A=1800p P=180u m=2
Cc2 \vcc2 \gnd cap_cmim w=30u l=60u A=1800p P=180u m=2
Cc3 \vcc3 \gnd cap_cmim w=30u l=60u A=1800p P=180u m=2

RRF \RFin \net2 rppd w=2u l=6.5u ps=0 b=0 m=1

RRC1 \vcc1 \net1 rppd w=8u l=4.5u ps=0 b=0 m=1
RRE2 \net2 \gnd rppd w=3u l=6u ps=0 b=0 m=1

RRC3 \vcc3 \RFout rsil w=4u l=14.5u ps=0 b=0 m=1
RRE3 \net3 \gnd rsil w=4u l=3u ps=0 b=0 m=1

Qq1 \net1 \RFin \gnd \gnd npn13G2 AE=0.063p PE=1.94u AB=63.456p PB=45.22u
+ AC=63.429884p PC=45.21u NE=10 m=10
Qq2 \vcc2 \net1 \net2 \gnd npn13G2 AE=0.063p PE=1.94u AB=31.9135p
+ PB=26.72u AC=31.896634p PC=26.71u NE=5 m=5
Qq3 \RFout \net2 \net3 \gnd npn13G2 AE=0.063p PE=1.94u AB=63.456p
+ PB=45.22u AC=63.429884p PC=45.21u NE=10 m=10

.ENDS TOP
