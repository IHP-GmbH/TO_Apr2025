* Extracted by KLayout with SG13G2 LVS runset on : 05/04/2025 05:22

.SUBCKT nmos_200_2
M$1 \$3 \$4 \$2 \$1 rfnmos L=0.36u W=200u AS=120.565p AD=120.565p PS=442.13u
+ PD=442.13u
M$201 \$3 \$6 \$5 \$1 rfnmos L=0.36u W=200u AS=120.565p AD=120.565p PS=442.13u
+ PD=442.13u
.ENDS nmos_200_2
