** sch_path: /home/noritsuna/LNA/202504/lvs/lna_npn_base_lvs.sch
.subckt lna_npn_base_lvs VDD IN OUT VSS VBIAS_IN VBIAS_OUT IBIAS_IN
*.PININFO VDD:B IN:I OUT:O VSS:B VBIAS_IN:B VBIAS_OUT:B IBIAS_IN:B
R2 VBIAS_OUT net1 rppd w=0.5e-6 l=3.6e-6 m=1 b=0
R1 net1 VDD rppd w=0.5e-6 l=1.8e-6 m=1 b=0
R3 net3 IN rsil w=0.5e-6 l=2.4e-6 m=1 b=0
C1 net3 VBIAS_OUT VSS rfcmim w=60.0e-6 l=55.0e-6 wfeed=5.0e-6
M3 net1 net1 VSS VSS rfnmos l=0.36u w=10.0u ng=5
Q1 OUT VDD net2 VSS npn13G2 le=900e-9 we=70.0n m=10
Q2 net2 VBIAS_IN IBIAS_IN VSS npn13G2 le=900e-9 we=70.0n m=10
Q3 OUT VDD net2 VSS npn13G2 le=900e-9 we=70.0n m=10
Q4 net2 VBIAS_IN IBIAS_IN VSS npn13G2 le=900e-9 we=70.0n m=10
Q5 OUT VDD net2 VSS npn13G2 le=900e-9 we=70.0n m=10
Q6 net2 VBIAS_IN IBIAS_IN VSS npn13G2 le=900e-9 we=70.0n m=10
Q7 OUT VDD net2 VSS npn13G2 le=900e-9 we=70.0n m=10
Q8 net2 VBIAS_IN IBIAS_IN VSS npn13G2 le=900e-9 we=70.0n m=10
Q9 OUT VDD net2 VSS npn13G2 le=900e-9 we=70.0n m=10
Q10 net2 VBIAS_IN IBIAS_IN VSS npn13G2 le=900e-9 we=70.0n m=10
Q11 OUT VDD net2 VSS npn13G2 le=900e-9 we=70.0n m=10
Q12 net2 VBIAS_IN IBIAS_IN VSS npn13G2 le=900e-9 we=70.0n m=10
.ends
.end
