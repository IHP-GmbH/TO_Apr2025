* Extracted by KLayout with SG13G2 LVS runset on : 10/04/2025 17:36

.SUBCKT FDM_QNC_00_LN_TIA
C$1 \$I94377 \$1 cap_cmim w=30u l=60u A=1800p P=180u m=2
C$2 \$I94382 \$1 cap_cmim w=30u l=60u A=1800p P=180u m=2
C$5 \$I94381 \$1 cap_cmim w=30u l=60u A=1800p P=180u m=2
R$7 \$I210262 \$I210263 rppd w=2u l=6.5u ps=0 b=0 m=1
R$8 \$1 \$I210266 rsil w=4u l=3u ps=0 b=0 m=1
R$9 \$I210264 \$I94381 rsil w=4u l=14.5u ps=0 b=0 m=1
R$10 \$1 \$I210263 rppd w=3u l=6u ps=0 b=0 m=1
Q$11 \$I94377 \$I210265 \$I210263 \$1 npn13G2 AE=0.063p PE=1.94u AB=31.9135p
+ PB=26.72u AC=31.896634p PC=26.71u NE=5 m=5
R$16 \$I94382 \$I210265 rppd w=8u l=4.5u ps=0 b=0 m=1
Q$17 \$I210264 \$I210263 \$I210266 \$1 npn13G2 AE=0.063p PE=1.94u AB=63.456p
+ PB=45.22u AC=63.429884p PC=45.21u NE=10 m=10
Q$27 \$I210265 \$I210262 \$1 \$1 npn13G2 AE=0.063p PE=1.94u AB=63.456p
+ PB=45.22u AC=63.429884p PC=45.21u NE=10 m=10
.ENDS FDM_QNC_00_LN_TIA
