* Extracted by KLayout with SG13G2 LVS runset on : 04/04/2025 06:36

.SUBCKT TOP
Q$1 \$10816 \$11051 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
Q$21 \$10842 \$11278 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=50.839p PB=37.82u AC=50.816584p PC=37.81u NE=16 m=16
Q$37 \$11022 \$11277 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=50.839p PB=37.82u AC=50.816584p PC=37.81u NE=16 m=16
Q$53 \$17270 \$17494 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=50.839p PB=37.82u AC=50.816584p PC=37.81u NE=16 m=16
Q$69 \$17282 \$17571 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
Q$89 \$17317 \$17495 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=50.839p PB=37.82u AC=50.816584p PC=37.81u NE=16 m=16
Q$105 \$24255 \$24680 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
Q$125 \$24404 \$24900 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=50.839p PB=37.82u AC=50.816584p PC=37.81u NE=16 m=16
Q$141 \$24461 \$24899 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=50.839p PB=37.82u AC=50.816584p PC=37.81u NE=16 m=16
Q$157 \$30799 \$30965 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=50.839p PB=37.82u AC=50.816584p PC=37.81u NE=16 m=16
Q$173 \$30962 \$31252 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=63.456p PB=45.22u AC=63.429884p PC=45.21u NE=20 m=20
Q$193 \$30966 \$31192 RFIN|RFOUT|VSS RFIN|RFOUT|VSS npn13G2 AE=0.063p PE=1.94u
+ AB=50.839p PB=37.82u AC=50.816584p PC=37.81u NE=16 m=16
R$209 \$11051 VBB2 rsil w=2u l=12u ps=0 b=0 m=1
R$210 \$11278 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$211 \$11277 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$212 RFIN|RFOUT|VSS RFIN|RFOUT|VSS rsil w=2.04u l=28u ps=0 b=0 m=6
R$214 VBB1 \$17494 rsil w=2u l=11u ps=0 b=0 m=1
R$215 VBB1 \$17495 rsil w=2u l=11u ps=0 b=0 m=1
R$216 VBB2 \$17571 rsil w=2u l=12u ps=0 b=0 m=1
R$219 \$24680 VBB2 rsil w=2u l=12u ps=0 b=0 m=1
R$220 \$24900 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$221 \$24899 VBB1 rsil w=2u l=11u ps=0 b=0 m=1
R$224 VBB1 \$30965 rsil w=2u l=11u ps=0 b=0 m=1
R$225 VBB1 \$31192 rsil w=2u l=11u ps=0 b=0 m=1
R$226 VBB2 \$31252 rsil w=2u l=12u ps=0 b=0 m=1
R$227 VCC2 \$10816 rppd w=35u l=0.5u ps=0 b=0 m=1
R$228 VCC1 \$10842 rppd w=35u l=0.5u ps=0 b=0 m=1
R$229 VCC1 \$11022 rppd w=35u l=0.5u ps=0 b=0 m=1
R$230 \$17270 VCC1$1 rppd w=35u l=0.5u ps=0 b=0 m=1
R$231 \$17317 VCC1$1 rppd w=35u l=0.5u ps=0 b=0 m=1
R$232 \$17282 VCC2 rppd w=35u l=0.5u ps=0 b=0 m=1
R$233 VCC2 \$24255 rppd w=35u l=0.5u ps=0 b=0 m=1
R$234 VCC1$1 \$24404 rppd w=35u l=0.5u ps=0 b=0 m=1
R$235 VCC1$1 \$24461 rppd w=35u l=0.5u ps=0 b=0 m=1
R$236 \$30799 VCC1$1 rppd w=35u l=0.5u ps=0 b=0 m=1
R$237 \$30966 VCC1$1 rppd w=35u l=0.5u ps=0 b=0 m=1
R$238 \$30962 VCC2$1 rppd w=35u l=0.5u ps=0 b=0 m=1
C$239 VCC1$1 RFIN|RFOUT|VSS cap_cmim w=15u l=30u A=450p P=90u m=16
C$242 VCC1 RFIN|RFOUT|VSS cap_cmim w=15u l=30u A=450p P=90u m=4
C$247 VCC2$1 RFIN|RFOUT|VSS cap_cmim w=15u l=30u A=450p P=90u m=2
C$249 VCC2 RFIN|RFOUT|VSS cap_cmim w=15u l=30u A=450p P=90u m=10
.ENDS TOP
