* Extracted by KLayout with SG13G2 LVS runset on : 05/04/2025 05:18

.SUBCKT INP_LVS
C$1 \$4 \$3 \$1 rfcmim w=60u l=55u A=3300p P=230u m=1 wfeed=5u
R$2 \$4 \$8 rsil w=0.5u l=2.4u ps=0 b=0 m=1
.ENDS INP_LVS
