* Qucs 25.1.0  /headless/QucsWorkspace/Ikram_prj/3_Stage_2nd_Design.sch
.SUBCKT Sub_SPfile_X3 1 2 3
R1N 1 10 -50
R1P 10 11 100
R2N 2 20 -50
R2P 20 21 100

A11 %vd(10 3) %vd(11, 12) xfer1
.model xfer1 xfer R_I=true table=[
+ 0Hz 0.00482376 0
+ 1e+08Hz 0.00482395 1.93737e-06
+ 2e+08Hz 0.00482452 3.86743e-06
+ 3e+08Hz 0.00482548 5.78289e-06
+ 4e+08Hz 0.00482681 7.67645e-06
+ 5e+08Hz 0.00482853 9.54082e-06
+ 6e+08Hz 0.00483063 1.13687e-05
+ 7e+08Hz 0.0048331 1.3153e-05
+ 8e+08Hz 0.00483596 1.48863e-05
+ 9e+08Hz 0.00483919 1.65614e-05
+ 1e+09Hz 0.0048428 1.81712e-05
+ 1.1e+09Hz 0.00484679 1.97086e-05
+ 1.2e+09Hz 0.00485114 2.11664e-05
+ 1.3e+09Hz 0.00485587 2.25375e-05
+ 1.4e+09Hz 0.00486097 2.3815e-05
+ 1.5e+09Hz 0.00486643 2.49917e-05
+ 1.6e+09Hz 0.00487226 2.60609e-05
+ 1.7e+09Hz 0.00487846 2.70156e-05
+ 1.8e+09Hz 0.00488501 2.78489e-05
+ 1.9e+09Hz 0.00489192 2.85541e-05
+ 2e+09Hz 0.00489919 2.91245e-05
+ 2.1e+09Hz 0.00490681 2.95534e-05
+ 2.2e+09Hz 0.00491478 2.98342e-05
+ 2.3e+09Hz 0.00492309 2.99605e-05
+ 2.4e+09Hz 0.00493175 2.99257e-05
+ 2.5e+09Hz 0.00494075 2.97235e-05
+ 2.6e+09Hz 0.00495008 2.93477e-05
+ 2.7e+09Hz 0.00495975 2.87919e-05
+ 2.8e+09Hz 0.00496975 2.80502e-05
+ 2.9e+09Hz 0.00498007 2.71164e-05
+ 3e+09Hz 0.00499071 2.59846e-05
+ 3.1e+09Hz 0.00500167 2.4649e-05
+ 3.2e+09Hz 0.00501294 2.31038e-05
+ 3.3e+09Hz 0.00502452 2.13433e-05
+ 3.4e+09Hz 0.0050364 1.93619e-05
+ 3.5e+09Hz 0.00504859 1.71543e-05
+ 3.6e+09Hz 0.00506107 1.4715e-05
+ 3.7e+09Hz 0.00507383 1.20388e-05
+ 3.8e+09Hz 0.00508689 9.12049e-06
+ 3.9e+09Hz 0.00510022 5.9551e-06
+ 4e+09Hz 0.00511383 2.53768e-06
+ 4.1e+09Hz 0.00512771 -1.13658e-06
+ 4.2e+09Hz 0.00514185 -5.07238e-06
+ 4.3e+09Hz 0.00515626 -9.2743e-06
+ 4.4e+09Hz 0.00517091 -1.37468e-05
+ 4.5e+09Hz 0.00518582 -1.84942e-05
+ 4.6e+09Hz 0.00520097 -2.35208e-05
+ 4.7e+09Hz 0.00521636 -2.88306e-05
+ 4.8e+09Hz 0.00523198 -3.44276e-05
+ 4.9e+09Hz 0.00524782 -4.03157e-05
+ 5e+09Hz 0.00526389 -4.64986e-05
+ 5.1e+09Hz 0.00528017 -5.29798e-05
+ 5.2e+09Hz 0.00529666 -5.97629e-05
+ 5.3e+09Hz 0.00531335 -6.68512e-05
+ 5.4e+09Hz 0.00533024 -7.42479e-05
+ 5.5e+09Hz 0.00534732 -8.1956e-05
+ 5.6e+09Hz 0.00536459 -8.99785e-05
+ 5.7e+09Hz 0.00538203 -9.83183e-05
+ 5.8e+09Hz 0.00539964 -0.000106978
+ 5.9e+09Hz 0.00541742 -0.00011596
+ 6e+09Hz 0.00543536 -0.000125267
+ 6.1e+09Hz 0.00545346 -0.000134901
+ 6.2e+09Hz 0.0054717 -0.000144864
+ 6.3e+09Hz 0.00549008 -0.000155159
+ 6.4e+09Hz 0.00550859 -0.000165787
+ 6.5e+09Hz 0.00552723 -0.00017675
+ 6.6e+09Hz 0.005546 -0.000188049
+ 6.7e+09Hz 0.00556488 -0.000199686
+ 6.8e+09Hz 0.00558387 -0.000211663
+ 6.9e+09Hz 0.00560296 -0.00022398
+ 7e+09Hz 0.00562214 -0.000236638
+ 7.1e+09Hz 0.00564142 -0.000249639
+ 7.2e+09Hz 0.00566077 -0.000262984
+ 7.3e+09Hz 0.00568021 -0.000276673
+ 7.4e+09Hz 0.00569971 -0.000290706
+ 7.5e+09Hz 0.00571928 -0.000305084
+ 7.6e+09Hz 0.00573891 -0.000319807
+ 7.7e+09Hz 0.00575858 -0.000334876
+ 7.8e+09Hz 0.0057783 -0.00035029
+ 7.9e+09Hz 0.00579806 -0.00036605
+ 8e+09Hz 0.00581785 -0.000382155
+ 8.1e+09Hz 0.00583767 -0.000398604
+ 8.2e+09Hz 0.00585751 -0.000415398
+ 8.3e+09Hz 0.00587736 -0.000432536
+ 8.4e+09Hz 0.00589721 -0.000450016
+ 8.5e+09Hz 0.00591707 -0.000467839
+ 8.6e+09Hz 0.00593692 -0.000486003
+ 8.7e+09Hz 0.00595676 -0.000504507
+ 8.8e+09Hz 0.00597658 -0.00052335
+ 8.9e+09Hz 0.00599638 -0.000542531
+ 9e+09Hz 0.00601615 -0.000562048
+ 9.1e+09Hz 0.00603589 -0.0005819
+ 9.2e+09Hz 0.00605558 -0.000602085
+ 9.3e+09Hz 0.00607523 -0.000622601
+ 9.4e+09Hz 0.00609483 -0.000643447
+ 9.5e+09Hz 0.00611437 -0.00066462
+ 9.6e+09Hz 0.00613384 -0.000686119
+ 9.7e+09Hz 0.00615324 -0.000707941
+ 9.8e+09Hz 0.00617257 -0.000730084
+ 9.9e+09Hz 0.00619183 -0.000752546
+ 1e+10Hz 0.00621099 -0.000775324
+ 1.01e+10Hz 0.00623007 -0.000798416
+ 1.02e+10Hz 0.00624905 -0.000821819
+ 1.03e+10Hz 0.00626793 -0.000845531
+ 1.04e+10Hz 0.0062867 -0.000869548
+ 1.05e+10Hz 0.00630536 -0.000893868
+ 1.06e+10Hz 0.00632391 -0.000918487
+ 1.07e+10Hz 0.00634234 -0.000943403
+ 1.08e+10Hz 0.00636064 -0.000968612
+ 1.09e+10Hz 0.00637881 -0.000994112
+ 1.1e+10Hz 0.00639685 -0.0010199
+ 1.11e+10Hz 0.00641475 -0.00104597
+ 1.12e+10Hz 0.00643251 -0.00107232
+ 1.13e+10Hz 0.00645012 -0.00109895
+ 1.14e+10Hz 0.00646758 -0.00112585
+ 1.15e+10Hz 0.00648489 -0.00115302
+ 1.16e+10Hz 0.00650203 -0.00118045
+ 1.17e+10Hz 0.00651902 -0.00120815
+ 1.18e+10Hz 0.00653583 -0.00123611
+ 1.19e+10Hz 0.00655248 -0.00126432
+ 1.2e+10Hz 0.00656895 -0.00129278
+ 1.21e+10Hz 0.00658524 -0.00132148
+ 1.22e+10Hz 0.00660135 -0.00135043
+ 1.23e+10Hz 0.00661728 -0.00137962
+ 1.24e+10Hz 0.00663302 -0.00140904
+ 1.25e+10Hz 0.00664857 -0.00143869
+ 1.26e+10Hz 0.00666392 -0.00146857
+ 1.27e+10Hz 0.00667908 -0.00149867
+ 1.28e+10Hz 0.00669404 -0.00152899
+ 1.29e+10Hz 0.00670879 -0.00155951
+ 1.3e+10Hz 0.00672335 -0.00159025
+ 1.31e+10Hz 0.00673769 -0.00162119
+ 1.32e+10Hz 0.00675182 -0.00165234
+ 1.33e+10Hz 0.00676574 -0.00168367
+ 1.34e+10Hz 0.00677945 -0.0017152
+ 1.35e+10Hz 0.00679294 -0.00174692
+ 1.36e+10Hz 0.00680621 -0.00177882
+ 1.37e+10Hz 0.00681926 -0.00181089
+ 1.38e+10Hz 0.00683208 -0.00184314
+ 1.39e+10Hz 0.00684468 -0.00187555
+ 1.4e+10Hz 0.00685706 -0.00190813
+ 1.41e+10Hz 0.00686921 -0.00194087
+ 1.42e+10Hz 0.00688113 -0.00197377
+ 1.43e+10Hz 0.00689282 -0.00200681
+ 1.44e+10Hz 0.00690427 -0.00204001
+ 1.45e+10Hz 0.0069155 -0.00207334
+ 1.46e+10Hz 0.00692649 -0.00210681
+ 1.47e+10Hz 0.00693724 -0.00214041
+ 1.48e+10Hz 0.00694776 -0.00217414
+ 1.49e+10Hz 0.00695804 -0.00220799
+ 1.5e+10Hz 0.00696809 -0.00224196
+ 1.51e+10Hz 0.0069779 -0.00227604
+ 1.52e+10Hz 0.00698746 -0.00231024
+ 1.53e+10Hz 0.00699679 -0.00234454
+ 1.54e+10Hz 0.00700588 -0.00237894
+ 1.55e+10Hz 0.00701474 -0.00241344
+ 1.56e+10Hz 0.00702335 -0.00244802
+ 1.57e+10Hz 0.00703172 -0.0024827
+ 1.58e+10Hz 0.00703985 -0.00251746
+ 1.59e+10Hz 0.00704774 -0.0025523
+ 1.6e+10Hz 0.0070554 -0.00258721
+ 1.61e+10Hz 0.00706281 -0.00262219
+ 1.62e+10Hz 0.00706999 -0.00265724
+ 1.63e+10Hz 0.00707693 -0.00269235
+ 1.64e+10Hz 0.00708363 -0.00272752
+ 1.65e+10Hz 0.00709009 -0.00276274
+ 1.66e+10Hz 0.00709632 -0.00279801
+ 1.67e+10Hz 0.00710231 -0.00283332
+ 1.68e+10Hz 0.00710806 -0.00286868
+ 1.69e+10Hz 0.00711359 -0.00290407
+ 1.7e+10Hz 0.00711888 -0.0029395
+ 1.71e+10Hz 0.00712393 -0.00297496
+ 1.72e+10Hz 0.00712876 -0.00301044
+ 1.73e+10Hz 0.00713336 -0.00304594
+ 1.74e+10Hz 0.00713773 -0.00308147
+ 1.75e+10Hz 0.00714187 -0.003117
+ 1.76e+10Hz 0.00714579 -0.00315255
+ 1.77e+10Hz 0.00714948 -0.0031881
+ 1.78e+10Hz 0.00715295 -0.00322366
+ 1.79e+10Hz 0.00715621 -0.00325922
+ 1.8e+10Hz 0.00715924 -0.00329477
+ 1.81e+10Hz 0.00716205 -0.00333032
+ 1.82e+10Hz 0.00716465 -0.00336586
+ 1.83e+10Hz 0.00716703 -0.00340138
+ 1.84e+10Hz 0.00716921 -0.00343689
+ 1.85e+10Hz 0.00717117 -0.00347238
+ 1.86e+10Hz 0.00717293 -0.00350784
+ 1.87e+10Hz 0.00717447 -0.00354328
+ 1.88e+10Hz 0.00717582 -0.00357869
+ 1.89e+10Hz 0.00717696 -0.00361407
+ 1.9e+10Hz 0.00717791 -0.00364941
+ 1.91e+10Hz 0.00717866 -0.00368472
+ 1.92e+10Hz 0.00717921 -0.00371999
+ 1.93e+10Hz 0.00717957 -0.00375522
+ 1.94e+10Hz 0.00717974 -0.0037904
+ 1.95e+10Hz 0.00717972 -0.00382553
+ 1.96e+10Hz 0.00717951 -0.00386061
+ 1.97e+10Hz 0.00717912 -0.00389564
+ 1.98e+10Hz 0.00717856 -0.00393062
+ 1.99e+10Hz 0.00717781 -0.00396554
+ 2e+10Hz 0.00717689 -0.0040004
+ 2.01e+10Hz 0.00717579 -0.0040352
+ 2.02e+10Hz 0.00717453 -0.00406994
+ 2.03e+10Hz 0.00717309 -0.00410461
+ 2.04e+10Hz 0.00717149 -0.00413921
+ 2.05e+10Hz 0.00716973 -0.00417375
+ 2.06e+10Hz 0.00716781 -0.00420822
+ 2.07e+10Hz 0.00716573 -0.00424261
+ 2.08e+10Hz 0.0071635 -0.00427693
+ 2.09e+10Hz 0.00716111 -0.00431118
+ 2.1e+10Hz 0.00715858 -0.00434535
+ 2.11e+10Hz 0.0071559 -0.00437944
+ 2.12e+10Hz 0.00715308 -0.00441345
+ 2.13e+10Hz 0.00715011 -0.00444738
+ 2.14e+10Hz 0.00714701 -0.00448123
+ 2.15e+10Hz 0.00714377 -0.004515
+ 2.16e+10Hz 0.0071404 -0.00454868
+ 2.17e+10Hz 0.0071369 -0.00458228
+ 2.18e+10Hz 0.00713327 -0.0046158
+ 2.19e+10Hz 0.00712952 -0.00464922
+ 2.2e+10Hz 0.00712565 -0.00468256
+ 2.21e+10Hz 0.00712165 -0.00471582
+ 2.22e+10Hz 0.00711755 -0.00474898
+ 2.23e+10Hz 0.00711332 -0.00478206
+ 2.24e+10Hz 0.00710899 -0.00481504
+ 2.25e+10Hz 0.00710455 -0.00484794
+ 2.26e+10Hz 0.00710001 -0.00488074
+ 2.27e+10Hz 0.00709536 -0.00491346
+ 2.28e+10Hz 0.00709061 -0.00494608
+ 2.29e+10Hz 0.00708577 -0.00497862
+ 2.3e+10Hz 0.00708083 -0.00501106
+ 2.31e+10Hz 0.00707579 -0.00504341
+ 2.32e+10Hz 0.00707067 -0.00507567
+ 2.33e+10Hz 0.00706546 -0.00510784
+ 2.34e+10Hz 0.00706017 -0.00513992
+ 2.35e+10Hz 0.0070548 -0.00517191
+ 2.36e+10Hz 0.00704934 -0.00520381
+ 2.37e+10Hz 0.00704381 -0.00523561
+ 2.38e+10Hz 0.00703821 -0.00526733
+ 2.39e+10Hz 0.00703253 -0.00529896
+ 2.4e+10Hz 0.00702678 -0.0053305
+ 2.41e+10Hz 0.00702097 -0.00536195
+ 2.42e+10Hz 0.00701509 -0.00539332
+ 2.43e+10Hz 0.00700915 -0.00542459
+ 2.44e+10Hz 0.00700315 -0.00545578
+ 2.45e+10Hz 0.00699709 -0.00548688
+ 2.46e+10Hz 0.00699097 -0.0055179
+ 2.47e+10Hz 0.0069848 -0.00554884
+ 2.48e+10Hz 0.00697857 -0.00557969
+ 2.49e+10Hz 0.0069723 -0.00561046
+ 2.5e+10Hz 0.00696598 -0.00564114
+ 2.51e+10Hz 0.00695961 -0.00567175
+ 2.52e+10Hz 0.0069532 -0.00570228
+ 2.53e+10Hz 0.00694675 -0.00573272
+ 2.54e+10Hz 0.00694026 -0.00576309
+ 2.55e+10Hz 0.00693372 -0.00579339
+ 2.56e+10Hz 0.00692716 -0.00582361
+ 2.57e+10Hz 0.00692055 -0.00585375
+ 2.58e+10Hz 0.00691392 -0.00588382
+ 2.59e+10Hz 0.00690725 -0.00591382
+ 2.6e+10Hz 0.00690055 -0.00594375
+ 2.61e+10Hz 0.00689382 -0.00597361
+ 2.62e+10Hz 0.00688707 -0.0060034
+ 2.63e+10Hz 0.00688029 -0.00603313
+ 2.64e+10Hz 0.00687348 -0.00606279
+ 2.65e+10Hz 0.00686665 -0.00609239
+ 2.66e+10Hz 0.0068598 -0.00612192
+ 2.67e+10Hz 0.00685293 -0.00615139
+ 2.68e+10Hz 0.00684605 -0.00618081
+ 2.69e+10Hz 0.00683914 -0.00621016
+ 2.7e+10Hz 0.00683221 -0.00623947
+ 2.71e+10Hz 0.00682527 -0.00626871
+ 2.72e+10Hz 0.00681832 -0.0062979
+ 2.73e+10Hz 0.00681135 -0.00632704
+ 2.74e+10Hz 0.00680436 -0.00635613
+ 2.75e+10Hz 0.00679737 -0.00638517
+ 2.76e+10Hz 0.00679036 -0.00641417
+ 2.77e+10Hz 0.00678335 -0.00644311
+ 2.78e+10Hz 0.00677632 -0.00647202
+ 2.79e+10Hz 0.00676928 -0.00650088
+ 2.8e+10Hz 0.00676224 -0.0065297
+ 2.81e+10Hz 0.00675518 -0.00655848
+ 2.82e+10Hz 0.00674812 -0.00658722
+ 2.83e+10Hz 0.00674105 -0.00661593
+ 2.84e+10Hz 0.00673398 -0.0066446
+ 2.85e+10Hz 0.00672689 -0.00667324
+ 2.86e+10Hz 0.0067198 -0.00670184
+ 2.87e+10Hz 0.00671271 -0.00673042
+ 2.88e+10Hz 0.00670561 -0.00675897
+ 2.89e+10Hz 0.00669851 -0.00678749
+ 2.9e+10Hz 0.00669139 -0.00681599
+ 2.91e+10Hz 0.00668428 -0.00684446
+ 2.92e+10Hz 0.00667716 -0.00687291
+ 2.93e+10Hz 0.00667003 -0.00690134
+ 2.94e+10Hz 0.0066629 -0.00692975
+ 2.95e+10Hz 0.00665576 -0.00695814
+ 2.96e+10Hz 0.00664862 -0.00698652
+ 2.97e+10Hz 0.00664148 -0.00701488
+ 2.98e+10Hz 0.00663432 -0.00704322
+ 2.99e+10Hz 0.00662716 -0.00707156
+ 3e+10Hz 0.00662 -0.00709988
+ 3.01e+10Hz 0.00661283 -0.0071282
+ 3.02e+10Hz 0.00660565 -0.00715651
+ 3.03e+10Hz 0.00659846 -0.00718481
+ 3.04e+10Hz 0.00659127 -0.0072131
+ 3.05e+10Hz 0.00658407 -0.00724139
+ 3.06e+10Hz 0.00657686 -0.00726968
+ 3.07e+10Hz 0.00656964 -0.00729797
+ 3.08e+10Hz 0.00656241 -0.00732626
+ 3.09e+10Hz 0.00655517 -0.00735454
+ 3.1e+10Hz 0.00654792 -0.00738283
+ 3.11e+10Hz 0.00654066 -0.00741113
+ 3.12e+10Hz 0.00653339 -0.00743943
+ 3.13e+10Hz 0.0065261 -0.00746773
+ 3.14e+10Hz 0.0065188 -0.00749604
+ 3.15e+10Hz 0.00651149 -0.00752436
+ 3.16e+10Hz 0.00650416 -0.00755268
+ 3.17e+10Hz 0.00649682 -0.00758102
+ 3.18e+10Hz 0.00648946 -0.00760937
+ 3.19e+10Hz 0.00648208 -0.00763772
+ 3.2e+10Hz 0.00647468 -0.00766609
+ 3.21e+10Hz 0.00646726 -0.00769448
+ 3.22e+10Hz 0.00645983 -0.00772288
+ 3.23e+10Hz 0.00645237 -0.00775129
+ 3.24e+10Hz 0.00644489 -0.00777972
+ 3.25e+10Hz 0.00643738 -0.00780816
+ 3.26e+10Hz 0.00642986 -0.00783662
+ 3.27e+10Hz 0.0064223 -0.0078651
+ 3.28e+10Hz 0.00641473 -0.0078936
+ 3.29e+10Hz 0.00640712 -0.00792212
+ 3.3e+10Hz 0.00639949 -0.00795065
+ 3.31e+10Hz 0.00639182 -0.00797921
+ 3.32e+10Hz 0.00638413 -0.00800779
+ 3.33e+10Hz 0.00637641 -0.00803639
+ 3.34e+10Hz 0.00636865 -0.008065
+ 3.35e+10Hz 0.00636086 -0.00809365
+ 3.36e+10Hz 0.00635303 -0.00812231
+ 3.37e+10Hz 0.00634517 -0.008151
+ 3.38e+10Hz 0.00633728 -0.0081797
+ 3.39e+10Hz 0.00632934 -0.00820844
+ 3.4e+10Hz 0.00632137 -0.00823719
+ 3.41e+10Hz 0.00631335 -0.00826597
+ 3.42e+10Hz 0.0063053 -0.00829477
+ 3.43e+10Hz 0.0062972 -0.0083236
+ 3.44e+10Hz 0.00628906 -0.00835245
+ 3.45e+10Hz 0.00628087 -0.00838133
+ 3.46e+10Hz 0.00627264 -0.00841022
+ 3.47e+10Hz 0.00626436 -0.00843915
+ 3.48e+10Hz 0.00625603 -0.00846809
+ 3.49e+10Hz 0.00624766 -0.00849706
+ 3.5e+10Hz 0.00623923 -0.00852606
+ 3.51e+10Hz 0.00623075 -0.00855508
+ 3.52e+10Hz 0.00622222 -0.00858412
+ 3.53e+10Hz 0.00621364 -0.00861318
+ 3.54e+10Hz 0.006205 -0.00864227
+ 3.55e+10Hz 0.00619631 -0.00867138
+ 3.56e+10Hz 0.00618756 -0.00870052
+ 3.57e+10Hz 0.00617875 -0.00872968
+ 3.58e+10Hz 0.00616989 -0.00875885
+ 3.59e+10Hz 0.00616096 -0.00878805
+ 3.6e+10Hz 0.00615198 -0.00881728
+ 3.61e+10Hz 0.00614293 -0.00884652
+ 3.62e+10Hz 0.00613382 -0.00887578
+ 3.63e+10Hz 0.00612464 -0.00890507
+ 3.64e+10Hz 0.00611541 -0.00893437
+ 3.65e+10Hz 0.0061061 -0.00896369
+ 3.66e+10Hz 0.00609673 -0.00899303
+ 3.67e+10Hz 0.00608729 -0.00902239
+ 3.68e+10Hz 0.00607778 -0.00905177
+ 3.69e+10Hz 0.00606821 -0.00908116
+ 3.7e+10Hz 0.00605856 -0.00911057
+ 3.71e+10Hz 0.00604885 -0.00913999
+ 3.72e+10Hz 0.00603906 -0.00916943
+ 3.73e+10Hz 0.0060292 -0.00919888
+ 3.74e+10Hz 0.00601926 -0.00922835
+ 3.75e+10Hz 0.00600926 -0.00925783
+ 3.76e+10Hz 0.00599917 -0.00928732
+ 3.77e+10Hz 0.00598901 -0.00931682
+ 3.78e+10Hz 0.00597878 -0.00934633
+ 3.79e+10Hz 0.00596847 -0.00937585
+ 3.8e+10Hz 0.00595808 -0.00940538
+ 3.81e+10Hz 0.00594761 -0.00943492
+ 3.82e+10Hz 0.00593707 -0.00946447
+ 3.83e+10Hz 0.00592644 -0.00949402
+ 3.84e+10Hz 0.00591574 -0.00952358
+ 3.85e+10Hz 0.00590495 -0.00955314
+ 3.86e+10Hz 0.00589408 -0.0095827
+ 3.87e+10Hz 0.00588314 -0.00961227
+ 3.88e+10Hz 0.00587211 -0.00964184
+ 3.89e+10Hz 0.00586099 -0.00967141
+ 3.9e+10Hz 0.0058498 -0.00970098
+ 3.91e+10Hz 0.00583852 -0.00973055
+ 3.92e+10Hz 0.00582716 -0.00976011
+ 3.93e+10Hz 0.00581571 -0.00978968
+ 3.94e+10Hz 0.00580418 -0.00981924
+ 3.95e+10Hz 0.00579257 -0.00984879
+ 3.96e+10Hz 0.00578087 -0.00987834
+ 3.97e+10Hz 0.00576908 -0.00990788
+ 3.98e+10Hz 0.00575722 -0.00993741
+ 3.99e+10Hz 0.00574526 -0.00996694
+ 4e+10Hz 0.00573322 -0.00999645
+ 4.01e+10Hz 0.00572109 -0.010026
+ 4.02e+10Hz 0.00570888 -0.0100554
+ 4.03e+10Hz 0.00569658 -0.0100849
+ 4.04e+10Hz 0.00568419 -0.0101144
+ 4.05e+10Hz 0.00567172 -0.0101438
+ 4.06e+10Hz 0.00565916 -0.0101733
+ 4.07e+10Hz 0.00564652 -0.0102027
+ 4.08e+10Hz 0.00563379 -0.0102321
+ 4.09e+10Hz 0.00562097 -0.0102615
+ 4.1e+10Hz 0.00560807 -0.0102908
+ 4.11e+10Hz 0.00559508 -0.0103202
+ 4.12e+10Hz 0.00558201 -0.0103495
+ 4.13e+10Hz 0.00556884 -0.0103788
+ 4.14e+10Hz 0.0055556 -0.010408
+ 4.15e+10Hz 0.00554227 -0.0104373
+ 4.16e+10Hz 0.00552885 -0.0104665
+ 4.17e+10Hz 0.00551534 -0.0104957
+ 4.18e+10Hz 0.00550176 -0.0105248
+ 4.19e+10Hz 0.00548809 -0.010554
+ 4.2e+10Hz 0.00547433 -0.0105831
+ 4.21e+10Hz 0.00546049 -0.0106121
+ 4.22e+10Hz 0.00544656 -0.0106412
+ 4.23e+10Hz 0.00543256 -0.0106702
+ 4.24e+10Hz 0.00541846 -0.0106992
+ 4.25e+10Hz 0.00540429 -0.0107281
+ 4.26e+10Hz 0.00539004 -0.010757
+ 4.27e+10Hz 0.0053757 -0.0107859
+ 4.28e+10Hz 0.00536128 -0.0108147
+ 4.29e+10Hz 0.00534678 -0.0108435
+ 4.3e+10Hz 0.0053322 -0.0108723
+ 4.31e+10Hz 0.00531754 -0.010901
+ 4.32e+10Hz 0.0053028 -0.0109297
+ 4.33e+10Hz 0.00528798 -0.0109583
+ 4.34e+10Hz 0.00527308 -0.0109869
+ 4.35e+10Hz 0.00525811 -0.0110154
+ 4.36e+10Hz 0.00524306 -0.0110439
+ 4.37e+10Hz 0.00522793 -0.0110724
+ 4.38e+10Hz 0.00521272 -0.0111008
+ 4.39e+10Hz 0.00519744 -0.0111292
+ 4.4e+10Hz 0.00518209 -0.0111575
+ 4.41e+10Hz 0.00516666 -0.0111858
+ 4.42e+10Hz 0.00515116 -0.011214
+ 4.43e+10Hz 0.00513558 -0.0112422
+ 4.44e+10Hz 0.00511993 -0.0112703
+ 4.45e+10Hz 0.00510421 -0.0112984
+ 4.46e+10Hz 0.00508842 -0.0113265
+ 4.47e+10Hz 0.00507256 -0.0113545
+ 4.48e+10Hz 0.00505663 -0.0113824
+ 4.49e+10Hz 0.00504063 -0.0114103
+ 4.5e+10Hz 0.00502457 -0.0114381
+ 4.51e+10Hz 0.00500843 -0.0114659
+ 4.52e+10Hz 0.00499223 -0.0114936
+ 4.53e+10Hz 0.00497597 -0.0115213
+ 4.54e+10Hz 0.00495964 -0.0115489
+ 4.55e+10Hz 0.00494324 -0.0115765
+ 4.56e+10Hz 0.00492678 -0.011604
+ 4.57e+10Hz 0.00491026 -0.0116314
+ 4.58e+10Hz 0.00489368 -0.0116588
+ 4.59e+10Hz 0.00487703 -0.0116862
+ 4.6e+10Hz 0.00486033 -0.0117135
+ 4.61e+10Hz 0.00484356 -0.0117407
+ 4.62e+10Hz 0.00482674 -0.0117679
+ 4.63e+10Hz 0.00480986 -0.011795
+ 4.64e+10Hz 0.00479292 -0.011822
+ 4.65e+10Hz 0.00477592 -0.011849
+ 4.66e+10Hz 0.00475887 -0.011876
+ 4.67e+10Hz 0.00474177 -0.0119029
+ 4.68e+10Hz 0.00472461 -0.0119297
+ 4.69e+10Hz 0.0047074 -0.0119565
+ 4.7e+10Hz 0.00469013 -0.0119832
+ 4.71e+10Hz 0.00467281 -0.0120098
+ 4.72e+10Hz 0.00465544 -0.0120364
+ 4.73e+10Hz 0.00463803 -0.012063
+ 4.74e+10Hz 0.00462056 -0.0120895
+ 4.75e+10Hz 0.00460304 -0.0121159
+ 4.76e+10Hz 0.00458548 -0.0121422
+ 4.77e+10Hz 0.00456787 -0.0121685
+ 4.78e+10Hz 0.00455021 -0.0121948
+ 4.79e+10Hz 0.00453251 -0.012221
+ 4.8e+10Hz 0.00451476 -0.0122471
+ 4.81e+10Hz 0.00449697 -0.0122732
+ 4.82e+10Hz 0.00447914 -0.0122992
+ 4.83e+10Hz 0.00446126 -0.0123251
+ 4.84e+10Hz 0.00444334 -0.012351
+ 4.85e+10Hz 0.00442538 -0.0123769
+ 4.86e+10Hz 0.00440738 -0.0124027
+ 4.87e+10Hz 0.00438934 -0.0124284
+ 4.88e+10Hz 0.00437126 -0.0124541
+ 4.89e+10Hz 0.00435314 -0.0124797
+ 4.9e+10Hz 0.00433498 -0.0125052
+ 4.91e+10Hz 0.00431679 -0.0125307
+ 4.92e+10Hz 0.00429856 -0.0125561
+ 4.93e+10Hz 0.0042803 -0.0125815
+ 4.94e+10Hz 0.004262 -0.0126068
+ 4.95e+10Hz 0.00424366 -0.0126321
+ 4.96e+10Hz 0.00422529 -0.0126573
+ 4.97e+10Hz 0.00420689 -0.0126825
+ 4.98e+10Hz 0.00418846 -0.0127076
+ 4.99e+10Hz 0.00416999 -0.0127326
+ 5e+10Hz 0.00415149 -0.0127576
+ 5.01e+10Hz 0.00413296 -0.0127826
+ 5.02e+10Hz 0.0041144 -0.0128074
+ 5.03e+10Hz 0.00409581 -0.0128323
+ 5.04e+10Hz 0.00407719 -0.0128571
+ 5.05e+10Hz 0.00405854 -0.0128818
+ 5.06e+10Hz 0.00403987 -0.0129065
+ 5.07e+10Hz 0.00402116 -0.0129311
+ 5.08e+10Hz 0.00400243 -0.0129556
+ 5.09e+10Hz 0.00398367 -0.0129802
+ 5.1e+10Hz 0.00396488 -0.0130046
+ 5.11e+10Hz 0.00394607 -0.013029
+ 5.12e+10Hz 0.00392723 -0.0130534
+ 5.13e+10Hz 0.00390836 -0.0130777
+ 5.14e+10Hz 0.00388947 -0.013102
+ 5.15e+10Hz 0.00387056 -0.0131262
+ 5.16e+10Hz 0.00385162 -0.0131504
+ 5.17e+10Hz 0.00383265 -0.0131745
+ 5.18e+10Hz 0.00381367 -0.0131986
+ 5.19e+10Hz 0.00379466 -0.0132226
+ 5.2e+10Hz 0.00377562 -0.0132466
+ 5.21e+10Hz 0.00375656 -0.0132705
+ 5.22e+10Hz 0.00373748 -0.0132944
+ 5.23e+10Hz 0.00371838 -0.0133183
+ 5.24e+10Hz 0.00369925 -0.0133421
+ 5.25e+10Hz 0.00368011 -0.0133658
+ 5.26e+10Hz 0.00366094 -0.0133896
+ 5.27e+10Hz 0.00364175 -0.0134132
+ 5.28e+10Hz 0.00362253 -0.0134369
+ 5.29e+10Hz 0.0036033 -0.0134604
+ 5.3e+10Hz 0.00358404 -0.013484
+ 5.31e+10Hz 0.00356477 -0.0135075
+ 5.32e+10Hz 0.00354547 -0.013531
+ 5.33e+10Hz 0.00352615 -0.0135544
+ 5.34e+10Hz 0.00350681 -0.0135778
+ 5.35e+10Hz 0.00348745 -0.0136011
+ 5.36e+10Hz 0.00346807 -0.0136244
+ 5.37e+10Hz 0.00344867 -0.0136477
+ 5.38e+10Hz 0.00342925 -0.0136709
+ 5.39e+10Hz 0.0034098 -0.0136941
+ 5.4e+10Hz 0.00339034 -0.0137172
+ 5.41e+10Hz 0.00337085 -0.0137403
+ 5.42e+10Hz 0.00335135 -0.0137634
+ 5.43e+10Hz 0.00333182 -0.0137865
+ 5.44e+10Hz 0.00331228 -0.0138095
+ 5.45e+10Hz 0.00329271 -0.0138324
+ 5.46e+10Hz 0.00327312 -0.0138554
+ 5.47e+10Hz 0.00325351 -0.0138783
+ 5.48e+10Hz 0.00323388 -0.0139011
+ 5.49e+10Hz 0.00321423 -0.013924
+ 5.5e+10Hz 0.00319455 -0.0139468
+ 5.51e+10Hz 0.00317486 -0.0139695
+ 5.52e+10Hz 0.00315514 -0.0139923
+ 5.53e+10Hz 0.0031354 -0.014015
+ 5.54e+10Hz 0.00311564 -0.0140376
+ 5.55e+10Hz 0.00309586 -0.0140603
+ 5.56e+10Hz 0.00307606 -0.0140829
+ 5.57e+10Hz 0.00305623 -0.0141055
+ 5.58e+10Hz 0.00303638 -0.014128
+ 5.59e+10Hz 0.00301651 -0.0141505
+ 5.6e+10Hz 0.00299662 -0.014173
+ 5.61e+10Hz 0.0029767 -0.0141955
+ 5.62e+10Hz 0.00295676 -0.0142179
+ 5.63e+10Hz 0.00293679 -0.0142403
+ 5.64e+10Hz 0.0029168 -0.0142626
+ 5.65e+10Hz 0.00289679 -0.014285
+ 5.66e+10Hz 0.00287675 -0.0143073
+ 5.67e+10Hz 0.00285669 -0.0143296
+ 5.68e+10Hz 0.0028366 -0.0143518
+ 5.69e+10Hz 0.00281649 -0.014374
+ 5.7e+10Hz 0.00279635 -0.0143962
+ 5.71e+10Hz 0.00277619 -0.0144184
+ 5.72e+10Hz 0.002756 -0.0144406
+ 5.73e+10Hz 0.00273579 -0.0144627
+ 5.74e+10Hz 0.00271554 -0.0144848
+ 5.75e+10Hz 0.00269527 -0.0145068
+ 5.76e+10Hz 0.00267498 -0.0145288
+ 5.77e+10Hz 0.00265465 -0.0145509
+ 5.78e+10Hz 0.0026343 -0.0145728
+ 5.79e+10Hz 0.00261392 -0.0145948
+ 5.8e+10Hz 0.00259351 -0.0146167
+ 5.81e+10Hz 0.00257308 -0.0146386
+ 5.82e+10Hz 0.00255261 -0.0146605
+ 5.83e+10Hz 0.00253212 -0.0146823
+ 5.84e+10Hz 0.00251159 -0.0147042
+ 5.85e+10Hz 0.00249104 -0.014726
+ 5.86e+10Hz 0.00247045 -0.0147477
+ 5.87e+10Hz 0.00244984 -0.0147695
+ 5.88e+10Hz 0.00242919 -0.0147912
+ 5.89e+10Hz 0.00240851 -0.0148129
+ 5.9e+10Hz 0.00238781 -0.0148345
+ 5.91e+10Hz 0.00236707 -0.0148562
+ 5.92e+10Hz 0.00234629 -0.0148778
+ 5.93e+10Hz 0.00232549 -0.0148994
+ 5.94e+10Hz 0.00230465 -0.0149209
+ 5.95e+10Hz 0.00228378 -0.0149425
+ 5.96e+10Hz 0.00226287 -0.014964
+ 5.97e+10Hz 0.00224194 -0.0149854
+ 5.98e+10Hz 0.00222096 -0.0150069
+ 5.99e+10Hz 0.00219996 -0.0150283
+ 6e+10Hz 0.00217892 -0.0150497
+ 6.01e+10Hz 0.00215784 -0.0150711
+ 6.02e+10Hz 0.00213673 -0.0150924
+ 6.03e+10Hz 0.00211559 -0.0151137
+ 6.04e+10Hz 0.00209441 -0.015135
+ 6.05e+10Hz 0.00207319 -0.0151563
+ 6.06e+10Hz 0.00205194 -0.0151775
+ 6.07e+10Hz 0.00203065 -0.0151987
+ 6.08e+10Hz 0.00200932 -0.0152199
+ 6.09e+10Hz 0.00198796 -0.015241
+ 6.1e+10Hz 0.00196656 -0.0152621
+ 6.11e+10Hz 0.00194512 -0.0152832
+ 6.12e+10Hz 0.00192364 -0.0153043
+ 6.13e+10Hz 0.00190213 -0.0153253
+ 6.14e+10Hz 0.00188058 -0.0153463
+ 6.15e+10Hz 0.00185899 -0.0153672
+ 6.16e+10Hz 0.00183736 -0.0153882
+ 6.17e+10Hz 0.0018157 -0.0154091
+ 6.18e+10Hz 0.00179399 -0.0154299
+ 6.19e+10Hz 0.00177225 -0.0154508
+ 6.2e+10Hz 0.00175047 -0.0154716
+ 6.21e+10Hz 0.00172865 -0.0154924
+ 6.22e+10Hz 0.00170678 -0.0155131
+ 6.23e+10Hz 0.00168488 -0.0155338
+ 6.24e+10Hz 0.00166294 -0.0155545
+ 6.25e+10Hz 0.00164096 -0.0155751
+ 6.26e+10Hz 0.00161894 -0.0155957
+ 6.27e+10Hz 0.00159688 -0.0156163
+ 6.28e+10Hz 0.00157478 -0.0156368
+ 6.29e+10Hz 0.00155264 -0.0156574
+ 6.3e+10Hz 0.00153046 -0.0156778
+ 6.31e+10Hz 0.00150824 -0.0156983
+ 6.32e+10Hz 0.00148597 -0.0157187
+ 6.33e+10Hz 0.00146367 -0.015739
+ 6.34e+10Hz 0.00144133 -0.0157593
+ 6.35e+10Hz 0.00141894 -0.0157796
+ 6.36e+10Hz 0.00139652 -0.0157999
+ 6.37e+10Hz 0.00137405 -0.0158201
+ 6.38e+10Hz 0.00135155 -0.0158403
+ 6.39e+10Hz 0.001329 -0.0158604
+ 6.4e+10Hz 0.00130641 -0.0158805
+ 6.41e+10Hz 0.00128378 -0.0159006
+ 6.42e+10Hz 0.00126111 -0.0159206
+ 6.43e+10Hz 0.00123841 -0.0159406
+ 6.44e+10Hz 0.00121566 -0.0159605
+ 6.45e+10Hz 0.00119286 -0.0159804
+ 6.46e+10Hz 0.00117003 -0.0160003
+ 6.47e+10Hz 0.00114716 -0.0160201
+ 6.48e+10Hz 0.00112425 -0.0160399
+ 6.49e+10Hz 0.0011013 -0.0160596
+ 6.5e+10Hz 0.0010783 -0.0160793
+ 6.51e+10Hz 0.00105527 -0.0160989
+ 6.52e+10Hz 0.0010322 -0.0161185
+ 6.53e+10Hz 0.00100909 -0.0161381
+ 6.54e+10Hz 0.000985935 -0.0161576
+ 6.55e+10Hz 0.000962743 -0.0161771
+ 6.56e+10Hz 0.000939512 -0.0161965
+ 6.57e+10Hz 0.000916242 -0.0162159
+ 6.58e+10Hz 0.000892933 -0.0162352
+ 6.59e+10Hz 0.000869584 -0.0162545
+ 6.6e+10Hz 0.000846197 -0.0162737
+ 6.61e+10Hz 0.000822772 -0.0162929
+ 6.62e+10Hz 0.000799308 -0.0163121
+ 6.63e+10Hz 0.000775805 -0.0163312
+ 6.64e+10Hz 0.000752265 -0.0163502
+ 6.65e+10Hz 0.000728688 -0.0163693
+ 6.66e+10Hz 0.000705072 -0.0163882
+ 6.67e+10Hz 0.00068142 -0.0164071
+ 6.68e+10Hz 0.00065773 -0.016426
+ 6.69e+10Hz 0.000634004 -0.0164448
+ 6.7e+10Hz 0.000610241 -0.0164636
+ 6.71e+10Hz 0.000586442 -0.0164823
+ 6.72e+10Hz 0.000562607 -0.0165009
+ 6.73e+10Hz 0.000538736 -0.0165195
+ 6.74e+10Hz 0.00051483 -0.0165381
+ 6.75e+10Hz 0.000490889 -0.0165566
+ 6.76e+10Hz 0.000466913 -0.0165751
+ 6.77e+10Hz 0.000442902 -0.0165935
+ 6.78e+10Hz 0.000418857 -0.0166118
+ 6.79e+10Hz 0.000394778 -0.0166301
+ 6.8e+10Hz 0.000370666 -0.0166484
+ 6.81e+10Hz 0.00034652 -0.0166666
+ 6.82e+10Hz 0.000322341 -0.0166847
+ 6.83e+10Hz 0.00029813 -0.0167028
+ 6.84e+10Hz 0.000273886 -0.0167209
+ 6.85e+10Hz 0.000249611 -0.0167388
+ 6.86e+10Hz 0.000225304 -0.0167568
+ 6.87e+10Hz 0.000200965 -0.0167747
+ 6.88e+10Hz 0.000176596 -0.0167925
+ 6.89e+10Hz 0.000152196 -0.0168102
+ 6.9e+10Hz 0.000127766 -0.016828
+ 6.91e+10Hz 0.000103306 -0.0168456
+ 6.92e+10Hz 7.88161e-05 -0.0168632
+ 6.93e+10Hz 5.42975e-05 -0.0168808
+ 6.94e+10Hz 2.97502e-05 -0.0168983
+ 6.95e+10Hz 5.17445e-06 -0.0169157
+ 6.96e+10Hz -1.94293e-05 -0.0169331
+ 6.97e+10Hz -4.40606e-05 -0.0169504
+ 6.98e+10Hz -6.87192e-05 -0.0169677
+ 6.99e+10Hz -9.34047e-05 -0.0169849
+ 7e+10Hz -0.000118117 -0.0170021
+ 7.01e+10Hz -0.000142855 -0.0170192
+ 7.02e+10Hz -0.000167619 -0.0170362
+ 7.03e+10Hz -0.000192408 -0.0170532
+ 7.04e+10Hz -0.000217222 -0.0170701
+ 7.05e+10Hz -0.00024206 -0.017087
+ 7.06e+10Hz -0.000266923 -0.0171039
+ 7.07e+10Hz -0.00029181 -0.0171206
+ 7.08e+10Hz -0.00031672 -0.0171373
+ 7.09e+10Hz -0.000341654 -0.017154
+ 7.1e+10Hz -0.000366609 -0.0171706
+ 7.11e+10Hz -0.000391588 -0.0171871
+ 7.12e+10Hz -0.000416588 -0.0172036
+ 7.13e+10Hz -0.000441609 -0.01722
+ 7.14e+10Hz -0.000466652 -0.0172364
+ 7.15e+10Hz -0.000491716 -0.0172527
+ 7.16e+10Hz -0.0005168 -0.017269
+ 7.17e+10Hz -0.000541904 -0.0172852
+ 7.18e+10Hz -0.000567028 -0.0173013
+ 7.19e+10Hz -0.000592171 -0.0173174
+ 7.2e+10Hz -0.000617333 -0.0173335
+ 7.21e+10Hz -0.000642514 -0.0173494
+ 7.22e+10Hz -0.000667713 -0.0173654
+ 7.23e+10Hz -0.000692929 -0.0173812
+ 7.24e+10Hz -0.000718164 -0.017397
+ 7.25e+10Hz -0.000743415 -0.0174128
+ 7.26e+10Hz -0.000768684 -0.0174285
+ 7.27e+10Hz -0.000793969 -0.0174441
+ 7.28e+10Hz -0.00081927 -0.0174597
+ 7.29e+10Hz -0.000844587 -0.0174752
+ 7.3e+10Hz -0.000869919 -0.0174907
+ 7.31e+10Hz -0.000895267 -0.0175061
+ 7.32e+10Hz -0.000920629 -0.0175215
+ 7.33e+10Hz -0.000946006 -0.0175368
+ 7.34e+10Hz -0.000971398 -0.017552
+ 7.35e+10Hz -0.000996803 -0.0175672
+ 7.36e+10Hz -0.00102222 -0.0175824
+ 7.37e+10Hz -0.00104765 -0.0175975
+ 7.38e+10Hz -0.0010731 -0.0176125
+ 7.39e+10Hz -0.00109856 -0.0176275
+ 7.4e+10Hz -0.00112403 -0.0176424
+ 7.41e+10Hz -0.00114951 -0.0176573
+ 7.42e+10Hz -0.00117501 -0.0176721
+ 7.43e+10Hz -0.00120051 -0.0176869
+ 7.44e+10Hz -0.00122603 -0.0177016
+ 7.45e+10Hz -0.00125156 -0.0177162
+ 7.46e+10Hz -0.0012771 -0.0177308
+ 7.47e+10Hz -0.00130265 -0.0177454
+ 7.48e+10Hz -0.00132821 -0.0177599
+ 7.49e+10Hz -0.00135379 -0.0177743
+ 7.5e+10Hz -0.00137937 -0.0177887
+ 7.51e+10Hz -0.00140496 -0.0178031
+ 7.52e+10Hz -0.00143056 -0.0178174
+ 7.53e+10Hz -0.00145617 -0.0178316
+ 7.54e+10Hz -0.00148179 -0.0178458
+ 7.55e+10Hz -0.00150742 -0.0178599
+ 7.56e+10Hz -0.00153306 -0.017874
+ 7.57e+10Hz -0.00155871 -0.0178881
+ 7.58e+10Hz -0.00158436 -0.0179021
+ 7.59e+10Hz -0.00161003 -0.017916
+ 7.6e+10Hz -0.0016357 -0.0179299
+ 7.61e+10Hz -0.00166138 -0.0179437
+ 7.62e+10Hz -0.00168707 -0.0179575
+ 7.63e+10Hz -0.00171277 -0.0179712
+ 7.64e+10Hz -0.00173847 -0.0179849
+ 7.65e+10Hz -0.00176418 -0.0179986
+ 7.66e+10Hz -0.0017899 -0.0180121
+ 7.67e+10Hz -0.00181563 -0.0180257
+ 7.68e+10Hz -0.00184136 -0.0180392
+ 7.69e+10Hz -0.0018671 -0.0180526
+ 7.7e+10Hz -0.00189285 -0.018066
+ 7.71e+10Hz -0.00191861 -0.0180794
+ 7.72e+10Hz -0.00194437 -0.0180927
+ 7.73e+10Hz -0.00197014 -0.0181059
+ 7.74e+10Hz -0.00199592 -0.0181191
+ 7.75e+10Hz -0.0020217 -0.0181323
+ 7.76e+10Hz -0.00204749 -0.0181454
+ 7.77e+10Hz -0.00207328 -0.0181585
+ 7.78e+10Hz -0.00209909 -0.0181715
+ 7.79e+10Hz -0.0021249 -0.0181845
+ 7.8e+10Hz -0.00215071 -0.0181974
+ 7.81e+10Hz -0.00217654 -0.0182103
+ 7.82e+10Hz -0.00220237 -0.0182231
+ 7.83e+10Hz -0.0022282 -0.0182359
+ 7.84e+10Hz -0.00225405 -0.0182487
+ 7.85e+10Hz -0.0022799 -0.0182614
+ 7.86e+10Hz -0.00230575 -0.018274
+ 7.87e+10Hz -0.00233162 -0.0182867
+ 7.88e+10Hz -0.00235749 -0.0182992
+ 7.89e+10Hz -0.00238336 -0.0183118
+ 7.9e+10Hz -0.00240925 -0.0183242
+ 7.91e+10Hz -0.00243514 -0.0183367
+ 7.92e+10Hz -0.00246103 -0.0183491
+ 7.93e+10Hz -0.00248694 -0.0183614
+ 7.94e+10Hz -0.00251285 -0.0183737
+ 7.95e+10Hz -0.00253876 -0.018386
+ 7.96e+10Hz -0.00256469 -0.0183982
+ 7.97e+10Hz -0.00259062 -0.0184104
+ 7.98e+10Hz -0.00261656 -0.0184226
+ 7.99e+10Hz -0.00264251 -0.0184347
+ 8e+10Hz -0.00266846 -0.0184467
+ 8.01e+10Hz -0.00269442 -0.0184587
+ 8.02e+10Hz -0.00272039 -0.0184707
+ 8.03e+10Hz -0.00274637 -0.0184826
+ 8.04e+10Hz -0.00277235 -0.0184945
+ 8.05e+10Hz -0.00279834 -0.0185064
+ 8.06e+10Hz -0.00282434 -0.0185182
+ 8.07e+10Hz -0.00285035 -0.0185299
+ 8.08e+10Hz -0.00287637 -0.0185417
+ 8.09e+10Hz -0.00290239 -0.0185534
+ 8.1e+10Hz -0.00292842 -0.018565
+ 8.11e+10Hz -0.00295446 -0.0185766
+ 8.12e+10Hz -0.00298051 -0.0185882
+ 8.13e+10Hz -0.00300657 -0.0185997
+ 8.14e+10Hz -0.00303264 -0.0186111
+ 8.15e+10Hz -0.00305872 -0.0186226
+ 8.16e+10Hz -0.0030848 -0.018634
+ 8.17e+10Hz -0.00311089 -0.0186453
+ 8.18e+10Hz -0.003137 -0.0186567
+ 8.19e+10Hz -0.00316311 -0.0186679
+ 8.2e+10Hz -0.00318923 -0.0186792
+ 8.21e+10Hz -0.00321537 -0.0186904
+ 8.22e+10Hz -0.00324151 -0.0187015
+ 8.23e+10Hz -0.00326766 -0.0187126
+ 8.24e+10Hz -0.00329382 -0.0187237
+ 8.25e+10Hz -0.00332 -0.0187347
+ 8.26e+10Hz -0.00334618 -0.0187457
+ 8.27e+10Hz -0.00337237 -0.0187567
+ 8.28e+10Hz -0.00339858 -0.0187676
+ 8.29e+10Hz -0.00342479 -0.0187784
+ 8.3e+10Hz -0.00345102 -0.0187893
+ 8.31e+10Hz -0.00347725 -0.0188001
+ 8.32e+10Hz -0.0035035 -0.0188108
+ 8.33e+10Hz -0.00352976 -0.0188215
+ 8.34e+10Hz -0.00355603 -0.0188322
+ 8.35e+10Hz -0.00358231 -0.0188428
+ 8.36e+10Hz -0.00360861 -0.0188534
+ 8.37e+10Hz -0.00363491 -0.0188639
+ 8.38e+10Hz -0.00366123 -0.0188744
+ 8.39e+10Hz -0.00368756 -0.0188849
+ 8.4e+10Hz -0.0037139 -0.0188953
+ 8.41e+10Hz -0.00374026 -0.0189057
+ 8.42e+10Hz -0.00376662 -0.018916
+ 8.43e+10Hz -0.003793 -0.0189263
+ 8.44e+10Hz -0.00381939 -0.0189366
+ 8.45e+10Hz -0.0038458 -0.0189468
+ 8.46e+10Hz -0.00387221 -0.018957
+ 8.47e+10Hz -0.00389864 -0.0189671
+ 8.48e+10Hz -0.00392508 -0.0189772
+ 8.49e+10Hz -0.00395154 -0.0189872
+ 8.5e+10Hz -0.00397801 -0.0189972
+ 8.51e+10Hz -0.00400449 -0.0190072
+ 8.52e+10Hz -0.00403099 -0.0190171
+ 8.53e+10Hz -0.00405749 -0.019027
+ 8.54e+10Hz -0.00408402 -0.0190368
+ 8.55e+10Hz -0.00411055 -0.0190466
+ 8.56e+10Hz -0.0041371 -0.0190563
+ 8.57e+10Hz -0.00416367 -0.019066
+ 8.58e+10Hz -0.00419024 -0.0190757
+ 8.59e+10Hz -0.00421683 -0.0190853
+ 8.6e+10Hz -0.00424344 -0.0190948
+ 8.61e+10Hz -0.00427006 -0.0191044
+ 8.62e+10Hz -0.00429669 -0.0191138
+ 8.63e+10Hz -0.00432333 -0.0191233
+ 8.64e+10Hz -0.00435 -0.0191327
+ 8.65e+10Hz -0.00437667 -0.019142
+ 8.66e+10Hz -0.00440336 -0.0191513
+ 8.67e+10Hz -0.00443006 -0.0191606
+ 8.68e+10Hz -0.00445678 -0.0191698
+ 8.69e+10Hz -0.00448351 -0.0191789
+ 8.7e+10Hz -0.00451025 -0.0191881
+ 8.71e+10Hz -0.00453701 -0.0191971
+ 8.72e+10Hz -0.00456379 -0.0192062
+ 8.73e+10Hz -0.00459057 -0.0192151
+ 8.74e+10Hz -0.00461738 -0.0192241
+ 8.75e+10Hz -0.00464419 -0.0192329
+ 8.76e+10Hz -0.00467102 -0.0192418
+ 8.77e+10Hz -0.00469786 -0.0192506
+ 8.78e+10Hz -0.00472472 -0.0192593
+ 8.79e+10Hz -0.00475159 -0.019268
+ 8.8e+10Hz -0.00477848 -0.0192766
+ 8.81e+10Hz -0.00480538 -0.0192852
+ 8.82e+10Hz -0.00483229 -0.0192938
+ 8.83e+10Hz -0.00485922 -0.0193023
+ 8.84e+10Hz -0.00488616 -0.0193107
+ 8.85e+10Hz -0.00491311 -0.0193191
+ 8.86e+10Hz -0.00494008 -0.0193275
+ 8.87e+10Hz -0.00496706 -0.0193358
+ 8.88e+10Hz -0.00499405 -0.019344
+ 8.89e+10Hz -0.00502106 -0.0193522
+ 8.9e+10Hz -0.00504808 -0.0193604
+ 8.91e+10Hz -0.00507512 -0.0193685
+ 8.92e+10Hz -0.00510216 -0.0193765
+ 8.93e+10Hz -0.00512922 -0.0193845
+ 8.94e+10Hz -0.00515629 -0.0193925
+ 8.95e+10Hz -0.00518338 -0.0194004
+ 8.96e+10Hz -0.00521047 -0.0194082
+ 8.97e+10Hz -0.00523758 -0.019416
+ 8.98e+10Hz -0.0052647 -0.0194237
+ 8.99e+10Hz -0.00529184 -0.0194314
+ 9e+10Hz -0.00531898 -0.019439
+ 9.01e+10Hz -0.00534614 -0.0194466
+ 9.02e+10Hz -0.0053733 -0.0194541
+ 9.03e+10Hz -0.00540048 -0.0194616
+ 9.04e+10Hz -0.00542767 -0.019469
+ 9.05e+10Hz -0.00545487 -0.0194764
+ 9.06e+10Hz -0.00548208 -0.0194837
+ 9.07e+10Hz -0.00550931 -0.0194909
+ 9.08e+10Hz -0.00553654 -0.0194981
+ 9.09e+10Hz -0.00556378 -0.0195053
+ 9.1e+10Hz -0.00559103 -0.0195124
+ 9.11e+10Hz -0.00561829 -0.0195194
+ 9.12e+10Hz -0.00564557 -0.0195264
+ 9.13e+10Hz -0.00567285 -0.0195333
+ 9.14e+10Hz -0.00570014 -0.0195402
+ 9.15e+10Hz -0.00572743 -0.019547
+ 9.16e+10Hz -0.00575474 -0.0195537
+ 9.17e+10Hz -0.00578206 -0.0195604
+ 9.18e+10Hz -0.00580938 -0.0195671
+ 9.19e+10Hz -0.00583671 -0.0195737
+ 9.2e+10Hz -0.00586405 -0.0195802
+ 9.21e+10Hz -0.0058914 -0.0195867
+ 9.22e+10Hz -0.00591875 -0.0195931
+ 9.23e+10Hz -0.00594611 -0.0195994
+ 9.24e+10Hz -0.00597347 -0.0196057
+ 9.25e+10Hz -0.00600085 -0.019612
+ 9.26e+10Hz -0.00602823 -0.0196182
+ 9.27e+10Hz -0.00605561 -0.0196243
+ 9.28e+10Hz -0.006083 -0.0196304
+ 9.29e+10Hz -0.00611039 -0.0196364
+ 9.3e+10Hz -0.00613779 -0.0196423
+ 9.31e+10Hz -0.0061652 -0.0196482
+ 9.32e+10Hz -0.00619261 -0.019654
+ 9.33e+10Hz -0.00622002 -0.0196598
+ 9.34e+10Hz -0.00624744 -0.0196655
+ 9.35e+10Hz -0.00627485 -0.0196712
+ 9.36e+10Hz -0.00630228 -0.0196768
+ 9.37e+10Hz -0.0063297 -0.0196823
+ 9.38e+10Hz -0.00635713 -0.0196878
+ 9.39e+10Hz -0.00638456 -0.0196932
+ 9.4e+10Hz -0.00641199 -0.0196986
+ 9.41e+10Hz -0.00643943 -0.0197039
+ 9.42e+10Hz -0.00646686 -0.0197091
+ 9.43e+10Hz -0.0064943 -0.0197143
+ 9.44e+10Hz -0.00652173 -0.0197194
+ 9.45e+10Hz -0.00654917 -0.0197245
+ 9.46e+10Hz -0.0065766 -0.0197295
+ 9.47e+10Hz -0.00660404 -0.0197344
+ 9.48e+10Hz -0.00663148 -0.0197393
+ 9.49e+10Hz -0.00665891 -0.0197441
+ 9.5e+10Hz -0.00668634 -0.0197489
+ 9.51e+10Hz -0.00671377 -0.0197536
+ 9.52e+10Hz -0.0067412 -0.0197582
+ 9.53e+10Hz -0.00676863 -0.0197628
+ 9.54e+10Hz -0.00679605 -0.0197673
+ 9.55e+10Hz -0.00682347 -0.0197718
+ 9.56e+10Hz -0.00685089 -0.0197762
+ 9.57e+10Hz -0.00687831 -0.0197805
+ 9.58e+10Hz -0.00690572 -0.0197848
+ 9.59e+10Hz -0.00693312 -0.019789
+ 9.6e+10Hz -0.00696052 -0.0197932
+ 9.61e+10Hz -0.00698792 -0.0197973
+ 9.62e+10Hz -0.00701531 -0.0198014
+ 9.63e+10Hz -0.0070427 -0.0198053
+ 9.64e+10Hz -0.00707008 -0.0198093
+ 9.65e+10Hz -0.00709745 -0.0198131
+ 9.66e+10Hz -0.00712482 -0.0198169
+ 9.67e+10Hz -0.00715218 -0.0198207
+ 9.68e+10Hz -0.00717953 -0.0198243
+ 9.69e+10Hz -0.00720688 -0.019828
+ 9.7e+10Hz -0.00723421 -0.0198315
+ 9.71e+10Hz -0.00726154 -0.019835
+ 9.72e+10Hz -0.00728887 -0.0198385
+ 9.73e+10Hz -0.00731618 -0.0198418
+ 9.74e+10Hz -0.00734348 -0.0198452
+ 9.75e+10Hz -0.00737078 -0.0198484
+ 9.76e+10Hz -0.00739806 -0.0198516
+ 9.77e+10Hz -0.00742533 -0.0198548
+ 9.78e+10Hz -0.0074526 -0.0198579
+ 9.79e+10Hz -0.00747985 -0.0198609
+ 9.8e+10Hz -0.0075071 -0.0198639
+ 9.81e+10Hz -0.00753433 -0.0198668
+ 9.82e+10Hz -0.00756155 -0.0198696
+ 9.83e+10Hz -0.00758876 -0.0198724
+ 9.84e+10Hz -0.00761595 -0.0198752
+ 9.85e+10Hz -0.00764314 -0.0198778
+ 9.86e+10Hz -0.00767031 -0.0198805
+ 9.87e+10Hz -0.00769747 -0.019883
+ 9.88e+10Hz -0.00772461 -0.0198855
+ 9.89e+10Hz -0.00775175 -0.019888
+ 9.9e+10Hz -0.00777887 -0.0198904
+ 9.91e+10Hz -0.00780597 -0.0198927
+ 9.92e+10Hz -0.00783306 -0.019895
+ 9.93e+10Hz -0.00786014 -0.0198972
+ 9.94e+10Hz -0.0078872 -0.0198993
+ 9.95e+10Hz -0.00791425 -0.0199014
+ 9.96e+10Hz -0.00794128 -0.0199035
+ 9.97e+10Hz -0.00796829 -0.0199055
+ 9.98e+10Hz -0.0079953 -0.0199074
+ 9.99e+10Hz -0.00802228 -0.0199093
+ 1e+11Hz -0.00804925 -0.0199111
+ 1.001e+11Hz -0.0080762 -0.0199129
+ 1.002e+11Hz -0.00810314 -0.0199146
+ 1.003e+11Hz -0.00813006 -0.0199162
+ 1.004e+11Hz -0.00815696 -0.0199178
+ 1.005e+11Hz -0.00818384 -0.0199194
+ 1.006e+11Hz -0.00821071 -0.0199209
+ 1.007e+11Hz -0.00823756 -0.0199223
+ 1.008e+11Hz -0.00826439 -0.0199237
+ 1.009e+11Hz -0.00829121 -0.019925
+ 1.01e+11Hz -0.008318 -0.0199263
+ 1.011e+11Hz -0.00834478 -0.0199275
+ 1.012e+11Hz -0.00837154 -0.0199287
+ 1.013e+11Hz -0.00839828 -0.0199298
+ 1.014e+11Hz -0.008425 -0.0199309
+ 1.015e+11Hz -0.0084517 -0.0199319
+ 1.016e+11Hz -0.00847838 -0.0199328
+ 1.017e+11Hz -0.00850504 -0.0199337
+ 1.018e+11Hz -0.00853169 -0.0199346
+ 1.019e+11Hz -0.00855831 -0.0199354
+ 1.02e+11Hz -0.00858491 -0.0199361
+ 1.021e+11Hz -0.0086115 -0.0199368
+ 1.022e+11Hz -0.00863806 -0.0199374
+ 1.023e+11Hz -0.0086646 -0.019938
+ 1.024e+11Hz -0.00869113 -0.0199386
+ 1.025e+11Hz -0.00871763 -0.019939
+ 1.026e+11Hz -0.00874411 -0.0199395
+ 1.027e+11Hz -0.00877057 -0.0199399
+ 1.028e+11Hz -0.00879701 -0.0199402
+ 1.029e+11Hz -0.00882343 -0.0199405
+ 1.03e+11Hz -0.00884982 -0.0199407
+ 1.031e+11Hz -0.0088762 -0.0199409
+ 1.032e+11Hz -0.00890255 -0.019941
+ 1.033e+11Hz -0.00892888 -0.0199411
+ 1.034e+11Hz -0.00895519 -0.0199412
+ 1.035e+11Hz -0.00898148 -0.0199412
+ 1.036e+11Hz -0.00900775 -0.0199411
+ 1.037e+11Hz -0.00903399 -0.019941
+ 1.038e+11Hz -0.00906022 -0.0199408
+ 1.039e+11Hz -0.00908642 -0.0199406
+ 1.04e+11Hz -0.0091126 -0.0199404
+ 1.041e+11Hz -0.00913875 -0.0199401
+ 1.042e+11Hz -0.00916489 -0.0199397
+ 1.043e+11Hz -0.009191 -0.0199393
+ 1.044e+11Hz -0.00921709 -0.0199389
+ 1.045e+11Hz -0.00924315 -0.0199384
+ 1.046e+11Hz -0.0092692 -0.0199378
+ 1.047e+11Hz -0.00929522 -0.0199373
+ 1.048e+11Hz -0.00932122 -0.0199366
+ 1.049e+11Hz -0.00934719 -0.0199359
+ 1.05e+11Hz -0.00937315 -0.0199352
+ 1.051e+11Hz -0.00939908 -0.0199345
+ 1.052e+11Hz -0.00942498 -0.0199336
+ 1.053e+11Hz -0.00945087 -0.0199328
+ 1.054e+11Hz -0.00947673 -0.0199319
+ 1.055e+11Hz -0.00950257 -0.0199309
+ 1.056e+11Hz -0.00952838 -0.0199299
+ 1.057e+11Hz -0.00955417 -0.0199289
+ 1.058e+11Hz -0.00957994 -0.0199278
+ 1.059e+11Hz -0.00960569 -0.0199267
+ 1.06e+11Hz -0.00963141 -0.0199255
+ 1.061e+11Hz -0.00965711 -0.0199243
+ 1.062e+11Hz -0.00968279 -0.019923
+ 1.063e+11Hz -0.00970844 -0.0199217
+ 1.064e+11Hz -0.00973407 -0.0199203
+ 1.065e+11Hz -0.00975968 -0.0199189
+ 1.066e+11Hz -0.00978526 -0.0199175
+ 1.067e+11Hz -0.00981082 -0.019916
+ 1.068e+11Hz -0.00983636 -0.0199145
+ 1.069e+11Hz -0.00986187 -0.0199129
+ 1.07e+11Hz -0.00988736 -0.0199113
+ 1.071e+11Hz -0.00991283 -0.0199096
+ 1.072e+11Hz -0.00993828 -0.019908
+ 1.073e+11Hz -0.0099637 -0.0199062
+ 1.074e+11Hz -0.00998909 -0.0199044
+ 1.075e+11Hz -0.0100145 -0.0199026
+ 1.076e+11Hz -0.0100398 -0.0199007
+ 1.077e+11Hz -0.0100651 -0.0198988
+ 1.078e+11Hz -0.0100905 -0.0198969
+ 1.079e+11Hz -0.0101157 -0.0198949
+ 1.08e+11Hz -0.010141 -0.0198928
+ 1.081e+11Hz -0.0101662 -0.0198908
+ 1.082e+11Hz -0.0101914 -0.0198886
+ 1.083e+11Hz -0.0102166 -0.0198865
+ 1.084e+11Hz -0.0102418 -0.0198843
+ 1.085e+11Hz -0.0102669 -0.019882
+ 1.086e+11Hz -0.0102921 -0.0198797
+ 1.087e+11Hz -0.0103172 -0.0198774
+ 1.088e+11Hz -0.0103422 -0.019875
+ 1.089e+11Hz -0.0103673 -0.0198726
+ 1.09e+11Hz -0.0103923 -0.0198702
+ 1.091e+11Hz -0.0104173 -0.0198677
+ 1.092e+11Hz -0.0104423 -0.0198652
+ 1.093e+11Hz -0.0104672 -0.0198626
+ 1.094e+11Hz -0.0104922 -0.01986
+ 1.095e+11Hz -0.0105171 -0.0198573
+ 1.096e+11Hz -0.010542 -0.0198546
+ 1.097e+11Hz -0.0105668 -0.0198519
+ 1.098e+11Hz -0.0105917 -0.0198491
+ 1.099e+11Hz -0.0106165 -0.0198463
+ 1.1e+11Hz -0.0106413 -0.0198434
+ 1.101e+11Hz -0.0106661 -0.0198405
+ 1.102e+11Hz -0.0106908 -0.0198376
+ 1.103e+11Hz -0.0107155 -0.0198346
+ 1.104e+11Hz -0.0107403 -0.0198316
+ 1.105e+11Hz -0.0107649 -0.0198285
+ 1.106e+11Hz -0.0107896 -0.0198254
+ 1.107e+11Hz -0.0108142 -0.0198223
+ 1.108e+11Hz -0.0108388 -0.0198191
+ 1.109e+11Hz -0.0108634 -0.0198159
+ 1.11e+11Hz -0.010888 -0.0198126
+ 1.111e+11Hz -0.0109125 -0.0198093
+ 1.112e+11Hz -0.010937 -0.019806
+ 1.113e+11Hz -0.0109615 -0.0198026
+ 1.114e+11Hz -0.010986 -0.0197992
+ 1.115e+11Hz -0.0110105 -0.0197957
+ 1.116e+11Hz -0.0110349 -0.0197922
+ 1.117e+11Hz -0.0110593 -0.0197887
+ 1.118e+11Hz -0.0110837 -0.0197851
+ 1.119e+11Hz -0.011108 -0.0197815
+ 1.12e+11Hz -0.0111324 -0.0197778
+ 1.121e+11Hz -0.0111567 -0.0197741
+ 1.122e+11Hz -0.011181 -0.0197704
+ 1.123e+11Hz -0.0112052 -0.0197666
+ 1.124e+11Hz -0.0112295 -0.0197628
+ 1.125e+11Hz -0.0112537 -0.0197589
+ 1.126e+11Hz -0.0112779 -0.019755
+ 1.127e+11Hz -0.011302 -0.0197511
+ 1.128e+11Hz -0.0113262 -0.0197471
+ 1.129e+11Hz -0.0113503 -0.0197431
+ 1.13e+11Hz -0.0113744 -0.019739
+ 1.131e+11Hz -0.0113985 -0.0197349
+ 1.132e+11Hz -0.0114225 -0.0197308
+ 1.133e+11Hz -0.0114466 -0.0197266
+ 1.134e+11Hz -0.0114706 -0.0197224
+ 1.135e+11Hz -0.0114945 -0.0197181
+ 1.136e+11Hz -0.0115185 -0.0197138
+ 1.137e+11Hz -0.0115424 -0.0197095
+ 1.138e+11Hz -0.0115663 -0.0197051
+ 1.139e+11Hz -0.0115902 -0.0197007
+ 1.14e+11Hz -0.0116141 -0.0196962
+ 1.141e+11Hz -0.0116379 -0.0196917
+ 1.142e+11Hz -0.0116617 -0.0196872
+ 1.143e+11Hz -0.0116855 -0.0196826
+ 1.144e+11Hz -0.0117093 -0.019678
+ 1.145e+11Hz -0.011733 -0.0196733
+ 1.146e+11Hz -0.0117567 -0.0196686
+ 1.147e+11Hz -0.0117804 -0.0196638
+ 1.148e+11Hz -0.0118041 -0.0196591
+ 1.149e+11Hz -0.0118277 -0.0196542
+ 1.15e+11Hz -0.0118513 -0.0196494
+ 1.151e+11Hz -0.0118749 -0.0196445
+ 1.152e+11Hz -0.0118985 -0.0196395
+ 1.153e+11Hz -0.011922 -0.0196345
+ 1.154e+11Hz -0.0119455 -0.0196295
+ 1.155e+11Hz -0.011969 -0.0196245
+ 1.156e+11Hz -0.0119925 -0.0196194
+ 1.157e+11Hz -0.0120159 -0.0196142
+ 1.158e+11Hz -0.0120393 -0.019609
+ 1.159e+11Hz -0.0120627 -0.0196038
+ 1.16e+11Hz -0.012086 -0.0195985
+ 1.161e+11Hz -0.0121094 -0.0195932
+ 1.162e+11Hz -0.0121327 -0.0195879
+ 1.163e+11Hz -0.0121559 -0.0195825
+ 1.164e+11Hz -0.0121792 -0.019577
+ 1.165e+11Hz -0.0122024 -0.0195716
+ 1.166e+11Hz -0.0122256 -0.0195661
+ 1.167e+11Hz -0.0122488 -0.0195605
+ 1.168e+11Hz -0.0122719 -0.0195549
+ 1.169e+11Hz -0.012295 -0.0195493
+ 1.17e+11Hz -0.0123181 -0.0195436
+ 1.171e+11Hz -0.0123412 -0.0195379
+ 1.172e+11Hz -0.0123642 -0.0195322
+ 1.173e+11Hz -0.0123872 -0.0195264
+ 1.174e+11Hz -0.0124102 -0.0195205
+ 1.175e+11Hz -0.0124331 -0.0195147
+ 1.176e+11Hz -0.012456 -0.0195087
+ 1.177e+11Hz -0.0124789 -0.0195028
+ 1.178e+11Hz -0.0125018 -0.0194968
+ 1.179e+11Hz -0.0125246 -0.0194908
+ 1.18e+11Hz -0.0125474 -0.0194847
+ 1.181e+11Hz -0.0125702 -0.0194786
+ 1.182e+11Hz -0.0125929 -0.0194724
+ 1.183e+11Hz -0.0126157 -0.0194662
+ 1.184e+11Hz -0.0126383 -0.01946
+ 1.185e+11Hz -0.012661 -0.0194537
+ 1.186e+11Hz -0.0126836 -0.0194474
+ 1.187e+11Hz -0.0127062 -0.019441
+ 1.188e+11Hz -0.0127288 -0.0194346
+ 1.189e+11Hz -0.0127513 -0.0194282
+ 1.19e+11Hz -0.0127738 -0.0194217
+ 1.191e+11Hz -0.0127963 -0.0194152
+ 1.192e+11Hz -0.0128187 -0.0194086
+ 1.193e+11Hz -0.0128411 -0.019402
+ 1.194e+11Hz -0.0128635 -0.0193954
+ 1.195e+11Hz -0.0128859 -0.0193887
+ 1.196e+11Hz -0.0129082 -0.019382
+ 1.197e+11Hz -0.0129304 -0.0193752
+ 1.198e+11Hz -0.0129527 -0.0193684
+ 1.199e+11Hz -0.0129749 -0.0193616
+ 1.2e+11Hz -0.0129971 -0.0193547
+ 1.201e+11Hz -0.0130192 -0.0193478
+ 1.202e+11Hz -0.0130414 -0.0193409
+ 1.203e+11Hz -0.0130635 -0.0193339
+ 1.204e+11Hz -0.0130855 -0.0193268
+ 1.205e+11Hz -0.0131075 -0.0193198
+ 1.206e+11Hz -0.0131295 -0.0193126
+ 1.207e+11Hz -0.0131515 -0.0193055
+ 1.208e+11Hz -0.0131734 -0.0192983
+ 1.209e+11Hz -0.0131953 -0.0192911
+ 1.21e+11Hz -0.0132171 -0.0192838
+ 1.211e+11Hz -0.0132389 -0.0192765
+ 1.212e+11Hz -0.0132607 -0.0192692
+ 1.213e+11Hz -0.0132824 -0.0192618
+ 1.214e+11Hz -0.0133041 -0.0192544
+ 1.215e+11Hz -0.0133258 -0.0192469
+ 1.216e+11Hz -0.0133475 -0.0192394
+ 1.217e+11Hz -0.0133691 -0.0192319
+ 1.218e+11Hz -0.0133906 -0.0192243
+ 1.219e+11Hz -0.0134122 -0.0192167
+ 1.22e+11Hz -0.0134336 -0.019209
+ 1.221e+11Hz -0.0134551 -0.0192013
+ 1.222e+11Hz -0.0134765 -0.0191936
+ 1.223e+11Hz -0.0134979 -0.0191859
+ 1.224e+11Hz -0.0135192 -0.0191781
+ 1.225e+11Hz -0.0135405 -0.0191702
+ 1.226e+11Hz -0.0135618 -0.0191624
+ 1.227e+11Hz -0.013583 -0.0191544
+ 1.228e+11Hz -0.0136042 -0.0191465
+ 1.229e+11Hz -0.0136254 -0.0191385
+ 1.23e+11Hz -0.0136465 -0.0191305
+ 1.231e+11Hz -0.0136676 -0.0191225
+ 1.232e+11Hz -0.0136886 -0.0191144
+ 1.233e+11Hz -0.0137096 -0.0191062
+ 1.234e+11Hz -0.0137306 -0.0190981
+ 1.235e+11Hz -0.0137515 -0.0190899
+ 1.236e+11Hz -0.0137724 -0.0190816
+ 1.237e+11Hz -0.0137932 -0.0190734
+ 1.238e+11Hz -0.013814 -0.0190651
+ 1.239e+11Hz -0.0138348 -0.0190567
+ 1.24e+11Hz -0.0138555 -0.0190484
+ 1.241e+11Hz -0.0138762 -0.01904
+ 1.242e+11Hz -0.0138969 -0.0190315
+ 1.243e+11Hz -0.0139175 -0.019023
+ 1.244e+11Hz -0.013938 -0.0190145
+ 1.245e+11Hz -0.0139585 -0.019006
+ 1.246e+11Hz -0.013979 -0.0189974
+ 1.247e+11Hz -0.0139995 -0.0189888
+ 1.248e+11Hz -0.0140199 -0.0189802
+ 1.249e+11Hz -0.0140402 -0.0189715
+ 1.25e+11Hz -0.0140605 -0.0189628
+ 1.251e+11Hz -0.0140808 -0.018954
+ 1.252e+11Hz -0.014101 -0.0189452
+ 1.253e+11Hz -0.0141212 -0.0189364
+ 1.254e+11Hz -0.0141414 -0.0189276
+ 1.255e+11Hz -0.0141615 -0.0189187
+ 1.256e+11Hz -0.0141815 -0.0189098
+ 1.257e+11Hz -0.0142015 -0.0189009
+ 1.258e+11Hz -0.0142215 -0.0188919
+ 1.259e+11Hz -0.0142414 -0.0188829
+ 1.26e+11Hz -0.0142613 -0.0188739
+ 1.261e+11Hz -0.0142812 -0.0188648
+ 1.262e+11Hz -0.014301 -0.0188557
+ 1.263e+11Hz -0.0143207 -0.0188466
+ 1.264e+11Hz -0.0143404 -0.0188375
+ 1.265e+11Hz -0.0143601 -0.0188283
+ 1.266e+11Hz -0.0143797 -0.0188191
+ 1.267e+11Hz -0.0143993 -0.0188098
+ 1.268e+11Hz -0.0144188 -0.0188006
+ 1.269e+11Hz -0.0144383 -0.0187913
+ 1.27e+11Hz -0.0144578 -0.018782
+ 1.271e+11Hz -0.0144772 -0.0187726
+ 1.272e+11Hz -0.0144965 -0.0187632
+ 1.273e+11Hz -0.0145159 -0.0187538
+ 1.274e+11Hz -0.0145351 -0.0187444
+ 1.275e+11Hz -0.0145543 -0.0187349
+ 1.276e+11Hz -0.0145735 -0.0187254
+ 1.277e+11Hz -0.0145926 -0.0187159
+ 1.278e+11Hz -0.0146117 -0.0187063
+ 1.279e+11Hz -0.0146308 -0.0186968
+ 1.28e+11Hz -0.0146498 -0.0186872
+ 1.281e+11Hz -0.0146687 -0.0186775
+ 1.282e+11Hz -0.0146876 -0.0186679
+ 1.283e+11Hz -0.0147065 -0.0186582
+ 1.284e+11Hz -0.0147253 -0.0186485
+ 1.285e+11Hz -0.0147441 -0.0186388
+ 1.286e+11Hz -0.0147628 -0.018629
+ 1.287e+11Hz -0.0147814 -0.0186192
+ 1.288e+11Hz -0.0148001 -0.0186094
+ 1.289e+11Hz -0.0148186 -0.0185996
+ 1.29e+11Hz -0.0148372 -0.0185897
+ 1.291e+11Hz -0.0148557 -0.0185799
+ 1.292e+11Hz -0.0148741 -0.01857
+ 1.293e+11Hz -0.0148925 -0.01856
+ 1.294e+11Hz -0.0149108 -0.0185501
+ 1.295e+11Hz -0.0149291 -0.0185401
+ 1.296e+11Hz -0.0149474 -0.0185301
+ 1.297e+11Hz -0.0149656 -0.0185201
+ 1.298e+11Hz -0.0149838 -0.0185101
+ 1.299e+11Hz -0.0150019 -0.0185
+ 1.3e+11Hz -0.0150199 -0.0184899
+ 1.301e+11Hz -0.0150379 -0.0184798
+ 1.302e+11Hz -0.0150559 -0.0184697
+ 1.303e+11Hz -0.0150738 -0.0184595
+ 1.304e+11Hz -0.0150917 -0.0184494
+ 1.305e+11Hz -0.0151095 -0.0184392
+ 1.306e+11Hz -0.0151273 -0.018429
+ 1.307e+11Hz -0.015145 -0.0184187
+ 1.308e+11Hz -0.0151627 -0.0184085
+ 1.309e+11Hz -0.0151804 -0.0183982
+ 1.31e+11Hz -0.0151979 -0.0183879
+ 1.311e+11Hz -0.0152155 -0.0183776
+ 1.312e+11Hz -0.015233 -0.0183673
+ 1.313e+11Hz -0.0152504 -0.018357
+ 1.314e+11Hz -0.0152678 -0.0183466
+ 1.315e+11Hz -0.0152852 -0.0183362
+ 1.316e+11Hz -0.0153025 -0.0183258
+ 1.317e+11Hz -0.0153197 -0.0183154
+ 1.318e+11Hz -0.0153369 -0.018305
+ 1.319e+11Hz -0.0153541 -0.0182945
+ 1.32e+11Hz -0.0153712 -0.018284
+ 1.321e+11Hz -0.0153883 -0.0182735
+ 1.322e+11Hz -0.0154053 -0.018263
+ 1.323e+11Hz -0.0154222 -0.0182525
+ 1.324e+11Hz -0.0154392 -0.018242
+ 1.325e+11Hz -0.015456 -0.0182314
+ 1.326e+11Hz -0.0154729 -0.0182209
+ 1.327e+11Hz -0.0154896 -0.0182103
+ 1.328e+11Hz -0.0155064 -0.0181997
+ 1.329e+11Hz -0.015523 -0.0181891
+ 1.33e+11Hz -0.0155397 -0.0181784
+ 1.331e+11Hz -0.0155562 -0.0181678
+ 1.332e+11Hz -0.0155728 -0.0181571
+ 1.333e+11Hz -0.0155893 -0.0181464
+ 1.334e+11Hz -0.0156057 -0.0181358
+ 1.335e+11Hz -0.0156221 -0.0181251
+ 1.336e+11Hz -0.0156384 -0.0181143
+ 1.337e+11Hz -0.0156547 -0.0181036
+ 1.338e+11Hz -0.015671 -0.0180929
+ 1.339e+11Hz -0.0156872 -0.0180821
+ 1.34e+11Hz -0.0157033 -0.0180714
+ 1.341e+11Hz -0.0157194 -0.0180606
+ 1.342e+11Hz -0.0157355 -0.0180498
+ 1.343e+11Hz -0.0157515 -0.018039
+ 1.344e+11Hz -0.0157674 -0.0180282
+ 1.345e+11Hz -0.0157833 -0.0180173
+ 1.346e+11Hz -0.0157992 -0.0180065
+ 1.347e+11Hz -0.015815 -0.0179956
+ 1.348e+11Hz -0.0158308 -0.0179848
+ 1.349e+11Hz -0.0158465 -0.0179739
+ 1.35e+11Hz -0.0158622 -0.017963
+ 1.351e+11Hz -0.0158778 -0.0179521
+ 1.352e+11Hz -0.0158933 -0.0179412
+ 1.353e+11Hz -0.0159089 -0.0179303
+ 1.354e+11Hz -0.0159243 -0.0179194
+ 1.355e+11Hz -0.0159398 -0.0179084
+ 1.356e+11Hz -0.0159552 -0.0178975
+ 1.357e+11Hz -0.0159705 -0.0178865
+ 1.358e+11Hz -0.0159858 -0.0178756
+ 1.359e+11Hz -0.016001 -0.0178646
+ 1.36e+11Hz -0.0160162 -0.0178536
+ 1.361e+11Hz -0.0160313 -0.0178426
+ 1.362e+11Hz -0.0160464 -0.0178316
+ 1.363e+11Hz -0.0160615 -0.0178206
+ 1.364e+11Hz -0.0160765 -0.0178096
+ 1.365e+11Hz -0.0160914 -0.0177986
+ 1.366e+11Hz -0.0161063 -0.0177876
+ 1.367e+11Hz -0.0161212 -0.0177765
+ 1.368e+11Hz -0.016136 -0.0177655
+ 1.369e+11Hz -0.0161507 -0.0177544
+ 1.37e+11Hz -0.0161654 -0.0177434
+ 1.371e+11Hz -0.0161801 -0.0177323
+ 1.372e+11Hz -0.0161947 -0.0177212
+ 1.373e+11Hz -0.0162093 -0.0177101
+ 1.374e+11Hz -0.0162238 -0.0176991
+ 1.375e+11Hz -0.0162383 -0.017688
+ 1.376e+11Hz -0.0162527 -0.0176769
+ 1.377e+11Hz -0.0162671 -0.0176658
+ 1.378e+11Hz -0.0162814 -0.0176547
+ 1.379e+11Hz -0.0162957 -0.0176436
+ 1.38e+11Hz -0.0163099 -0.0176324
+ 1.381e+11Hz -0.0163241 -0.0176213
+ 1.382e+11Hz -0.0163382 -0.0176102
+ 1.383e+11Hz -0.0163523 -0.0175991
+ 1.384e+11Hz -0.0163663 -0.0175879
+ 1.385e+11Hz -0.0163803 -0.0175768
+ 1.386e+11Hz -0.0163943 -0.0175656
+ 1.387e+11Hz -0.0164082 -0.0175545
+ 1.388e+11Hz -0.016422 -0.0175433
+ 1.389e+11Hz -0.0164358 -0.0175322
+ 1.39e+11Hz -0.0164495 -0.017521
+ 1.391e+11Hz -0.0164633 -0.0175099
+ 1.392e+11Hz -0.0164769 -0.0174987
+ 1.393e+11Hz -0.0164905 -0.0174875
+ 1.394e+11Hz -0.0165041 -0.0174764
+ 1.395e+11Hz -0.0165176 -0.0174652
+ 1.396e+11Hz -0.016531 -0.017454
+ 1.397e+11Hz -0.0165445 -0.0174429
+ 1.398e+11Hz -0.0165578 -0.0174317
+ 1.399e+11Hz -0.0165711 -0.0174205
+ 1.4e+11Hz -0.0165844 -0.0174093
+ 1.401e+11Hz -0.0165976 -0.0173981
+ 1.402e+11Hz -0.0166108 -0.017387
+ 1.403e+11Hz -0.0166239 -0.0173758
+ 1.404e+11Hz -0.016637 -0.0173646
+ 1.405e+11Hz -0.0166501 -0.0173534
+ 1.406e+11Hz -0.016663 -0.0173422
+ 1.407e+11Hz -0.016676 -0.017331
+ 1.408e+11Hz -0.0166889 -0.0173199
+ 1.409e+11Hz -0.0167017 -0.0173087
+ 1.41e+11Hz -0.0167145 -0.0172975
+ 1.411e+11Hz -0.0167272 -0.0172863
+ 1.412e+11Hz -0.0167399 -0.0172751
+ 1.413e+11Hz -0.0167526 -0.017264
+ 1.414e+11Hz -0.0167652 -0.0172528
+ 1.415e+11Hz -0.0167777 -0.0172416
+ 1.416e+11Hz -0.0167902 -0.0172304
+ 1.417e+11Hz -0.0168027 -0.0172193
+ 1.418e+11Hz -0.0168151 -0.0172081
+ 1.419e+11Hz -0.0168274 -0.0171969
+ 1.42e+11Hz -0.0168398 -0.0171858
+ 1.421e+11Hz -0.016852 -0.0171746
+ 1.422e+11Hz -0.0168642 -0.0171634
+ 1.423e+11Hz -0.0168764 -0.0171523
+ 1.424e+11Hz -0.0168885 -0.0171411
+ 1.425e+11Hz -0.0169006 -0.01713
+ 1.426e+11Hz -0.0169126 -0.0171189
+ 1.427e+11Hz -0.0169246 -0.0171077
+ 1.428e+11Hz -0.0169365 -0.0170966
+ 1.429e+11Hz -0.0169484 -0.0170855
+ 1.43e+11Hz -0.0169602 -0.0170743
+ 1.431e+11Hz -0.016972 -0.0170632
+ 1.432e+11Hz -0.0169837 -0.0170521
+ 1.433e+11Hz -0.0169954 -0.017041
+ 1.434e+11Hz -0.017007 -0.0170299
+ 1.435e+11Hz -0.0170186 -0.0170188
+ 1.436e+11Hz -0.0170301 -0.0170077
+ 1.437e+11Hz -0.0170416 -0.0169966
+ 1.438e+11Hz -0.017053 -0.0169856
+ 1.439e+11Hz -0.0170644 -0.0169745
+ 1.44e+11Hz -0.0170757 -0.0169634
+ 1.441e+11Hz -0.017087 -0.0169524
+ 1.442e+11Hz -0.0170983 -0.0169413
+ 1.443e+11Hz -0.0171094 -0.0169303
+ 1.444e+11Hz -0.0171206 -0.0169193
+ 1.445e+11Hz -0.0171317 -0.0169083
+ 1.446e+11Hz -0.0171427 -0.0168973
+ 1.447e+11Hz -0.0171537 -0.0168863
+ 1.448e+11Hz -0.0171646 -0.0168753
+ 1.449e+11Hz -0.0171755 -0.0168643
+ 1.45e+11Hz -0.0171864 -0.0168533
+ 1.451e+11Hz -0.0171972 -0.0168424
+ 1.452e+11Hz -0.0172079 -0.0168314
+ 1.453e+11Hz -0.0172186 -0.0168205
+ 1.454e+11Hz -0.0172293 -0.0168096
+ 1.455e+11Hz -0.0172399 -0.0167987
+ 1.456e+11Hz -0.0172504 -0.0167878
+ 1.457e+11Hz -0.0172609 -0.0167769
+ 1.458e+11Hz -0.0172714 -0.016766
+ 1.459e+11Hz -0.0172818 -0.0167551
+ 1.46e+11Hz -0.0172921 -0.0167443
+ 1.461e+11Hz -0.0173024 -0.0167335
+ 1.462e+11Hz -0.0173127 -0.0167227
+ 1.463e+11Hz -0.0173229 -0.0167119
+ 1.464e+11Hz -0.017333 -0.0167011
+ 1.465e+11Hz -0.0173432 -0.0166903
+ 1.466e+11Hz -0.0173532 -0.0166795
+ 1.467e+11Hz -0.0173632 -0.0166688
+ 1.468e+11Hz -0.0173732 -0.0166581
+ 1.469e+11Hz -0.0173831 -0.0166474
+ 1.47e+11Hz -0.017393 -0.0166367
+ 1.471e+11Hz -0.0174028 -0.016626
+ 1.472e+11Hz -0.0174125 -0.0166154
+ 1.473e+11Hz -0.0174222 -0.0166047
+ 1.474e+11Hz -0.0174319 -0.0165941
+ 1.475e+11Hz -0.0174415 -0.0165835
+ 1.476e+11Hz -0.0174511 -0.0165729
+ 1.477e+11Hz -0.0174606 -0.0165624
+ 1.478e+11Hz -0.0174701 -0.0165518
+ 1.479e+11Hz -0.0174795 -0.0165413
+ 1.48e+11Hz -0.0174889 -0.0165308
+ 1.481e+11Hz -0.0174982 -0.0165203
+ 1.482e+11Hz -0.0175074 -0.0165099
+ 1.483e+11Hz -0.0175167 -0.0164994
+ 1.484e+11Hz -0.0175258 -0.016489
+ 1.485e+11Hz -0.017535 -0.0164787
+ 1.486e+11Hz -0.0175441 -0.0164683
+ 1.487e+11Hz -0.0175531 -0.0164579
+ 1.488e+11Hz -0.0175621 -0.0164476
+ 1.489e+11Hz -0.017571 -0.0164373
+ 1.49e+11Hz -0.0175799 -0.0164271
+ 1.491e+11Hz -0.0175887 -0.0164168
+ 1.492e+11Hz -0.0175975 -0.0164066
+ 1.493e+11Hz -0.0176063 -0.0163964
+ 1.494e+11Hz -0.0176149 -0.0163863
+ 1.495e+11Hz -0.0176236 -0.0163762
+ 1.496e+11Hz -0.0176322 -0.016366
+ 1.497e+11Hz -0.0176407 -0.016356
+ 1.498e+11Hz -0.0176492 -0.0163459
+ 1.499e+11Hz -0.0176577 -0.0163359
+ 1.5e+11Hz -0.0176661 -0.0163259
+ 1.501e+11Hz -0.0176745 -0.016316
+ 1.502e+11Hz -0.0176828 -0.016306
+ 1.503e+11Hz -0.0176911 -0.0162961
+ 1.504e+11Hz -0.0176993 -0.0162863
+ 1.505e+11Hz -0.0177075 -0.0162764
+ 1.506e+11Hz -0.0177156 -0.0162666
+ 1.507e+11Hz -0.0177237 -0.0162569
+ 1.508e+11Hz -0.0177317 -0.0162471
+ 1.509e+11Hz -0.0177397 -0.0162374
+ 1.51e+11Hz -0.0177477 -0.0162278
+ 1.511e+11Hz -0.0177556 -0.0162181
+ 1.512e+11Hz -0.0177634 -0.0162085
+ 1.513e+11Hz -0.0177713 -0.016199
+ 1.514e+11Hz -0.017779 -0.0161895
+ 1.515e+11Hz -0.0177868 -0.01618
+ 1.516e+11Hz -0.0177944 -0.0161705
+ 1.517e+11Hz -0.0178021 -0.0161611
+ 1.518e+11Hz -0.0178097 -0.0161518
+ 1.519e+11Hz -0.0178172 -0.0161424
+ 1.52e+11Hz -0.0178247 -0.0161331
+ 1.521e+11Hz -0.0178322 -0.0161239
+ 1.522e+11Hz -0.0178396 -0.0161147
+ 1.523e+11Hz -0.017847 -0.0161055
+ 1.524e+11Hz -0.0178544 -0.0160964
+ 1.525e+11Hz -0.0178617 -0.0160873
+ 1.526e+11Hz -0.0178689 -0.0160782
+ 1.527e+11Hz -0.0178762 -0.0160692
+ 1.528e+11Hz -0.0178833 -0.0160603
+ 1.529e+11Hz -0.0178905 -0.0160513
+ 1.53e+11Hz -0.0178976 -0.0160425
+ 1.531e+11Hz -0.0179046 -0.0160336
+ 1.532e+11Hz -0.0179117 -0.0160249
+ 1.533e+11Hz -0.0179187 -0.0160161
+ 1.534e+11Hz -0.0179256 -0.0160074
+ 1.535e+11Hz -0.0179325 -0.0159988
+ 1.536e+11Hz -0.0179394 -0.0159902
+ 1.537e+11Hz -0.0179462 -0.0159817
+ 1.538e+11Hz -0.017953 -0.0159732
+ 1.539e+11Hz -0.0179598 -0.0159647
+ 1.54e+11Hz -0.0179665 -0.0159563
+ 1.541e+11Hz -0.0179732 -0.015948
+ 1.542e+11Hz -0.0179799 -0.0159397
+ 1.543e+11Hz -0.0179865 -0.0159314
+ 1.544e+11Hz -0.0179931 -0.0159232
+ 1.545e+11Hz -0.0179996 -0.0159151
+ 1.546e+11Hz -0.0180062 -0.015907
+ 1.547e+11Hz -0.0180126 -0.0158989
+ 1.548e+11Hz -0.0180191 -0.0158909
+ 1.549e+11Hz -0.0180255 -0.015883
+ 1.55e+11Hz -0.0180319 -0.0158751
+ 1.551e+11Hz -0.0180383 -0.0158673
+ 1.552e+11Hz -0.0180446 -0.0158595
+ 1.553e+11Hz -0.0180509 -0.0158518
+ 1.554e+11Hz -0.0180572 -0.0158442
+ 1.555e+11Hz -0.0180635 -0.0158366
+ 1.556e+11Hz -0.0180697 -0.015829
+ 1.557e+11Hz -0.0180759 -0.0158215
+ 1.558e+11Hz -0.0180821 -0.0158141
+ 1.559e+11Hz -0.0180882 -0.0158067
+ 1.56e+11Hz -0.0180943 -0.0157994
+ 1.561e+11Hz -0.0181004 -0.0157922
+ 1.562e+11Hz -0.0181065 -0.015785
+ 1.563e+11Hz -0.0181126 -0.0157779
+ 1.564e+11Hz -0.0181186 -0.0157708
+ 1.565e+11Hz -0.0181246 -0.0157638
+ 1.566e+11Hz -0.0181306 -0.0157568
+ 1.567e+11Hz -0.0181365 -0.0157499
+ 1.568e+11Hz -0.0181425 -0.0157431
+ 1.569e+11Hz -0.0181484 -0.0157364
+ 1.57e+11Hz -0.0181543 -0.0157297
+ 1.571e+11Hz -0.0181602 -0.015723
+ 1.572e+11Hz -0.0181661 -0.0157164
+ 1.573e+11Hz -0.0181719 -0.0157099
+ 1.574e+11Hz -0.0181778 -0.0157035
+ 1.575e+11Hz -0.0181836 -0.0156971
+ 1.576e+11Hz -0.0181894 -0.0156908
+ 1.577e+11Hz -0.0181952 -0.0156845
+ 1.578e+11Hz -0.018201 -0.0156784
+ 1.579e+11Hz -0.0182068 -0.0156722
+ 1.58e+11Hz -0.0182125 -0.0156662
+ 1.581e+11Hz -0.0182183 -0.0156602
+ 1.582e+11Hz -0.018224 -0.0156543
+ 1.583e+11Hz -0.0182298 -0.0156484
+ 1.584e+11Hz -0.0182355 -0.0156427
+ 1.585e+11Hz -0.0182412 -0.0156369
+ 1.586e+11Hz -0.0182469 -0.0156313
+ 1.587e+11Hz -0.0182526 -0.0156257
+ 1.588e+11Hz -0.0182583 -0.0156202
+ 1.589e+11Hz -0.018264 -0.0156148
+ 1.59e+11Hz -0.0182697 -0.0156094
+ 1.591e+11Hz -0.0182754 -0.0156041
+ 1.592e+11Hz -0.0182811 -0.0155988
+ 1.593e+11Hz -0.0182868 -0.0155937
+ 1.594e+11Hz -0.0182925 -0.0155886
+ 1.595e+11Hz -0.0182982 -0.0155835
+ 1.596e+11Hz -0.0183039 -0.0155786
+ 1.597e+11Hz -0.0183096 -0.0155737
+ 1.598e+11Hz -0.0183153 -0.0155689
+ 1.599e+11Hz -0.018321 -0.0155641
+ 1.6e+11Hz -0.0183267 -0.0155595
+ 1.601e+11Hz -0.0183325 -0.0155549
+ 1.602e+11Hz -0.0183382 -0.0155503
+ 1.603e+11Hz -0.0183439 -0.0155459
+ 1.604e+11Hz -0.0183497 -0.0155415
+ 1.605e+11Hz -0.0183555 -0.0155371
+ 1.606e+11Hz -0.0183612 -0.0155329
+ 1.607e+11Hz -0.018367 -0.0155287
+ 1.608e+11Hz -0.0183728 -0.0155246
+ 1.609e+11Hz -0.0183786 -0.0155206
+ 1.61e+11Hz -0.0183845 -0.0155166
+ 1.611e+11Hz -0.0183903 -0.0155127
+ 1.612e+11Hz -0.0183962 -0.0155089
+ 1.613e+11Hz -0.0184021 -0.0155051
+ 1.614e+11Hz -0.018408 -0.0155014
+ 1.615e+11Hz -0.0184139 -0.0154978
+ 1.616e+11Hz -0.0184199 -0.0154943
+ 1.617e+11Hz -0.0184258 -0.0154908
+ 1.618e+11Hz -0.0184318 -0.0154874
+ 1.619e+11Hz -0.0184378 -0.0154841
+ 1.62e+11Hz -0.0184439 -0.0154808
+ 1.621e+11Hz -0.0184499 -0.0154776
+ 1.622e+11Hz -0.018456 -0.0154745
+ 1.623e+11Hz -0.0184622 -0.0154714
+ 1.624e+11Hz -0.0184683 -0.0154684
+ 1.625e+11Hz -0.0184745 -0.0154655
+ 1.626e+11Hz -0.0184807 -0.0154627
+ 1.627e+11Hz -0.018487 -0.0154599
+ 1.628e+11Hz -0.0184933 -0.0154572
+ 1.629e+11Hz -0.0184996 -0.0154546
+ 1.63e+11Hz -0.0185059 -0.015452
+ 1.631e+11Hz -0.0185123 -0.0154495
+ 1.632e+11Hz -0.0185187 -0.0154471
+ 1.633e+11Hz -0.0185252 -0.0154447
+ 1.634e+11Hz -0.0185317 -0.0154424
+ 1.635e+11Hz -0.0185383 -0.0154402
+ 1.636e+11Hz -0.0185448 -0.015438
+ 1.637e+11Hz -0.0185515 -0.0154359
+ 1.638e+11Hz -0.0185582 -0.0154339
+ 1.639e+11Hz -0.0185649 -0.0154319
+ 1.64e+11Hz -0.0185716 -0.01543
+ 1.641e+11Hz -0.0185785 -0.0154281
+ 1.642e+11Hz -0.0185853 -0.0154264
+ 1.643e+11Hz -0.0185922 -0.0154247
+ 1.644e+11Hz -0.0185992 -0.015423
+ 1.645e+11Hz -0.0186062 -0.0154214
+ 1.646e+11Hz -0.0186132 -0.0154199
+ 1.647e+11Hz -0.0186204 -0.0154184
+ 1.648e+11Hz -0.0186275 -0.015417
+ 1.649e+11Hz -0.0186347 -0.0154157
+ 1.65e+11Hz -0.018642 -0.0154144
+ 1.651e+11Hz -0.0186494 -0.0154132
+ 1.652e+11Hz -0.0186567 -0.015412
+ 1.653e+11Hz -0.0186642 -0.0154109
+ 1.654e+11Hz -0.0186717 -0.0154098
+ 1.655e+11Hz -0.0186793 -0.0154088
+ 1.656e+11Hz -0.0186869 -0.0154079
+ 1.657e+11Hz -0.0186946 -0.015407
+ 1.658e+11Hz -0.0187023 -0.0154062
+ 1.659e+11Hz -0.0187102 -0.0154054
+ 1.66e+11Hz -0.0187181 -0.0154047
+ 1.661e+11Hz -0.018726 -0.015404
+ 1.662e+11Hz -0.018734 -0.0154034
+ 1.663e+11Hz -0.0187421 -0.0154028
+ 1.664e+11Hz -0.0187503 -0.0154023
+ 1.665e+11Hz -0.0187585 -0.0154018
+ 1.666e+11Hz -0.0187668 -0.0154014
+ 1.667e+11Hz -0.0187751 -0.0154011
+ 1.668e+11Hz -0.0187836 -0.0154007
+ 1.669e+11Hz -0.0187921 -0.0154005
+ 1.67e+11Hz -0.0188007 -0.0154002
+ 1.671e+11Hz -0.0188093 -0.0154
+ 1.672e+11Hz -0.0188181 -0.0153999
+ 1.673e+11Hz -0.0188269 -0.0153998
+ 1.674e+11Hz -0.0188358 -0.0153997
+ 1.675e+11Hz -0.0188447 -0.0153997
+ 1.676e+11Hz -0.0188538 -0.0153997
+ 1.677e+11Hz -0.0188629 -0.0153998
+ 1.678e+11Hz -0.0188721 -0.0153999
+ 1.679e+11Hz -0.0188814 -0.0154
+ 1.68e+11Hz -0.0188908 -0.0154002
+ 1.681e+11Hz -0.0189002 -0.0154004
+ 1.682e+11Hz -0.0189097 -0.0154007
+ 1.683e+11Hz -0.0189194 -0.015401
+ 1.684e+11Hz -0.0189291 -0.0154013
+ 1.685e+11Hz -0.0189388 -0.0154016
+ 1.686e+11Hz -0.0189487 -0.015402
+ 1.687e+11Hz -0.0189587 -0.0154024
+ 1.688e+11Hz -0.0189687 -0.0154028
+ 1.689e+11Hz -0.0189789 -0.0154033
+ 1.69e+11Hz -0.0189891 -0.0154037
+ 1.691e+11Hz -0.0189994 -0.0154043
+ 1.692e+11Hz -0.0190098 -0.0154048
+ 1.693e+11Hz -0.0190203 -0.0154053
+ 1.694e+11Hz -0.0190309 -0.0154059
+ 1.695e+11Hz -0.0190415 -0.0154065
+ 1.696e+11Hz -0.0190523 -0.0154071
+ 1.697e+11Hz -0.0190632 -0.0154078
+ 1.698e+11Hz -0.0190741 -0.0154084
+ 1.699e+11Hz -0.0190852 -0.0154091
+ 1.7e+11Hz -0.0190963 -0.0154098
+ 1.701e+11Hz -0.0191075 -0.0154105
+ 1.702e+11Hz -0.0191189 -0.0154112
+ 1.703e+11Hz -0.0191303 -0.0154119
+ 1.704e+11Hz -0.0191418 -0.0154126
+ 1.705e+11Hz -0.0191534 -0.0154133
+ 1.706e+11Hz -0.0191651 -0.0154141
+ 1.707e+11Hz -0.0191769 -0.0154148
+ 1.708e+11Hz -0.0191889 -0.0154156
+ 1.709e+11Hz -0.0192009 -0.0154163
+ 1.71e+11Hz -0.019213 -0.0154171
+ 1.711e+11Hz -0.0192252 -0.0154179
+ 1.712e+11Hz -0.0192375 -0.0154186
+ 1.713e+11Hz -0.0192499 -0.0154194
+ 1.714e+11Hz -0.0192623 -0.0154201
+ 1.715e+11Hz -0.0192749 -0.0154209
+ 1.716e+11Hz -0.0192876 -0.0154216
+ 1.717e+11Hz -0.0193004 -0.0154224
+ 1.718e+11Hz -0.0193133 -0.0154231
+ 1.719e+11Hz -0.0193263 -0.0154238
+ 1.72e+11Hz -0.0193394 -0.0154246
+ 1.721e+11Hz -0.0193526 -0.0154253
+ 1.722e+11Hz -0.0193659 -0.015426
+ 1.723e+11Hz -0.0193793 -0.0154266
+ 1.724e+11Hz -0.0193928 -0.0154273
+ 1.725e+11Hz -0.0194064 -0.0154279
+ 1.726e+11Hz -0.0194201 -0.0154285
+ 1.727e+11Hz -0.0194339 -0.0154292
+ 1.728e+11Hz -0.0194478 -0.0154297
+ 1.729e+11Hz -0.0194618 -0.0154303
+ 1.73e+11Hz -0.0194759 -0.0154308
+ 1.731e+11Hz -0.0194901 -0.0154313
+ 1.732e+11Hz -0.0195044 -0.0154318
+ 1.733e+11Hz -0.0195188 -0.0154323
+ 1.734e+11Hz -0.0195334 -0.0154327
+ 1.735e+11Hz -0.019548 -0.0154331
+ 1.736e+11Hz -0.0195627 -0.0154335
+ 1.737e+11Hz -0.0195775 -0.0154338
+ 1.738e+11Hz -0.0195924 -0.0154341
+ 1.739e+11Hz -0.0196074 -0.0154343
+ 1.74e+11Hz -0.0196225 -0.0154346
+ 1.741e+11Hz -0.0196377 -0.0154348
+ 1.742e+11Hz -0.019653 -0.0154349
+ 1.743e+11Hz -0.0196684 -0.015435
+ 1.744e+11Hz -0.0196839 -0.0154351
+ 1.745e+11Hz -0.0196995 -0.0154351
+ 1.746e+11Hz -0.0197153 -0.015435
+ 1.747e+11Hz -0.0197311 -0.015435
+ 1.748e+11Hz -0.019747 -0.0154348
+ 1.749e+11Hz -0.019763 -0.0154347
+ 1.75e+11Hz -0.019779 -0.0154344
+ 1.751e+11Hz -0.0197952 -0.0154342
+ 1.752e+11Hz -0.0198115 -0.0154338
+ 1.753e+11Hz -0.0198279 -0.0154335
+ 1.754e+11Hz -0.0198444 -0.015433
+ 1.755e+11Hz -0.019861 -0.0154325
+ 1.756e+11Hz -0.0198776 -0.015432
+ 1.757e+11Hz -0.0198944 -0.0154313
+ 1.758e+11Hz -0.0199112 -0.0154307
+ 1.759e+11Hz -0.0199282 -0.0154299
+ 1.76e+11Hz -0.0199452 -0.0154291
+ 1.761e+11Hz -0.0199624 -0.0154283
+ 1.762e+11Hz -0.0199796 -0.0154273
+ 1.763e+11Hz -0.0199969 -0.0154263
+ 1.764e+11Hz -0.0200143 -0.0154252
+ 1.765e+11Hz -0.0200318 -0.0154241
+ 1.766e+11Hz -0.0200494 -0.0154229
+ 1.767e+11Hz -0.020067 -0.0154216
+ 1.768e+11Hz -0.0200848 -0.0154202
+ 1.769e+11Hz -0.0201026 -0.0154188
+ 1.77e+11Hz -0.0201206 -0.0154173
+ 1.771e+11Hz -0.0201386 -0.0154157
+ 1.772e+11Hz -0.0201567 -0.015414
+ 1.773e+11Hz -0.0201749 -0.0154123
+ 1.774e+11Hz -0.0201931 -0.0154105
+ 1.775e+11Hz -0.0202115 -0.0154086
+ 1.776e+11Hz -0.0202299 -0.0154066
+ 1.777e+11Hz -0.0202484 -0.0154045
+ 1.778e+11Hz -0.020267 -0.0154023
+ 1.779e+11Hz -0.0202857 -0.0154001
+ 1.78e+11Hz -0.0203044 -0.0153977
+ 1.781e+11Hz -0.0203232 -0.0153953
+ 1.782e+11Hz -0.0203421 -0.0153928
+ 1.783e+11Hz -0.0203611 -0.0153902
+ 1.784e+11Hz -0.0203801 -0.0153875
+ 1.785e+11Hz -0.0203993 -0.0153847
+ 1.786e+11Hz -0.0204184 -0.0153818
+ 1.787e+11Hz -0.0204377 -0.0153788
+ 1.788e+11Hz -0.020457 -0.0153757
+ 1.789e+11Hz -0.0204764 -0.0153726
+ 1.79e+11Hz -0.0204959 -0.0153693
+ 1.791e+11Hz -0.0205154 -0.0153659
+ 1.792e+11Hz -0.020535 -0.0153624
+ 1.793e+11Hz -0.0205547 -0.0153589
+ 1.794e+11Hz -0.0205744 -0.0153552
+ 1.795e+11Hz -0.0205942 -0.0153514
+ 1.796e+11Hz -0.0206141 -0.0153475
+ 1.797e+11Hz -0.020634 -0.0153435
+ 1.798e+11Hz -0.020654 -0.0153394
+ 1.799e+11Hz -0.020674 -0.0153352
+ 1.8e+11Hz -0.0206941 -0.0153309
+ 1.801e+11Hz -0.0207143 -0.0153265
+ 1.802e+11Hz -0.0207345 -0.015322
+ 1.803e+11Hz -0.0207547 -0.0153174
+ 1.804e+11Hz -0.020775 -0.0153126
+ 1.805e+11Hz -0.0207954 -0.0153078
+ 1.806e+11Hz -0.0208158 -0.0153028
+ 1.807e+11Hz -0.0208363 -0.0152977
+ 1.808e+11Hz -0.0208568 -0.0152925
+ 1.809e+11Hz -0.0208773 -0.0152872
+ 1.81e+11Hz -0.0208979 -0.0152818
+ 1.811e+11Hz -0.0209186 -0.0152762
+ 1.812e+11Hz -0.0209392 -0.0152706
+ 1.813e+11Hz -0.02096 -0.0152648
+ 1.814e+11Hz -0.0209807 -0.0152589
+ 1.815e+11Hz -0.0210015 -0.0152529
+ 1.816e+11Hz -0.0210224 -0.0152467
+ 1.817e+11Hz -0.0210433 -0.0152405
+ 1.818e+11Hz -0.0210642 -0.0152341
+ 1.819e+11Hz -0.0210851 -0.0152276
+ 1.82e+11Hz -0.0211061 -0.015221
+ 1.821e+11Hz -0.0211271 -0.0152143
+ 1.822e+11Hz -0.0211481 -0.0152074
+ 1.823e+11Hz -0.0211692 -0.0152004
+ 1.824e+11Hz -0.0211903 -0.0151933
+ 1.825e+11Hz -0.0212114 -0.0151861
+ 1.826e+11Hz -0.0212325 -0.0151787
+ 1.827e+11Hz -0.0212537 -0.0151712
+ 1.828e+11Hz -0.0212749 -0.0151636
+ 1.829e+11Hz -0.0212961 -0.0151559
+ 1.83e+11Hz -0.0213173 -0.015148
+ 1.831e+11Hz -0.0213385 -0.0151401
+ 1.832e+11Hz -0.0213598 -0.015132
+ 1.833e+11Hz -0.021381 -0.0151237
+ 1.834e+11Hz -0.0214023 -0.0151154
+ 1.835e+11Hz -0.0214236 -0.0151069
+ 1.836e+11Hz -0.0214449 -0.0150982
+ 1.837e+11Hz -0.0214662 -0.0150895
+ 1.838e+11Hz -0.0214875 -0.0150806
+ 1.839e+11Hz -0.0215088 -0.0150716
+ 1.84e+11Hz -0.0215301 -0.0150625
+ 1.841e+11Hz -0.0215515 -0.0150532
+ 1.842e+11Hz -0.0215728 -0.0150438
+ 1.843e+11Hz -0.0215941 -0.0150343
+ 1.844e+11Hz -0.0216154 -0.0150247
+ 1.845e+11Hz -0.0216367 -0.0150149
+ 1.846e+11Hz -0.021658 -0.015005
+ 1.847e+11Hz -0.0216793 -0.014995
+ 1.848e+11Hz -0.0217006 -0.0149848
+ 1.849e+11Hz -0.0217219 -0.0149745
+ 1.85e+11Hz -0.0217432 -0.0149641
+ 1.851e+11Hz -0.0217644 -0.0149536
+ 1.852e+11Hz -0.0217857 -0.0149429
+ 1.853e+11Hz -0.0218069 -0.0149321
+ 1.854e+11Hz -0.0218281 -0.0149212
+ 1.855e+11Hz -0.0218493 -0.0149101
+ 1.856e+11Hz -0.0218705 -0.0148989
+ 1.857e+11Hz -0.0218916 -0.0148876
+ 1.858e+11Hz -0.0219128 -0.0148761
+ 1.859e+11Hz -0.0219339 -0.0148646
+ 1.86e+11Hz -0.0219549 -0.0148529
+ 1.861e+11Hz -0.021976 -0.014841
+ 1.862e+11Hz -0.021997 -0.0148291
+ 1.863e+11Hz -0.022018 -0.014817
+ 1.864e+11Hz -0.022039 -0.0148048
+ 1.865e+11Hz -0.0220599 -0.0147925
+ 1.866e+11Hz -0.0220808 -0.01478
+ 1.867e+11Hz -0.0221016 -0.0147674
+ 1.868e+11Hz -0.0221224 -0.0147547
+ 1.869e+11Hz -0.0221432 -0.0147419
+ 1.87e+11Hz -0.0221639 -0.0147289
+ 1.871e+11Hz -0.0221846 -0.0147158
+ 1.872e+11Hz -0.0222053 -0.0147026
+ 1.873e+11Hz -0.0222259 -0.0146893
+ 1.874e+11Hz -0.0222464 -0.0146758
+ 1.875e+11Hz -0.0222669 -0.0146623
+ 1.876e+11Hz -0.0222874 -0.0146486
+ 1.877e+11Hz -0.0223078 -0.0146348
+ 1.878e+11Hz -0.0223282 -0.0146208
+ 1.879e+11Hz -0.0223485 -0.0146068
+ 1.88e+11Hz -0.0223687 -0.0145926
+ 1.881e+11Hz -0.0223889 -0.0145783
+ 1.882e+11Hz -0.022409 -0.0145639
+ 1.883e+11Hz -0.0224291 -0.0145494
+ 1.884e+11Hz -0.0224491 -0.0145347
+ 1.885e+11Hz -0.0224691 -0.01452
+ 1.886e+11Hz -0.022489 -0.0145051
+ 1.887e+11Hz -0.0225088 -0.0144901
+ 1.888e+11Hz -0.0225286 -0.014475
+ 1.889e+11Hz -0.0225482 -0.0144598
+ 1.89e+11Hz -0.0225679 -0.0144445
+ 1.891e+11Hz -0.0225874 -0.0144291
+ 1.892e+11Hz -0.0226069 -0.0144135
+ 1.893e+11Hz -0.0226263 -0.0143979
+ 1.894e+11Hz -0.0226457 -0.0143821
+ 1.895e+11Hz -0.0226649 -0.0143663
+ 1.896e+11Hz -0.0226841 -0.0143503
+ 1.897e+11Hz -0.0227032 -0.0143342
+ 1.898e+11Hz -0.0227223 -0.014318
+ 1.899e+11Hz -0.0227412 -0.0143017
+ 1.9e+11Hz -0.0227601 -0.0142854
+ 1.901e+11Hz -0.0227789 -0.0142689
+ 1.902e+11Hz -0.0227976 -0.0142523
+ 1.903e+11Hz -0.0228162 -0.0142356
+ 1.904e+11Hz -0.0228348 -0.0142188
+ 1.905e+11Hz -0.0228532 -0.0142019
+ 1.906e+11Hz -0.0228716 -0.014185
+ 1.907e+11Hz -0.0228899 -0.0141679
+ 1.908e+11Hz -0.0229081 -0.0141507
+ 1.909e+11Hz -0.0229262 -0.0141335
+ 1.91e+11Hz -0.0229442 -0.0141161
+ 1.911e+11Hz -0.0229621 -0.0140987
+ 1.912e+11Hz -0.0229799 -0.0140812
+ 1.913e+11Hz -0.0229976 -0.0140635
+ 1.914e+11Hz -0.0230153 -0.0140458
+ 1.915e+11Hz -0.0230328 -0.014028
+ 1.916e+11Hz -0.0230503 -0.0140102
+ 1.917e+11Hz -0.0230676 -0.0139922
+ 1.918e+11Hz -0.0230848 -0.0139742
+ 1.919e+11Hz -0.023102 -0.0139561
+ 1.92e+11Hz -0.023119 -0.0139379
+ 1.921e+11Hz -0.023136 -0.0139196
+ 1.922e+11Hz -0.0231528 -0.0139013
+ 1.923e+11Hz -0.0231695 -0.0138828
+ 1.924e+11Hz -0.0231862 -0.0138644
+ 1.925e+11Hz -0.0232027 -0.0138458
+ 1.926e+11Hz -0.0232191 -0.0138271
+ 1.927e+11Hz -0.0232354 -0.0138084
+ 1.928e+11Hz -0.0232516 -0.0137897
+ 1.929e+11Hz -0.0232677 -0.0137708
+ 1.93e+11Hz -0.0232837 -0.0137519
+ 1.931e+11Hz -0.0232996 -0.013733
+ 1.932e+11Hz -0.0233154 -0.0137139
+ 1.933e+11Hz -0.0233311 -0.0136948
+ 1.934e+11Hz -0.0233466 -0.0136757
+ 1.935e+11Hz -0.0233621 -0.0136565
+ 1.936e+11Hz -0.0233774 -0.0136372
+ 1.937e+11Hz -0.0233926 -0.0136179
+ 1.938e+11Hz -0.0234077 -0.0135985
+ 1.939e+11Hz -0.0234227 -0.0135791
+ 1.94e+11Hz -0.0234376 -0.0135596
+ 1.941e+11Hz -0.0234523 -0.0135401
+ 1.942e+11Hz -0.023467 -0.0135206
+ 1.943e+11Hz -0.0234815 -0.0135009
+ 1.944e+11Hz -0.0234959 -0.0134813
+ 1.945e+11Hz -0.0235102 -0.0134616
+ 1.946e+11Hz -0.0235244 -0.0134419
+ 1.947e+11Hz -0.0235385 -0.0134221
+ 1.948e+11Hz -0.0235525 -0.0134023
+ 1.949e+11Hz -0.0235663 -0.0133824
+ 1.95e+11Hz -0.02358 -0.0133625
+ 1.951e+11Hz -0.0235936 -0.0133426
+ 1.952e+11Hz -0.0236071 -0.0133227
+ 1.953e+11Hz -0.0236205 -0.0133027
+ 1.954e+11Hz -0.0236337 -0.0132827
+ 1.955e+11Hz -0.0236469 -0.0132627
+ 1.956e+11Hz -0.0236599 -0.0132426
+ 1.957e+11Hz -0.0236728 -0.0132226
+ 1.958e+11Hz -0.0236856 -0.0132025
+ 1.959e+11Hz -0.0236982 -0.0131824
+ 1.96e+11Hz -0.0237108 -0.0131622
+ 1.961e+11Hz -0.0237232 -0.0131421
+ 1.962e+11Hz -0.0237355 -0.0131219
+ 1.963e+11Hz -0.0237477 -0.0131018
+ 1.964e+11Hz -0.0237598 -0.0130816
+ 1.965e+11Hz -0.0237718 -0.0130614
+ 1.966e+11Hz -0.0237836 -0.0130412
+ 1.967e+11Hz -0.0237953 -0.013021
+ 1.968e+11Hz -0.0238069 -0.0130008
+ 1.969e+11Hz -0.0238184 -0.0129806
+ 1.97e+11Hz -0.0238298 -0.0129604
+ 1.971e+11Hz -0.0238411 -0.0129402
+ 1.972e+11Hz -0.0238522 -0.01292
+ 1.973e+11Hz -0.0238633 -0.0128998
+ 1.974e+11Hz -0.0238742 -0.0128796
+ 1.975e+11Hz -0.023885 -0.0128594
+ 1.976e+11Hz -0.0238957 -0.0128392
+ 1.977e+11Hz -0.0239063 -0.012819
+ 1.978e+11Hz -0.0239168 -0.0127989
+ 1.979e+11Hz -0.0239271 -0.0127787
+ 1.98e+11Hz -0.0239374 -0.0127586
+ 1.981e+11Hz -0.0239475 -0.0127385
+ 1.982e+11Hz -0.0239575 -0.0127184
+ 1.983e+11Hz -0.0239675 -0.0126984
+ 1.984e+11Hz -0.0239773 -0.0126783
+ 1.985e+11Hz -0.023987 -0.0126583
+ 1.986e+11Hz -0.0239966 -0.0126383
+ 1.987e+11Hz -0.0240061 -0.0126183
+ 1.988e+11Hz -0.0240155 -0.0125984
+ 1.989e+11Hz -0.0240247 -0.0125785
+ 1.99e+11Hz -0.0240339 -0.0125586
+ 1.991e+11Hz -0.024043 -0.0125388
+ 1.992e+11Hz -0.024052 -0.012519
+ 1.993e+11Hz -0.0240608 -0.0124992
+ 1.994e+11Hz -0.0240696 -0.0124795
+ 1.995e+11Hz -0.0240783 -0.0124598
+ 1.996e+11Hz -0.0240869 -0.0124401
+ 1.997e+11Hz -0.0240954 -0.0124205
+ 1.998e+11Hz -0.0241037 -0.0124009
+ 1.999e+11Hz -0.024112 -0.0123814
+ 2e+11Hz -0.0241202 -0.0123619
+ 2.001e+11Hz -0.0241283 -0.0123425
+ 2.002e+11Hz -0.0241364 -0.0123231
+ 2.003e+11Hz -0.0241443 -0.0123038
+ 2.004e+11Hz -0.0241521 -0.0122845
+ 2.005e+11Hz -0.0241599 -0.0122653
+ 2.006e+11Hz -0.0241675 -0.0122461
+ 2.007e+11Hz -0.0241751 -0.012227
+ 2.008e+11Hz -0.0241826 -0.0122079
+ 2.009e+11Hz -0.02419 -0.0121889
+ 2.01e+11Hz -0.0241974 -0.01217
+ 2.011e+11Hz -0.0242046 -0.0121511
+ 2.012e+11Hz -0.0242118 -0.0121323
+ 2.013e+11Hz -0.0242189 -0.0121136
+ 2.014e+11Hz -0.024226 -0.0120949
+ 2.015e+11Hz -0.0242329 -0.0120762
+ 2.016e+11Hz -0.0242398 -0.0120577
+ 2.017e+11Hz -0.0242466 -0.0120392
+ 2.018e+11Hz -0.0242534 -0.0120208
+ 2.019e+11Hz -0.0242601 -0.0120024
+ 2.02e+11Hz -0.0242667 -0.0119841
+ 2.021e+11Hz -0.0242732 -0.0119659
+ 2.022e+11Hz -0.0242797 -0.0119478
+ 2.023e+11Hz -0.0242861 -0.0119297
+ 2.024e+11Hz -0.0242925 -0.0119118
+ 2.025e+11Hz -0.0242988 -0.0118938
+ 2.026e+11Hz -0.0243051 -0.011876
+ 2.027e+11Hz -0.0243113 -0.0118582
+ 2.028e+11Hz -0.0243175 -0.0118406
+ 2.029e+11Hz -0.0243236 -0.011823
+ 2.03e+11Hz -0.0243296 -0.0118054
+ 2.031e+11Hz -0.0243357 -0.011788
+ 2.032e+11Hz -0.0243416 -0.0117706
+ 2.033e+11Hz -0.0243476 -0.0117533
+ 2.034e+11Hz -0.0243535 -0.0117361
+ 2.035e+11Hz -0.0243593 -0.011719
+ 2.036e+11Hz -0.0243651 -0.011702
+ 2.037e+11Hz -0.0243709 -0.011685
+ 2.038e+11Hz -0.0243767 -0.0116682
+ 2.039e+11Hz -0.0243824 -0.0116514
+ 2.04e+11Hz -0.0243881 -0.0116347
+ 2.041e+11Hz -0.0243938 -0.0116181
+ 2.042e+11Hz -0.0243994 -0.0116016
+ 2.043e+11Hz -0.024405 -0.0115851
+ 2.044e+11Hz -0.0244106 -0.0115688
+ 2.045e+11Hz -0.0244162 -0.0115525
+ 2.046e+11Hz -0.0244218 -0.0115363
+ 2.047e+11Hz -0.0244273 -0.0115202
+ 2.048e+11Hz -0.0244329 -0.0115042
+ 2.049e+11Hz -0.0244384 -0.0114883
+ 2.05e+11Hz -0.0244439 -0.0114724
+ 2.051e+11Hz -0.0244495 -0.0114567
+ 2.052e+11Hz -0.024455 -0.011441
+ 2.053e+11Hz -0.0244605 -0.0114254
+ 2.054e+11Hz -0.024466 -0.0114099
+ 2.055e+11Hz -0.0244715 -0.0113945
+ 2.056e+11Hz -0.0244771 -0.0113792
+ 2.057e+11Hz -0.0244826 -0.011364
+ 2.058e+11Hz -0.0244881 -0.0113489
+ 2.059e+11Hz -0.0244937 -0.0113338
+ 2.06e+11Hz -0.0244993 -0.0113188
+ 2.061e+11Hz -0.0245049 -0.0113039
+ 2.062e+11Hz -0.0245105 -0.0112891
+ 2.063e+11Hz -0.0245161 -0.0112744
+ 2.064e+11Hz -0.0245217 -0.0112598
+ 2.065e+11Hz -0.0245274 -0.0112452
+ 2.066e+11Hz -0.0245331 -0.0112307
+ 2.067e+11Hz -0.0245389 -0.0112163
+ 2.068e+11Hz -0.0245446 -0.011202
+ 2.069e+11Hz -0.0245504 -0.0111878
+ 2.07e+11Hz -0.0245563 -0.0111737
+ 2.071e+11Hz -0.0245621 -0.0111596
+ 2.072e+11Hz -0.024568 -0.0111456
+ 2.073e+11Hz -0.024574 -0.0111317
+ 2.074e+11Hz -0.02458 -0.0111178
+ 2.075e+11Hz -0.0245861 -0.0111041
+ 2.076e+11Hz -0.0245921 -0.0110904
+ 2.077e+11Hz -0.0245983 -0.0110768
+ 2.078e+11Hz -0.0246045 -0.0110632
+ 2.079e+11Hz -0.0246107 -0.0110497
+ 2.08e+11Hz -0.0246171 -0.0110363
+ 2.081e+11Hz -0.0246234 -0.011023
+ 2.082e+11Hz -0.0246299 -0.0110097
+ 2.083e+11Hz -0.0246364 -0.0109965
+ 2.084e+11Hz -0.0246429 -0.0109834
+ 2.085e+11Hz -0.0246496 -0.0109703
+ 2.086e+11Hz -0.0246563 -0.0109573
+ 2.087e+11Hz -0.024663 -0.0109444
+ 2.088e+11Hz -0.0246699 -0.0109315
+ 2.089e+11Hz -0.0246768 -0.0109186
+ 2.09e+11Hz -0.0246838 -0.0109058
+ 2.091e+11Hz -0.0246909 -0.0108931
+ 2.092e+11Hz -0.024698 -0.0108804
+ 2.093e+11Hz -0.0247053 -0.0108678
+ 2.094e+11Hz -0.0247126 -0.0108553
+ 2.095e+11Hz -0.02472 -0.0108427
+ 2.096e+11Hz -0.0247275 -0.0108302
+ 2.097e+11Hz -0.0247351 -0.0108178
+ 2.098e+11Hz -0.0247428 -0.0108054
+ 2.099e+11Hz -0.0247505 -0.0107931
+ 2.1e+11Hz -0.0247584 -0.0107807
+ 2.101e+11Hz -0.0247664 -0.0107685
+ 2.102e+11Hz -0.0247744 -0.0107562
+ 2.103e+11Hz -0.0247826 -0.010744
+ 2.104e+11Hz -0.0247909 -0.0107318
+ 2.105e+11Hz -0.0247992 -0.0107197
+ 2.106e+11Hz -0.0248077 -0.0107075
+ 2.107e+11Hz -0.0248163 -0.0106954
+ 2.108e+11Hz -0.024825 -0.0106833
+ 2.109e+11Hz -0.0248338 -0.0106712
+ 2.11e+11Hz -0.0248427 -0.0106592
+ 2.111e+11Hz -0.0248517 -0.0106472
+ 2.112e+11Hz -0.0248608 -0.0106351
+ 2.113e+11Hz -0.02487 -0.0106231
+ 2.114e+11Hz -0.0248794 -0.0106111
+ 2.115e+11Hz -0.0248889 -0.0105991
+ 2.116e+11Hz -0.0248985 -0.0105871
+ 2.117e+11Hz -0.0249082 -0.0105751
+ 2.118e+11Hz -0.024918 -0.010563
+ 2.119e+11Hz -0.024928 -0.010551
+ 2.12e+11Hz -0.024938 -0.010539
+ 2.121e+11Hz -0.0249482 -0.0105269
+ 2.122e+11Hz -0.0249586 -0.0105149
+ 2.123e+11Hz -0.024969 -0.0105028
+ 2.124e+11Hz -0.0249796 -0.0104907
+ 2.125e+11Hz -0.0249903 -0.0104786
+ 2.126e+11Hz -0.0250011 -0.0104665
+ 2.127e+11Hz -0.025012 -0.0104543
+ 2.128e+11Hz -0.0250231 -0.0104421
+ 2.129e+11Hz -0.0250343 -0.0104299
+ 2.13e+11Hz -0.0250456 -0.0104176
+ 2.131e+11Hz -0.0250571 -0.0104053
+ 2.132e+11Hz -0.0250687 -0.0103929
+ 2.133e+11Hz -0.0250804 -0.0103805
+ 2.134e+11Hz -0.0250923 -0.0103681
+ 2.135e+11Hz -0.0251043 -0.0103556
+ 2.136e+11Hz -0.0251164 -0.010343
+ 2.137e+11Hz -0.0251286 -0.0103304
+ 2.138e+11Hz -0.025141 -0.0103177
+ 2.139e+11Hz -0.0251535 -0.010305
+ 2.14e+11Hz -0.0251661 -0.0102922
+ 2.141e+11Hz -0.0251789 -0.0102793
+ 2.142e+11Hz -0.0251918 -0.0102663
+ 2.143e+11Hz -0.0252048 -0.0102533
+ 2.144e+11Hz -0.025218 -0.0102402
+ 2.145e+11Hz -0.0252313 -0.010227
+ 2.146e+11Hz -0.0252447 -0.0102137
+ 2.147e+11Hz -0.0252583 -0.0102004
+ 2.148e+11Hz -0.0252719 -0.0101869
+ 2.149e+11Hz -0.0252857 -0.0101733
+ 2.15e+11Hz -0.0252997 -0.0101597
+ 2.151e+11Hz -0.0253137 -0.0101459
+ 2.152e+11Hz -0.0253279 -0.0101321
+ 2.153e+11Hz -0.0253422 -0.0101181
+ 2.154e+11Hz -0.0253567 -0.010104
+ 2.155e+11Hz -0.0253713 -0.0100898
+ 2.156e+11Hz -0.0253859 -0.0100755
+ 2.157e+11Hz -0.0254008 -0.0100611
+ 2.158e+11Hz -0.0254157 -0.0100466
+ 2.159e+11Hz -0.0254307 -0.0100319
+ 2.16e+11Hz -0.0254459 -0.0100171
+ 2.161e+11Hz -0.0254612 -0.0100021
+ 2.162e+11Hz -0.0254766 -0.00998704
+ 2.163e+11Hz -0.0254921 -0.00997182
+ 2.164e+11Hz -0.0255078 -0.00995646
+ 2.165e+11Hz -0.0255235 -0.00994096
+ 2.166e+11Hz -0.0255394 -0.0099253
+ 2.167e+11Hz -0.0255553 -0.00990949
+ 2.168e+11Hz -0.0255714 -0.00989353
+ 2.169e+11Hz -0.0255876 -0.00987741
+ 2.17e+11Hz -0.0256039 -0.00986113
+ 2.171e+11Hz -0.0256203 -0.00984469
+ 2.172e+11Hz -0.0256368 -0.00982807
+ 2.173e+11Hz -0.0256533 -0.00981129
+ 2.174e+11Hz -0.02567 -0.00979434
+ 2.175e+11Hz -0.0256868 -0.00977721
+ 2.176e+11Hz -0.0257037 -0.0097599
+ 2.177e+11Hz -0.0257206 -0.00974241
+ 2.178e+11Hz -0.0257377 -0.00972474
+ 2.179e+11Hz -0.0257548 -0.00970688
+ 2.18e+11Hz -0.025772 -0.00968883
+ 2.181e+11Hz -0.0257893 -0.00967059
+ 2.182e+11Hz -0.0258067 -0.00965215
+ 2.183e+11Hz -0.0258242 -0.00963351
+ 2.184e+11Hz -0.0258417 -0.00961468
+ 2.185e+11Hz -0.0258593 -0.00959564
+ 2.186e+11Hz -0.025877 -0.00957639
+ 2.187e+11Hz -0.0258947 -0.00955694
+ 2.188e+11Hz -0.0259125 -0.00953728
+ 2.189e+11Hz -0.0259304 -0.0095174
+ 2.19e+11Hz -0.0259483 -0.00949731
+ 2.191e+11Hz -0.0259663 -0.00947699
+ 2.192e+11Hz -0.0259843 -0.00945646
+ 2.193e+11Hz -0.0260024 -0.00943571
+ 2.194e+11Hz -0.0260205 -0.00941473
+ 2.195e+11Hz -0.0260386 -0.00939352
+ 2.196e+11Hz -0.0260568 -0.00937209
+ 2.197e+11Hz -0.0260751 -0.00935042
+ 2.198e+11Hz -0.0260933 -0.00932852
+ 2.199e+11Hz -0.0261116 -0.00930638
+ 2.2e+11Hz -0.02613 -0.00928401
+ 2.201e+11Hz -0.0261483 -0.00926139
+ 2.202e+11Hz -0.0261667 -0.00923854
+ 2.203e+11Hz -0.0261851 -0.00921544
+ 2.204e+11Hz -0.0262035 -0.00919209
+ 2.205e+11Hz -0.0262219 -0.0091685
+ 2.206e+11Hz -0.0262403 -0.00914466
+ 2.207e+11Hz -0.0262587 -0.00912057
+ 2.208e+11Hz -0.0262771 -0.00909623
+ 2.209e+11Hz -0.0262955 -0.00907164
+ 2.21e+11Hz -0.0263139 -0.00904679
+ 2.211e+11Hz -0.0263323 -0.00902169
+ 2.212e+11Hz -0.0263506 -0.00899633
+ 2.213e+11Hz -0.026369 -0.00897071
+ 2.214e+11Hz -0.0263873 -0.00894483
+ 2.215e+11Hz -0.0264056 -0.00891869
+ 2.216e+11Hz -0.0264238 -0.00889229
+ 2.217e+11Hz -0.026442 -0.00886562
+ 2.218e+11Hz -0.0264602 -0.00883869
+ 2.219e+11Hz -0.0264783 -0.0088115
+ 2.22e+11Hz -0.0264964 -0.00878404
+ 2.221e+11Hz -0.0265144 -0.00875631
+ 2.222e+11Hz -0.0265324 -0.00872832
+ 2.223e+11Hz -0.0265503 -0.00870006
+ 2.224e+11Hz -0.0265682 -0.00867153
+ 2.225e+11Hz -0.0265859 -0.00864274
+ 2.226e+11Hz -0.0266036 -0.00861367
+ 2.227e+11Hz -0.0266213 -0.00858434
+ 2.228e+11Hz -0.0266388 -0.00855473
+ 2.229e+11Hz -0.0266563 -0.00852486
+ 2.23e+11Hz -0.0266736 -0.00849471
+ 2.231e+11Hz -0.0266909 -0.0084643
+ 2.232e+11Hz -0.0267081 -0.00843362
+ 2.233e+11Hz -0.0267251 -0.00840266
+ 2.234e+11Hz -0.0267421 -0.00837144
+ 2.235e+11Hz -0.0267589 -0.00833994
+ 2.236e+11Hz -0.0267757 -0.00830818
+ 2.237e+11Hz -0.0267923 -0.00827615
+ 2.238e+11Hz -0.0268087 -0.00824385
+ 2.239e+11Hz -0.0268251 -0.00821128
+ 2.24e+11Hz -0.0268413 -0.00817845
+ 2.241e+11Hz -0.0268574 -0.00814535
+ 2.242e+11Hz -0.0268733 -0.00811198
+ 2.243e+11Hz -0.0268891 -0.00807835
+ 2.244e+11Hz -0.0269047 -0.00804445
+ 2.245e+11Hz -0.0269202 -0.00801029
+ 2.246e+11Hz -0.0269355 -0.00797587
+ 2.247e+11Hz -0.0269507 -0.00794119
+ 2.248e+11Hz -0.0269657 -0.00790625
+ 2.249e+11Hz -0.0269805 -0.00787105
+ 2.25e+11Hz -0.0269951 -0.00783559
+ 2.251e+11Hz -0.0270096 -0.00779987
+ 2.252e+11Hz -0.0270238 -0.00776391
+ 2.253e+11Hz -0.0270379 -0.00772769
+ 2.254e+11Hz -0.0270518 -0.00769121
+ 2.255e+11Hz -0.0270655 -0.00765449
+ 2.256e+11Hz -0.027079 -0.00761752
+ 2.257e+11Hz -0.0270922 -0.00758031
+ 2.258e+11Hz -0.0271053 -0.00754285
+ 2.259e+11Hz -0.0271182 -0.00750515
+ 2.26e+11Hz -0.0271308 -0.00746721
+ 2.261e+11Hz -0.0271432 -0.00742904
+ 2.262e+11Hz -0.0271554 -0.00739062
+ 2.263e+11Hz -0.0271673 -0.00735198
+ 2.264e+11Hz -0.027179 -0.0073131
+ 2.265e+11Hz -0.0271905 -0.007274
+ 2.266e+11Hz -0.0272017 -0.00723467
+ 2.267e+11Hz -0.0272127 -0.00719512
+ 2.268e+11Hz -0.0272234 -0.00715534
+ 2.269e+11Hz -0.0272339 -0.00711535
+ 2.27e+11Hz -0.0272441 -0.00707515
+ 2.271e+11Hz -0.027254 -0.00703473
+ 2.272e+11Hz -0.0272637 -0.0069941
+ 2.273e+11Hz -0.0272731 -0.00695327
+ 2.274e+11Hz -0.0272823 -0.00691223
+ 2.275e+11Hz -0.0272911 -0.00687099
+ 2.276e+11Hz -0.0272997 -0.00682956
+ 2.277e+11Hz -0.027308 -0.00678793
+ 2.278e+11Hz -0.027316 -0.00674611
+ 2.279e+11Hz -0.0273237 -0.00670411
+ 2.28e+11Hz -0.0273311 -0.00666192
+ 2.281e+11Hz -0.0273383 -0.00661955
+ 2.282e+11Hz -0.0273451 -0.00657701
+ 2.283e+11Hz -0.0273516 -0.00653429
+ 2.284e+11Hz -0.0273578 -0.0064914
+ 2.285e+11Hz -0.0273637 -0.00644835
+ 2.286e+11Hz -0.0273693 -0.00640514
+ 2.287e+11Hz -0.0273746 -0.00636176
+ 2.288e+11Hz -0.0273795 -0.00631824
+ 2.289e+11Hz -0.0273841 -0.00627456
+ 2.29e+11Hz -0.0273884 -0.00623074
+ 2.291e+11Hz -0.0273924 -0.00618678
+ 2.292e+11Hz -0.0273961 -0.00614267
+ 2.293e+11Hz -0.0273994 -0.00609844
+ 2.294e+11Hz -0.0274024 -0.00605407
+ 2.295e+11Hz -0.027405 -0.00600958
+ 2.296e+11Hz -0.0274073 -0.00596497
+ 2.297e+11Hz -0.0274092 -0.00592024
+ 2.298e+11Hz -0.0274109 -0.0058754
+ 2.299e+11Hz -0.0274121 -0.00583045
+ 2.3e+11Hz -0.027413 -0.00578539
+ 2.301e+11Hz -0.0274136 -0.00574024
+ 2.302e+11Hz -0.0274138 -0.00569499
+ 2.303e+11Hz -0.0274137 -0.00564965
+ 2.304e+11Hz -0.0274131 -0.00560423
+ 2.305e+11Hz -0.0274123 -0.00555873
+ 2.306e+11Hz -0.0274111 -0.00551315
+ 2.307e+11Hz -0.0274095 -0.0054675
+ 2.308e+11Hz -0.0274075 -0.00542178
+ 2.309e+11Hz -0.0274052 -0.005376
+ 2.31e+11Hz -0.0274025 -0.00533016
+ 2.311e+11Hz -0.0273995 -0.00528427
+ 2.312e+11Hz -0.0273961 -0.00523833
+ 2.313e+11Hz -0.0273923 -0.00519235
+ 2.314e+11Hz -0.0273881 -0.00514633
+ 2.315e+11Hz -0.0273836 -0.00510028
+ 2.316e+11Hz -0.0273787 -0.0050542
+ 2.317e+11Hz -0.0273734 -0.0050081
+ 2.318e+11Hz -0.0273678 -0.00496198
+ 2.319e+11Hz -0.0273617 -0.00491584
+ 2.32e+11Hz -0.0273553 -0.0048697
+ 2.321e+11Hz -0.0273485 -0.00482355
+ 2.322e+11Hz -0.0273414 -0.00477741
+ 2.323e+11Hz -0.0273339 -0.00473127
+ 2.324e+11Hz -0.0273259 -0.00468514
+ 2.325e+11Hz -0.0273177 -0.00463904
+ 2.326e+11Hz -0.027309 -0.00459295
+ 2.327e+11Hz -0.0272999 -0.00454689
+ 2.328e+11Hz -0.0272905 -0.00450086
+ 2.329e+11Hz -0.0272807 -0.00445486
+ 2.33e+11Hz -0.0272705 -0.00440891
+ 2.331e+11Hz -0.02726 -0.00436301
+ 2.332e+11Hz -0.027249 -0.00431716
+ 2.333e+11Hz -0.0272377 -0.00427136
+ 2.334e+11Hz -0.0272261 -0.00422563
+ 2.335e+11Hz -0.027214 -0.00417996
+ 2.336e+11Hz -0.0272016 -0.00413437
+ 2.337e+11Hz -0.0271888 -0.00408885
+ 2.338e+11Hz -0.0271756 -0.00404342
+ 2.339e+11Hz -0.027162 -0.00399807
+ 2.34e+11Hz -0.0271481 -0.00395281
+ 2.341e+11Hz -0.0271338 -0.00390765
+ 2.342e+11Hz -0.0271191 -0.00386259
+ 2.343e+11Hz -0.0271041 -0.00381764
+ 2.344e+11Hz -0.0270887 -0.00377279
+ 2.345e+11Hz -0.027073 -0.00372807
+ 2.346e+11Hz -0.0270568 -0.00368346
+ 2.347e+11Hz -0.0270404 -0.00363898
+ 2.348e+11Hz -0.0270235 -0.00359464
+ 2.349e+11Hz -0.0270063 -0.00355042
+ 2.35e+11Hz -0.0269888 -0.00350635
+ 2.351e+11Hz -0.0269709 -0.00346242
+ 2.352e+11Hz -0.0269526 -0.00341864
+ 2.353e+11Hz -0.026934 -0.00337501
+ 2.354e+11Hz -0.026915 -0.00333154
+ 2.355e+11Hz -0.0268957 -0.00328823
+ 2.356e+11Hz -0.0268761 -0.00324509
+ 2.357e+11Hz -0.0268561 -0.00320213
+ 2.358e+11Hz -0.0268357 -0.00315934
+ 2.359e+11Hz -0.0268151 -0.00311673
+ 2.36e+11Hz -0.0267941 -0.0030743
+ 2.361e+11Hz -0.0267727 -0.00303206
+ 2.362e+11Hz -0.0267511 -0.00299002
+ 2.363e+11Hz -0.0267291 -0.00294817
+ 2.364e+11Hz -0.0267068 -0.00290653
+ 2.365e+11Hz -0.0266842 -0.00286509
+ 2.366e+11Hz -0.0266612 -0.00282386
+ 2.367e+11Hz -0.026638 -0.00278284
+ 2.368e+11Hz -0.0266144 -0.00274204
+ 2.369e+11Hz -0.0265905 -0.00270146
+ 2.37e+11Hz -0.0265663 -0.00266111
+ 2.371e+11Hz -0.0265418 -0.00262099
+ 2.372e+11Hz -0.026517 -0.0025811
+ 2.373e+11Hz -0.026492 -0.00254144
+ 2.374e+11Hz -0.0264666 -0.00250203
+ 2.375e+11Hz -0.0264409 -0.00246286
+ 2.376e+11Hz -0.026415 -0.00242394
+ 2.377e+11Hz -0.0263888 -0.00238526
+ 2.378e+11Hz -0.0263623 -0.00234684
+ 2.379e+11Hz -0.0263355 -0.00230868
+ 2.38e+11Hz -0.0263084 -0.00227078
+ 2.381e+11Hz -0.0262811 -0.00223314
+ 2.382e+11Hz -0.0262535 -0.00219577
+ 2.383e+11Hz -0.0262257 -0.00215867
+ 2.384e+11Hz -0.0261976 -0.00212184
+ 2.385e+11Hz -0.0261693 -0.00208528
+ 2.386e+11Hz -0.0261407 -0.00204901
+ 2.387e+11Hz -0.0261119 -0.00201301
+ 2.388e+11Hz -0.0260828 -0.0019773
+ 2.389e+11Hz -0.0260535 -0.00194187
+ 2.39e+11Hz -0.0260239 -0.00190674
+ 2.391e+11Hz -0.0259942 -0.00187189
+ 2.392e+11Hz -0.0259642 -0.00183734
+ 2.393e+11Hz -0.025934 -0.00180309
+ 2.394e+11Hz -0.0259036 -0.00176913
+ 2.395e+11Hz -0.0258729 -0.00173548
+ 2.396e+11Hz -0.0258421 -0.00170213
+ 2.397e+11Hz -0.0258111 -0.00166908
+ 2.398e+11Hz -0.0257798 -0.00163634
+ 2.399e+11Hz -0.0257484 -0.0016039
+ 2.4e+11Hz -0.0257168 -0.00157178
+ 2.401e+11Hz -0.025685 -0.00153997
+ 2.402e+11Hz -0.025653 -0.00150848
+ 2.403e+11Hz -0.0256209 -0.0014773
+ 2.404e+11Hz -0.0255886 -0.00144644
+ 2.405e+11Hz -0.0255561 -0.00141589
+ 2.406e+11Hz -0.0255234 -0.00138567
+ 2.407e+11Hz -0.0254906 -0.00135577
+ 2.408e+11Hz -0.0254577 -0.00132619
+ 2.409e+11Hz -0.0254246 -0.00129693
+ 2.41e+11Hz -0.0253913 -0.001268
+ 2.411e+11Hz -0.0253579 -0.0012394
+ 2.412e+11Hz -0.0253244 -0.00121112
+ 2.413e+11Hz -0.0252908 -0.00118317
+ 2.414e+11Hz -0.025257 -0.00115555
+ 2.415e+11Hz -0.0252231 -0.00112826
+ 2.416e+11Hz -0.0251891 -0.00110129
+ 2.417e+11Hz -0.025155 -0.00107466
+ 2.418e+11Hz -0.0251207 -0.00104836
+ 2.419e+11Hz -0.0250864 -0.00102239
+ 2.42e+11Hz -0.025052 -0.000996754
+ 2.421e+11Hz -0.0250174 -0.000971449
+ 2.422e+11Hz -0.0249828 -0.000946475
+ 2.423e+11Hz -0.0249481 -0.000921835
+ 2.424e+11Hz -0.0249134 -0.000897527
+ 2.425e+11Hz -0.0248785 -0.000873551
+ 2.426e+11Hz -0.0248436 -0.000849908
+ 2.427e+11Hz -0.0248086 -0.000826598
+ 2.428e+11Hz -0.0247735 -0.000803619
+ 2.429e+11Hz -0.0247384 -0.000780973
+ 2.43e+11Hz -0.0247033 -0.000758658
+ 2.431e+11Hz -0.0246681 -0.000736674
+ 2.432e+11Hz -0.0246328 -0.000715021
+ 2.433e+11Hz -0.0245975 -0.000693698
+ 2.434e+11Hz -0.0245622 -0.000672704
+ 2.435e+11Hz -0.0245268 -0.000652039
+ 2.436e+11Hz -0.0244914 -0.000631703
+ 2.437e+11Hz -0.024456 -0.000611694
+ 2.438e+11Hz -0.0244206 -0.000592011
+ 2.439e+11Hz -0.0243851 -0.000572654
+ 2.44e+11Hz -0.0243497 -0.000553621
+ 2.441e+11Hz -0.0243142 -0.000534912
+ 2.442e+11Hz -0.0242788 -0.000516525
+ 2.443e+11Hz -0.0242433 -0.000498459
+ 2.444e+11Hz -0.0242078 -0.000480714
+ 2.445e+11Hz -0.0241724 -0.000463287
+ 2.446e+11Hz -0.024137 -0.000446178
+ 2.447e+11Hz -0.0241015 -0.000429384
+ 2.448e+11Hz -0.0240662 -0.000412905
+ 2.449e+11Hz -0.0240308 -0.00039674
+ 2.45e+11Hz -0.0239955 -0.000380885
+ 2.451e+11Hz -0.0239601 -0.000365341
+ 2.452e+11Hz -0.0239249 -0.000350105
+ 2.453e+11Hz -0.0238897 -0.000335176
+ 2.454e+11Hz -0.0238545 -0.000320551
+ 2.455e+11Hz -0.0238193 -0.000306229
+ 2.456e+11Hz -0.0237843 -0.000292209
+ 2.457e+11Hz -0.0237492 -0.000278487
+ 2.458e+11Hz -0.0237143 -0.000265063
+ 2.459e+11Hz -0.0236794 -0.000251935
+ 2.46e+11Hz -0.0236445 -0.000239099
+ 2.461e+11Hz -0.0236097 -0.000226555
+ 2.462e+11Hz -0.023575 -0.0002143
+ 2.463e+11Hz -0.0235404 -0.000202332
+ 2.464e+11Hz -0.0235059 -0.000190649
+ 2.465e+11Hz -0.0234714 -0.000179248
+ 2.466e+11Hz -0.023437 -0.000168128
+ 2.467e+11Hz -0.0234027 -0.000157285
+ 2.468e+11Hz -0.0233685 -0.000146718
+ 2.469e+11Hz -0.0233344 -0.000136425
+ 2.47e+11Hz -0.0233004 -0.000126402
+ 2.471e+11Hz -0.0232665 -0.000116648
+ 2.472e+11Hz -0.0232327 -0.00010716
+ 2.473e+11Hz -0.023199 -9.7935e-05
+ 2.474e+11Hz -0.0231654 -8.89712e-05
+ 2.475e+11Hz -0.023132 -8.02658e-05
+ 2.476e+11Hz -0.0230986 -7.18163e-05
+ 2.477e+11Hz -0.0230653 -6.36199e-05
+ 2.478e+11Hz -0.0230322 -5.56742e-05
+ 2.479e+11Hz -0.0229992 -4.79764e-05
+ 2.48e+11Hz -0.0229663 -4.05238e-05
+ 2.481e+11Hz -0.0229336 -3.33139e-05
+ 2.482e+11Hz -0.0229009 -2.63438e-05
+ 2.483e+11Hz -0.0228684 -1.96108e-05
+ 2.484e+11Hz -0.0228361 -1.31123e-05
+ 2.485e+11Hz -0.0228038 -6.84528e-06
+ 2.486e+11Hz -0.0227717 -8.0713e-07
+ 2.487e+11Hz -0.0227398 5.005e-06
+ 2.488e+11Hz -0.022708 1.05939e-05
+ 2.489e+11Hz -0.0226763 1.59625e-05
+ 2.49e+11Hz -0.0226448 2.11135e-05
+ 2.491e+11Hz -0.0226134 2.60498e-05
+ 2.492e+11Hz -0.0225822 3.07743e-05
+ 2.493e+11Hz -0.0225511 3.52899e-05
+ 2.494e+11Hz -0.0225202 3.95994e-05
+ 2.495e+11Hz -0.0224894 4.37058e-05
+ 2.496e+11Hz -0.0224588 4.76118e-05
+ 2.497e+11Hz -0.0224284 5.13205e-05
+ 2.498e+11Hz -0.0223981 5.48347e-05
+ 2.499e+11Hz -0.0223679 5.81574e-05
+ 2.5e+11Hz -0.022338 6.12915e-05
+ 2.501e+11Hz -0.0223082 6.42398e-05
+ 2.502e+11Hz -0.0222785 6.70053e-05
+ 2.503e+11Hz -0.022249 6.9591e-05
+ 2.504e+11Hz -0.0222197 7.19997e-05
+ 2.505e+11Hz -0.0221906 7.42343e-05
+ 2.506e+11Hz -0.0221616 7.62979e-05
+ 2.507e+11Hz -0.0221328 7.81932e-05
+ 2.508e+11Hz -0.0221042 7.99233e-05
+ 2.509e+11Hz -0.0220758 8.1491e-05
+ 2.51e+11Hz -0.0220475 8.28993e-05
+ 2.511e+11Hz -0.0220194 8.4151e-05
+ 2.512e+11Hz -0.0219915 8.52491e-05
+ 2.513e+11Hz -0.0219637 8.61964e-05
+ 2.514e+11Hz -0.0219362 8.69958e-05
+ 2.515e+11Hz -0.0219088 8.76503e-05
+ 2.516e+11Hz -0.0218816 8.81626e-05
+ 2.517e+11Hz -0.0218545 8.85356e-05
+ 2.518e+11Hz -0.0218277 8.87723e-05
+ 2.519e+11Hz -0.021801 8.88754e-05
+ 2.52e+11Hz -0.0217745 8.88478e-05
+ 2.521e+11Hz -0.0217482 8.86923e-05
+ 2.522e+11Hz -0.0217221 8.84117e-05
+ 2.523e+11Hz -0.0216962 8.80088e-05
+ 2.524e+11Hz -0.0216704 8.74864e-05
+ 2.525e+11Hz -0.0216449 8.68474e-05
+ 2.526e+11Hz -0.0216195 8.60944e-05
+ 2.527e+11Hz -0.0215943 8.52302e-05
+ 2.528e+11Hz -0.0215693 8.42576e-05
+ 2.529e+11Hz -0.0215445 8.31793e-05
+ 2.53e+11Hz -0.0215198 8.1998e-05
+ 2.531e+11Hz -0.0214954 8.07164e-05
+ 2.532e+11Hz -0.0214711 7.93372e-05
+ 2.533e+11Hz -0.0214471 7.78631e-05
+ 2.534e+11Hz -0.0214232 7.62967e-05
+ 2.535e+11Hz -0.0213995 7.46407e-05
+ 2.536e+11Hz -0.021376 7.28978e-05
+ 2.537e+11Hz -0.0213526 7.10704e-05
+ 2.538e+11Hz -0.0213295 6.91612e-05
+ 2.539e+11Hz -0.0213066 6.71729e-05
+ 2.54e+11Hz -0.0212838 6.5108e-05
+ 2.541e+11Hz -0.0212612 6.29689e-05
+ 2.542e+11Hz -0.0212389 6.07584e-05
+ 2.543e+11Hz -0.0212167 5.84788e-05
+ 2.544e+11Hz -0.0211947 5.61327e-05
+ 2.545e+11Hz -0.0211728 5.37226e-05
+ 2.546e+11Hz -0.0211512 5.1251e-05
+ 2.547e+11Hz -0.0211298 4.87203e-05
+ 2.548e+11Hz -0.0211085 4.61329e-05
+ 2.549e+11Hz -0.0210874 4.34914e-05
+ 2.55e+11Hz -0.0210665 4.0798e-05
+ 2.551e+11Hz -0.0210458 3.80552e-05
+ 2.552e+11Hz -0.0210253 3.52655e-05
+ 2.553e+11Hz -0.021005 3.2431e-05
+ 2.554e+11Hz -0.0209849 2.95543e-05
+ 2.555e+11Hz -0.0209649 2.66376e-05
+ 2.556e+11Hz -0.0209451 2.36832e-05
+ 2.557e+11Hz -0.0209255 2.06935e-05
+ 2.558e+11Hz -0.0209061 1.76707e-05
+ 2.559e+11Hz -0.0208869 1.46172e-05
+ 2.56e+11Hz -0.0208679 1.15352e-05
+ 2.561e+11Hz -0.020849 8.42689e-06
+ 2.562e+11Hz -0.0208303 5.29458e-06
+ 2.563e+11Hz -0.0208119 2.14047e-06
+ 2.564e+11Hz -0.0207935 -1.03323e-06
+ 2.565e+11Hz -0.0207754 -4.22433e-06
+ 2.566e+11Hz -0.0207575 -7.43064e-06
+ 2.567e+11Hz -0.0207397 -1.065e-05
+ 2.568e+11Hz -0.0207221 -1.38802e-05
+ 2.569e+11Hz -0.0207047 -1.71192e-05
+ 2.57e+11Hz -0.0206875 -2.03647e-05
+ 2.571e+11Hz -0.0206704 -2.36147e-05
+ 2.572e+11Hz -0.0206535 -2.68671e-05
+ 2.573e+11Hz -0.0206368 -3.01198e-05
+ 2.574e+11Hz -0.0206203 -3.33706e-05
+ 2.575e+11Hz -0.020604 -3.66174e-05
+ 2.576e+11Hz -0.0205878 -3.98583e-05
+ 2.577e+11Hz -0.0205718 -4.30911e-05
+ 2.578e+11Hz -0.020556 -4.63138e-05
+ 2.579e+11Hz -0.0205403 -4.95243e-05
+ 2.58e+11Hz -0.0205248 -5.27206e-05
+ 2.581e+11Hz -0.0205095 -5.59006e-05
+ 2.582e+11Hz -0.0204944 -5.90624e-05
+ 2.583e+11Hz -0.0204794 -6.22039e-05
+ 2.584e+11Hz -0.0204646 -6.53231e-05
+ 2.585e+11Hz -0.02045 -6.8418e-05
+ 2.586e+11Hz -0.0204355 -7.14866e-05
+ 2.587e+11Hz -0.0204212 -7.45269e-05
+ 2.588e+11Hz -0.0204071 -7.75369e-05
+ 2.589e+11Hz -0.0203931 -8.05147e-05
+ 2.59e+11Hz -0.0203793 -8.34582e-05
+ 2.591e+11Hz -0.0203657 -8.63655e-05
+ 2.592e+11Hz -0.0203522 -8.92346e-05
+ 2.593e+11Hz -0.0203389 -9.20635e-05
+ 2.594e+11Hz -0.0203258 -9.48504e-05
+ 2.595e+11Hz -0.0203128 -9.75931e-05
+ 2.596e+11Hz -0.0203 -0.00010029
+ 2.597e+11Hz -0.0202874 -0.000102939
+ 2.598e+11Hz -0.0202749 -0.000105537
+ 2.599e+11Hz -0.0202625 -0.000108084
+ 2.6e+11Hz -0.0202503 -0.000110577
+ 2.601e+11Hz -0.0202383 -0.000113014
+ 2.602e+11Hz -0.0202264 -0.000115394
+ 2.603e+11Hz -0.0202147 -0.000117713
+ 2.604e+11Hz -0.0202032 -0.000119971
+ 2.605e+11Hz -0.0201917 -0.000122166
+ 2.606e+11Hz -0.0201805 -0.000124295
+ 2.607e+11Hz -0.0201694 -0.000126356
+ 2.608e+11Hz -0.0201584 -0.000128348
+ 2.609e+11Hz -0.0201476 -0.000130269
+ 2.61e+11Hz -0.020137 -0.000132116
+ 2.611e+11Hz -0.0201265 -0.000133888
+ 2.612e+11Hz -0.0201161 -0.000135583
+ 2.613e+11Hz -0.0201059 -0.000137198
+ 2.614e+11Hz -0.0200958 -0.000138732
+ 2.615e+11Hz -0.0200859 -0.000140183
+ 2.616e+11Hz -0.0200761 -0.00014155
+ 2.617e+11Hz -0.0200664 -0.000142829
+ 2.618e+11Hz -0.0200569 -0.000144019
+ 2.619e+11Hz -0.0200476 -0.000145118
+ 2.62e+11Hz -0.0200383 -0.000146124
+ 2.621e+11Hz -0.0200292 -0.000147035
+ 2.622e+11Hz -0.0200203 -0.000147849
+ 2.623e+11Hz -0.0200115 -0.000148565
+ 2.624e+11Hz -0.0200028 -0.000149179
+ 2.625e+11Hz -0.0199942 -0.000149691
+ 2.626e+11Hz -0.0199858 -0.000150098
+ 2.627e+11Hz -0.0199775 -0.000150399
+ 2.628e+11Hz -0.0199693 -0.00015059
+ 2.629e+11Hz -0.0199613 -0.000150671
+ 2.63e+11Hz -0.0199534 -0.00015064
+ 2.631e+11Hz -0.0199456 -0.000150493
+ 2.632e+11Hz -0.0199379 -0.00015023
+ 2.633e+11Hz -0.0199303 -0.000149848
+ 2.634e+11Hz -0.0199229 -0.000149346
+ 2.635e+11Hz -0.0199156 -0.000148721
+ 2.636e+11Hz -0.0199084 -0.000147972
+ 2.637e+11Hz -0.0199013 -0.000147096
+ 2.638e+11Hz -0.0198943 -0.000146091
+ 2.639e+11Hz -0.0198875 -0.000144956
+ 2.64e+11Hz -0.0198807 -0.000143689
+ 2.641e+11Hz -0.0198741 -0.000142287
+ 2.642e+11Hz -0.0198676 -0.000140749
+ 2.643e+11Hz -0.0198611 -0.000139072
+ 2.644e+11Hz -0.0198548 -0.000137255
+ 2.645e+11Hz -0.0198486 -0.000135296
+ 2.646e+11Hz -0.0198425 -0.000133192
+ 2.647e+11Hz -0.0198364 -0.000130943
+ 2.648e+11Hz -0.0198305 -0.000128545
+ 2.649e+11Hz -0.0198247 -0.000125997
+ 2.65e+11Hz -0.0198189 -0.000123297
+ 2.651e+11Hz -0.0198133 -0.000120444
+ 2.652e+11Hz -0.0198077 -0.000117434
+ 2.653e+11Hz -0.0198022 -0.000114267
+ 2.654e+11Hz -0.0197968 -0.00011094
+ 2.655e+11Hz -0.0197915 -0.000107452
+ 2.656e+11Hz -0.0197863 -0.0001038
+ 2.657e+11Hz -0.0197811 -9.99837e-05
+ 2.658e+11Hz -0.019776 -9.59999e-05
+ 2.659e+11Hz -0.019771 -9.18472e-05
+ 2.66e+11Hz -0.0197661 -8.75239e-05
+ 2.661e+11Hz -0.0197612 -8.30281e-05
+ 2.662e+11Hz -0.0197564 -7.83581e-05
+ 2.663e+11Hz -0.0197517 -7.3512e-05
+ 2.664e+11Hz -0.019747 -6.84882e-05
+ 2.665e+11Hz -0.0197424 -6.32849e-05
+ 2.666e+11Hz -0.0197378 -5.79003e-05
+ 2.667e+11Hz -0.0197333 -5.23329e-05
+ 2.668e+11Hz -0.0197288 -4.65809e-05
+ 2.669e+11Hz -0.0197244 -4.06428e-05
+ 2.67e+11Hz -0.01972 -3.45167e-05
+ 2.671e+11Hz -0.0197157 -2.82013e-05
+ 2.672e+11Hz -0.0197114 -2.16949e-05
+ 2.673e+11Hz -0.0197072 -1.49959e-05
+ 2.674e+11Hz -0.0197029 -8.10288e-06
+ 2.675e+11Hz -0.0196988 -1.0143e-06
+ 2.676e+11Hz -0.0196946 6.27128e-06
+ 2.677e+11Hz -0.0196905 1.37553e-05
+ 2.678e+11Hz -0.0196863 2.14392e-05
+ 2.679e+11Hz -0.0196822 2.93242e-05
+ 2.68e+11Hz -0.0196782 3.74118e-05
+ 2.681e+11Hz -0.0196741 4.57032e-05
+ 2.682e+11Hz -0.01967 5.41997e-05
+ 2.683e+11Hz -0.019666 6.29025e-05
+ 2.684e+11Hz -0.0196619 7.18128e-05
+ 2.685e+11Hz -0.0196579 8.09317e-05
+ 2.686e+11Hz -0.0196538 9.02604e-05
+ 2.687e+11Hz -0.0196498 9.97999e-05
+ 2.688e+11Hz -0.0196457 0.000109551
+ 2.689e+11Hz -0.0196416 0.000119515
+ 2.69e+11Hz -0.0196375 0.000129693
+ 2.691e+11Hz -0.0196334 0.000140086
+ 2.692e+11Hz -0.0196292 0.000150694
+ 2.693e+11Hz -0.019625 0.000161518
+ 2.694e+11Hz -0.0196208 0.000172559
+ 2.695e+11Hz -0.0196166 0.000183818
+ 2.696e+11Hz -0.0196123 0.000195295
+ 2.697e+11Hz -0.019608 0.000206992
+ 2.698e+11Hz -0.0196036 0.000218907
+ 2.699e+11Hz -0.0195992 0.000231043
+ 2.7e+11Hz -0.0195947 0.000243399
+ 2.701e+11Hz -0.0195901 0.000255975
+ 2.702e+11Hz -0.0195855 0.000268773
+ 2.703e+11Hz -0.0195808 0.000281792
+ 2.704e+11Hz -0.0195761 0.000295032
+ 2.705e+11Hz -0.0195713 0.000308494
+ 2.706e+11Hz -0.0195664 0.000322178
+ 2.707e+11Hz -0.0195614 0.000336083
+ 2.708e+11Hz -0.0195563 0.00035021
+ 2.709e+11Hz -0.0195511 0.000364558
+ 2.71e+11Hz -0.0195459 0.000379128
+ 2.711e+11Hz -0.0195405 0.000393918
+ 2.712e+11Hz -0.0195351 0.00040893
+ 2.713e+11Hz -0.0195295 0.000424161
+ 2.714e+11Hz -0.0195238 0.000439612
+ 2.715e+11Hz -0.019518 0.000455283
+ 2.716e+11Hz -0.0195121 0.000471172
+ 2.717e+11Hz -0.019506 0.000487279
+ 2.718e+11Hz -0.0194999 0.000503603
+ 2.719e+11Hz -0.0194936 0.000520144
+ 2.72e+11Hz -0.0194871 0.000536899
+ 2.721e+11Hz -0.0194805 0.00055387
+ 2.722e+11Hz -0.0194738 0.000571054
+ 2.723e+11Hz -0.0194669 0.000588449
+ 2.724e+11Hz -0.0194599 0.000606056
+ 2.725e+11Hz -0.0194527 0.000623873
+ 2.726e+11Hz -0.0194453 0.000641898
+ 2.727e+11Hz -0.0194378 0.00066013
+ 2.728e+11Hz -0.01943 0.000678567
+ 2.729e+11Hz -0.0194222 0.000697208
+ 2.73e+11Hz -0.0194141 0.00071605
+ 2.731e+11Hz -0.0194058 0.000735093
+ 2.732e+11Hz -0.0193974 0.000754334
+ 2.733e+11Hz -0.0193888 0.000773772
+ 2.734e+11Hz -0.0193799 0.000793404
+ 2.735e+11Hz -0.0193709 0.000813228
+ 2.736e+11Hz -0.0193616 0.000833242
+ 2.737e+11Hz -0.0193522 0.000853444
+ 2.738e+11Hz -0.0193425 0.000873831
+ 2.739e+11Hz -0.0193326 0.000894401
+ 2.74e+11Hz -0.0193225 0.000915151
+ 2.741e+11Hz -0.0193121 0.000936079
+ 2.742e+11Hz -0.0193016 0.000957182
+ 2.743e+11Hz -0.0192907 0.000978457
+ 2.744e+11Hz -0.0192797 0.000999901
+ 2.745e+11Hz -0.0192684 0.00102151
+ 2.746e+11Hz -0.0192568 0.00104328
+ 2.747e+11Hz -0.019245 0.00106522
+ 2.748e+11Hz -0.0192329 0.00108731
+ 2.749e+11Hz -0.0192206 0.00110955
+ 2.75e+11Hz -0.019208 0.00113195
+ 2.751e+11Hz -0.0191951 0.00115449
+ 2.752e+11Hz -0.019182 0.00117717
+ 2.753e+11Hz -0.0191686 0.0012
+ 2.754e+11Hz -0.0191549 0.00122295
+ 2.755e+11Hz -0.0191409 0.00124604
+ 2.756e+11Hz -0.0191266 0.00126926
+ 2.757e+11Hz -0.0191121 0.00129261
+ 2.758e+11Hz -0.0190972 0.00131607
+ 2.759e+11Hz -0.0190821 0.00133965
+ 2.76e+11Hz -0.0190666 0.00136333
+ 2.761e+11Hz -0.0190509 0.00138713
+ 2.762e+11Hz -0.0190348 0.00141103
+ 2.763e+11Hz -0.0190184 0.00143503
+ 2.764e+11Hz -0.0190017 0.00145912
+ 2.765e+11Hz -0.0189847 0.0014833
+ 2.766e+11Hz -0.0189674 0.00150756
+ 2.767e+11Hz -0.0189497 0.00153191
+ 2.768e+11Hz -0.0189317 0.00155633
+ 2.769e+11Hz -0.0189134 0.00158082
+ 2.77e+11Hz -0.0188947 0.00160537
+ 2.771e+11Hz -0.0188757 0.00162998
+ 2.772e+11Hz -0.0188564 0.00165465
+ 2.773e+11Hz -0.0188367 0.00167937
+ 2.774e+11Hz -0.0188167 0.00170413
+ 2.775e+11Hz -0.0187964 0.00172893
+ 2.776e+11Hz -0.0187757 0.00175376
+ 2.777e+11Hz -0.0187546 0.00177862
+ 2.778e+11Hz -0.0187332 0.00180351
+ 2.779e+11Hz -0.0187114 0.00182841
+ 2.78e+11Hz -0.0186893 0.00185332
+ 2.781e+11Hz -0.0186668 0.00187824
+ 2.782e+11Hz -0.018644 0.00190316
+ 2.783e+11Hz -0.0186208 0.00192807
+ 2.784e+11Hz -0.0185972 0.00195297
+ 2.785e+11Hz -0.0185733 0.00197785
+ 2.786e+11Hz -0.018549 0.00200271
+ 2.787e+11Hz -0.0185243 0.00202753
+ 2.788e+11Hz -0.0184993 0.00205232
+ 2.789e+11Hz -0.0184739 0.00207707
+ 2.79e+11Hz -0.0184482 0.00210178
+ 2.791e+11Hz -0.018422 0.00212642
+ 2.792e+11Hz -0.0183955 0.00215101
+ 2.793e+11Hz -0.0183686 0.00217553
+ 2.794e+11Hz -0.0183414 0.00219998
+ 2.795e+11Hz -0.0183137 0.00222435
+ 2.796e+11Hz -0.0182857 0.00224863
+ 2.797e+11Hz -0.0182574 0.00227282
+ 2.798e+11Hz -0.0182286 0.00229692
+ 2.799e+11Hz -0.0181995 0.0023209
+ 2.8e+11Hz -0.01817 0.00234478
+ 2.801e+11Hz -0.0181401 0.00236854
+ 2.802e+11Hz -0.0181099 0.00239218
+ 2.803e+11Hz -0.0180793 0.00241568
+ 2.804e+11Hz -0.0180483 0.00243905
+ 2.805e+11Hz -0.018017 0.00246227
+ 2.806e+11Hz -0.0179852 0.00248535
+ 2.807e+11Hz -0.0179531 0.00250826
+ 2.808e+11Hz -0.0179207 0.00253102
+ 2.809e+11Hz -0.0178879 0.00255361
+ 2.81e+11Hz -0.0178547 0.00257602
+ 2.811e+11Hz -0.0178211 0.00259824
+ 2.812e+11Hz -0.0177872 0.00262028
+ 2.813e+11Hz -0.017753 0.00264213
+ 2.814e+11Hz -0.0177183 0.00266377
+ 2.815e+11Hz -0.0176833 0.0026852
+ 2.816e+11Hz -0.017648 0.00270642
+ 2.817e+11Hz -0.0176123 0.00272742
+ 2.818e+11Hz -0.0175763 0.00274819
+ 2.819e+11Hz -0.0175399 0.00276873
+ 2.82e+11Hz -0.0175032 0.00278903
+ 2.821e+11Hz -0.0174661 0.00280908
+ 2.822e+11Hz -0.0174287 0.00282888
+ 2.823e+11Hz -0.017391 0.00284842
+ 2.824e+11Hz -0.0173529 0.00286769
+ 2.825e+11Hz -0.0173146 0.0028867
+ 2.826e+11Hz -0.0172758 0.00290543
+ 2.827e+11Hz -0.0172368 0.00292387
+ 2.828e+11Hz -0.0171975 0.00294203
+ 2.829e+11Hz -0.0171578 0.00295989
+ 2.83e+11Hz -0.0171178 0.00297745
+ 2.831e+11Hz -0.0170775 0.00299471
+ 2.832e+11Hz -0.0170369 0.00301165
+ 2.833e+11Hz -0.0169961 0.00302828
+ 2.834e+11Hz -0.0169549 0.00304458
+ 2.835e+11Hz -0.0169134 0.00306056
+ 2.836e+11Hz -0.0168717 0.0030762
+ 2.837e+11Hz -0.0168297 0.0030915
+ 2.838e+11Hz -0.0167874 0.00310645
+ 2.839e+11Hz -0.0167448 0.00312106
+ 2.84e+11Hz -0.016702 0.00313531
+ 2.841e+11Hz -0.0166589 0.0031492
+ 2.842e+11Hz -0.0166156 0.00316272
+ 2.843e+11Hz -0.016572 0.00317587
+ 2.844e+11Hz -0.0165281 0.00318865
+ 2.845e+11Hz -0.0164841 0.00320105
+ 2.846e+11Hz -0.0164398 0.00321307
+ 2.847e+11Hz -0.0163952 0.0032247
+ 2.848e+11Hz -0.0163505 0.00323593
+ 2.849e+11Hz -0.0163055 0.00324677
+ 2.85e+11Hz -0.0162604 0.0032572
+ 2.851e+11Hz -0.016215 0.00326723
+ 2.852e+11Hz -0.0161694 0.00327685
+ 2.853e+11Hz -0.0161237 0.00328606
+ 2.854e+11Hz -0.0160777 0.00329485
+ 2.855e+11Hz -0.0160316 0.00330322
+ 2.856e+11Hz -0.0159853 0.00331116
+ 2.857e+11Hz -0.0159389 0.00331868
+ 2.858e+11Hz -0.0158923 0.00332577
+ 2.859e+11Hz -0.0158455 0.00333242
+ 2.86e+11Hz -0.0157986 0.00333863
+ 2.861e+11Hz -0.0157516 0.00334441
+ 2.862e+11Hz -0.0157044 0.00334974
+ 2.863e+11Hz -0.0156571 0.00335463
+ 2.864e+11Hz -0.0156097 0.00335906
+ 2.865e+11Hz -0.0155622 0.00336305
+ 2.866e+11Hz -0.0155146 0.00336659
+ 2.867e+11Hz -0.0154669 0.00336967
+ 2.868e+11Hz -0.0154191 0.00337229
+ 2.869e+11Hz -0.0153712 0.00337446
+ 2.87e+11Hz -0.0153233 0.00337616
+ 2.871e+11Hz -0.0152753 0.00337741
+ 2.872e+11Hz -0.0152272 0.00337819
+ 2.873e+11Hz -0.0151791 0.0033785
+ 2.874e+11Hz -0.0151309 0.00337835
+ 2.875e+11Hz -0.0150827 0.00337774
+ 2.876e+11Hz -0.0150345 0.00337665
+ 2.877e+11Hz -0.0149863 0.0033751
+ 2.878e+11Hz -0.014938 0.00337308
+ 2.879e+11Hz -0.0148898 0.00337059
+ 2.88e+11Hz -0.0148415 0.00336763
+ 2.881e+11Hz -0.0147933 0.0033642
+ 2.882e+11Hz -0.0147451 0.0033603
+ 2.883e+11Hz -0.0146969 0.00335593
+ 2.884e+11Hz -0.0146487 0.00335109
+ 2.885e+11Hz -0.0146006 0.00334578
+ 2.886e+11Hz -0.0145525 0.00334001
+ 2.887e+11Hz -0.0145045 0.00333376
+ 2.888e+11Hz -0.0144566 0.00332705
+ 2.889e+11Hz -0.0144087 0.00331988
+ 2.89e+11Hz -0.0143609 0.00331224
+ 2.891e+11Hz -0.0143132 0.00330414
+ 2.892e+11Hz -0.0142656 0.00329557
+ 2.893e+11Hz -0.0142181 0.00328655
+ 2.894e+11Hz -0.0141707 0.00327707
+ 2.895e+11Hz -0.0141234 0.00326713
+ 2.896e+11Hz -0.0140763 0.00325674
+ 2.897e+11Hz -0.0140293 0.0032459
+ 2.898e+11Hz -0.0139824 0.00323461
+ 2.899e+11Hz -0.0139357 0.00322287
+ 2.9e+11Hz -0.0138891 0.00321068
+ 2.901e+11Hz -0.0138427 0.00319805
+ 2.902e+11Hz -0.0137964 0.00318499
+ 2.903e+11Hz -0.0137504 0.00317149
+ 2.904e+11Hz -0.0137045 0.00315756
+ 2.905e+11Hz -0.0136588 0.0031432
+ 2.906e+11Hz -0.0136133 0.00312841
+ 2.907e+11Hz -0.013568 0.0031132
+ 2.908e+11Hz -0.0135229 0.00309757
+ 2.909e+11Hz -0.013478 0.00308153
+ 2.91e+11Hz -0.0134334 0.00306507
+ 2.911e+11Hz -0.013389 0.00304821
+ 2.912e+11Hz -0.0133448 0.00303095
+ 2.913e+11Hz -0.0133009 0.00301329
+ 2.914e+11Hz -0.0132572 0.00299524
+ 2.915e+11Hz -0.0132138 0.0029768
+ 2.916e+11Hz -0.0131706 0.00295797
+ 2.917e+11Hz -0.0131277 0.00293877
+ 2.918e+11Hz -0.0130851 0.00291919
+ 2.919e+11Hz -0.0130427 0.00289924
+ 2.92e+11Hz -0.0130007 0.00287893
+ 2.921e+11Hz -0.0129589 0.00285826
+ 2.922e+11Hz -0.0129174 0.00283723
+ 2.923e+11Hz -0.0128763 0.00281586
+ 2.924e+11Hz -0.0128354 0.00279415
+ 2.925e+11Hz -0.0127949 0.0027721
+ 2.926e+11Hz -0.0127546 0.00274972
+ 2.927e+11Hz -0.0127147 0.00272701
+ 2.928e+11Hz -0.0126751 0.00270398
+ 2.929e+11Hz -0.0126359 0.00268065
+ 2.93e+11Hz -0.012597 0.002657
+ 2.931e+11Hz -0.0125584 0.00263305
+ 2.932e+11Hz -0.0125202 0.00260882
+ 2.933e+11Hz -0.0124823 0.00258429
+ 2.934e+11Hz -0.0124448 0.00255948
+ 2.935e+11Hz -0.0124076 0.0025344
+ 2.936e+11Hz -0.0123708 0.00250904
+ 2.937e+11Hz -0.0123344 0.00248343
+ 2.938e+11Hz -0.0122983 0.00245756
+ 2.939e+11Hz -0.0122626 0.00243145
+ 2.94e+11Hz -0.0122273 0.00240509
+ 2.941e+11Hz -0.0121923 0.0023785
+ 2.942e+11Hz -0.0121578 0.00235168
+ 2.943e+11Hz -0.0121236 0.00232464
+ 2.944e+11Hz -0.0120898 0.00229738
+ 2.945e+11Hz -0.0120564 0.00226993
+ 2.946e+11Hz -0.0120234 0.00224227
+ 2.947e+11Hz -0.0119908 0.00221442
+ 2.948e+11Hz -0.0119585 0.00218638
+ 2.949e+11Hz -0.0119267 0.00215817
+ 2.95e+11Hz -0.0118953 0.00212979
+ 2.951e+11Hz -0.0118642 0.00210124
+ 2.952e+11Hz -0.0118336 0.00207254
+ 2.953e+11Hz -0.0118034 0.00204369
+ 2.954e+11Hz -0.0117736 0.0020147
+ 2.955e+11Hz -0.0117442 0.00198558
+ 2.956e+11Hz -0.0117152 0.00195633
+ 2.957e+11Hz -0.0116866 0.00192696
+ 2.958e+11Hz -0.0116584 0.00189747
+ 2.959e+11Hz -0.0116306 0.00186789
+ 2.96e+11Hz -0.0116033 0.0018382
+ 2.961e+11Hz -0.0115763 0.00180843
+ 2.962e+11Hz -0.0115498 0.00177858
+ 2.963e+11Hz -0.0115237 0.00174865
+ 2.964e+11Hz -0.0114979 0.00171865
+ 2.965e+11Hz -0.0114726 0.00168859
+ 2.966e+11Hz -0.0114477 0.00165848
+ 2.967e+11Hz -0.0114232 0.00162832
+ 2.968e+11Hz -0.0113991 0.00159812
+ 2.969e+11Hz -0.0113754 0.00156789
+ 2.97e+11Hz -0.0113522 0.00153764
+ 2.971e+11Hz -0.0113293 0.00150737
+ 2.972e+11Hz -0.0113068 0.00147708
+ 2.973e+11Hz -0.0112848 0.0014468
+ 2.974e+11Hz -0.0112631 0.00141651
+ 2.975e+11Hz -0.0112418 0.00138624
+ 2.976e+11Hz -0.0112209 0.00135598
+ 2.977e+11Hz -0.0112004 0.00132575
+ 2.978e+11Hz -0.0111804 0.00129555
+ 2.979e+11Hz -0.0111607 0.00126538
+ 2.98e+11Hz -0.0111413 0.00123526
+ 2.981e+11Hz -0.0111224 0.00120519
+ 2.982e+11Hz -0.0111039 0.00117517
+ 2.983e+11Hz -0.0110857 0.00114522
+ 2.984e+11Hz -0.0110679 0.00111534
+ 2.985e+11Hz -0.0110505 0.00108553
+ 2.986e+11Hz -0.0110334 0.0010558
+ 2.987e+11Hz -0.0110167 0.00102616
+ 2.988e+11Hz -0.0110004 0.000996611
+ 2.989e+11Hz -0.0109844 0.000967163
+ 2.99e+11Hz -0.0109688 0.000937819
+ 2.991e+11Hz -0.0109536 0.000908586
+ 2.992e+11Hz -0.0109387 0.000879469
+ 2.993e+11Hz -0.0109241 0.000850473
+ 2.994e+11Hz -0.0109099 0.000821604
+ 2.995e+11Hz -0.010896 0.000792867
+ 2.996e+11Hz -0.0108824 0.000764267
+ 2.997e+11Hz -0.0108692 0.00073581
+ 2.998e+11Hz -0.0108563 0.000707499
+ 2.999e+11Hz -0.0108437 0.000679341
+ 3e+11Hz -0.0108314 0.00065134
+ ]

A12 %vd(20 3) %vd(12, 3) xfer2
.model xfer2 xfer R_I=true table=[
+ 0Hz 0.995436 0
+ 1e+08Hz 0.995435 -0.000814178
+ 2e+08Hz 0.995433 -0.00162834
+ 3e+08Hz 0.99543 -0.00244247
+ 4e+08Hz 0.995425 -0.00325656
+ 5e+08Hz 0.99542 -0.00407058
+ 6e+08Hz 0.995412 -0.00488452
+ 7e+08Hz 0.995404 -0.00569837
+ 8e+08Hz 0.995394 -0.00651211
+ 9e+08Hz 0.995383 -0.00732573
+ 1e+09Hz 0.995371 -0.0081392
+ 1.1e+09Hz 0.995358 -0.00895252
+ 1.2e+09Hz 0.995343 -0.00976567
+ 1.3e+09Hz 0.995327 -0.0105786
+ 1.4e+09Hz 0.99531 -0.0113914
+ 1.5e+09Hz 0.995291 -0.012204
+ 1.6e+09Hz 0.995271 -0.0130163
+ 1.7e+09Hz 0.99525 -0.0138284
+ 1.8e+09Hz 0.995228 -0.0146402
+ 1.9e+09Hz 0.995204 -0.0154517
+ 2e+09Hz 0.99518 -0.016263
+ 2.1e+09Hz 0.995154 -0.017074
+ 2.2e+09Hz 0.995126 -0.0178846
+ 2.3e+09Hz 0.995098 -0.0186949
+ 2.4e+09Hz 0.995068 -0.0195049
+ 2.5e+09Hz 0.995038 -0.0203146
+ 2.6e+09Hz 0.995006 -0.0211238
+ 2.7e+09Hz 0.994973 -0.0219327
+ 2.8e+09Hz 0.994938 -0.0227412
+ 2.9e+09Hz 0.994903 -0.0235493
+ 3e+09Hz 0.994866 -0.024357
+ 3.1e+09Hz 0.994829 -0.0251643
+ 3.2e+09Hz 0.99479 -0.0259711
+ 3.3e+09Hz 0.99475 -0.0267775
+ 3.4e+09Hz 0.994709 -0.0275834
+ 3.5e+09Hz 0.994667 -0.0283889
+ 3.6e+09Hz 0.994624 -0.0291939
+ 3.7e+09Hz 0.994579 -0.0299984
+ 3.8e+09Hz 0.994534 -0.0308024
+ 3.9e+09Hz 0.994488 -0.031606
+ 4e+09Hz 0.994441 -0.032409
+ 4.1e+09Hz 0.994392 -0.0332114
+ 4.2e+09Hz 0.994343 -0.0340134
+ 4.3e+09Hz 0.994292 -0.0348148
+ 4.4e+09Hz 0.994241 -0.0356157
+ 4.5e+09Hz 0.994189 -0.036416
+ 4.6e+09Hz 0.994136 -0.0372158
+ 4.7e+09Hz 0.994081 -0.038015
+ 4.8e+09Hz 0.994026 -0.0388137
+ 4.9e+09Hz 0.99397 -0.0396118
+ 5e+09Hz 0.993913 -0.0404093
+ 5.1e+09Hz 0.993856 -0.0412062
+ 5.2e+09Hz 0.993797 -0.0420026
+ 5.3e+09Hz 0.993737 -0.0427983
+ 5.4e+09Hz 0.993677 -0.0435935
+ 5.5e+09Hz 0.993616 -0.044388
+ 5.6e+09Hz 0.993554 -0.045182
+ 5.7e+09Hz 0.993491 -0.0459753
+ 5.8e+09Hz 0.993427 -0.0467681
+ 5.9e+09Hz 0.993363 -0.0475602
+ 6e+09Hz 0.993298 -0.0483518
+ 6.1e+09Hz 0.993232 -0.0491427
+ 6.2e+09Hz 0.993165 -0.049933
+ 6.3e+09Hz 0.993098 -0.0507227
+ 6.4e+09Hz 0.99303 -0.0515118
+ 6.5e+09Hz 0.992961 -0.0523003
+ 6.6e+09Hz 0.992892 -0.0530882
+ 6.7e+09Hz 0.992821 -0.0538755
+ 6.8e+09Hz 0.992751 -0.0546622
+ 6.9e+09Hz 0.992679 -0.0554482
+ 7e+09Hz 0.992607 -0.0562337
+ 7.1e+09Hz 0.992535 -0.0570185
+ 7.2e+09Hz 0.992461 -0.0578028
+ 7.3e+09Hz 0.992387 -0.0585865
+ 7.4e+09Hz 0.992313 -0.0593695
+ 7.5e+09Hz 0.992238 -0.060152
+ 7.6e+09Hz 0.992162 -0.0609339
+ 7.7e+09Hz 0.992086 -0.0617152
+ 7.8e+09Hz 0.99201 -0.062496
+ 7.9e+09Hz 0.991933 -0.0632762
+ 8e+09Hz 0.991855 -0.0640558
+ 8.1e+09Hz 0.991777 -0.0648348
+ 8.2e+09Hz 0.991698 -0.0656133
+ 8.3e+09Hz 0.991619 -0.0663912
+ 8.4e+09Hz 0.99154 -0.0671686
+ 8.5e+09Hz 0.991459 -0.0679455
+ 8.6e+09Hz 0.991379 -0.0687218
+ 8.7e+09Hz 0.991298 -0.0694976
+ 8.8e+09Hz 0.991217 -0.0702728
+ 8.9e+09Hz 0.991135 -0.0710476
+ 9e+09Hz 0.991053 -0.0718218
+ 9.1e+09Hz 0.99097 -0.0725956
+ 9.2e+09Hz 0.990888 -0.0733689
+ 9.3e+09Hz 0.990804 -0.0741417
+ 9.4e+09Hz 0.990721 -0.074914
+ 9.5e+09Hz 0.990637 -0.0756858
+ 9.6e+09Hz 0.990552 -0.0764572
+ 9.7e+09Hz 0.990467 -0.0772282
+ 9.8e+09Hz 0.990382 -0.0779987
+ 9.9e+09Hz 0.990297 -0.0787687
+ 1e+10Hz 0.990211 -0.0795384
+ 1.01e+10Hz 0.990125 -0.0803076
+ 1.02e+10Hz 0.990039 -0.0810764
+ 1.03e+10Hz 0.989952 -0.0818449
+ 1.04e+10Hz 0.989865 -0.0826129
+ 1.05e+10Hz 0.989778 -0.0833806
+ 1.06e+10Hz 0.98969 -0.0841479
+ 1.07e+10Hz 0.989603 -0.0849148
+ 1.08e+10Hz 0.989514 -0.0856814
+ 1.09e+10Hz 0.989426 -0.0864477
+ 1.1e+10Hz 0.989337 -0.0872136
+ 1.11e+10Hz 0.989248 -0.0879793
+ 1.12e+10Hz 0.989159 -0.0887446
+ 1.13e+10Hz 0.98907 -0.0895096
+ 1.14e+10Hz 0.98898 -0.0902743
+ 1.15e+10Hz 0.98889 -0.0910387
+ 1.16e+10Hz 0.9888 -0.0918029
+ 1.17e+10Hz 0.988709 -0.0925668
+ 1.18e+10Hz 0.988618 -0.0933304
+ 1.19e+10Hz 0.988527 -0.0940938
+ 1.2e+10Hz 0.988436 -0.094857
+ 1.21e+10Hz 0.988344 -0.09562
+ 1.22e+10Hz 0.988253 -0.0963827
+ 1.23e+10Hz 0.988161 -0.0971453
+ 1.24e+10Hz 0.988068 -0.0979076
+ 1.25e+10Hz 0.987976 -0.0986698
+ 1.26e+10Hz 0.987883 -0.0994318
+ 1.27e+10Hz 0.98779 -0.100194
+ 1.28e+10Hz 0.987697 -0.100955
+ 1.29e+10Hz 0.987603 -0.101717
+ 1.3e+10Hz 0.987509 -0.102478
+ 1.31e+10Hz 0.987415 -0.10324
+ 1.32e+10Hz 0.987321 -0.104001
+ 1.33e+10Hz 0.987226 -0.104762
+ 1.34e+10Hz 0.987131 -0.105523
+ 1.35e+10Hz 0.987036 -0.106283
+ 1.36e+10Hz 0.986941 -0.107044
+ 1.37e+10Hz 0.986845 -0.107805
+ 1.38e+10Hz 0.986749 -0.108566
+ 1.39e+10Hz 0.986653 -0.109326
+ 1.4e+10Hz 0.986556 -0.110087
+ 1.41e+10Hz 0.986459 -0.110847
+ 1.42e+10Hz 0.986362 -0.111607
+ 1.43e+10Hz 0.986265 -0.112368
+ 1.44e+10Hz 0.986167 -0.113128
+ 1.45e+10Hz 0.986069 -0.113888
+ 1.46e+10Hz 0.985971 -0.114649
+ 1.47e+10Hz 0.985872 -0.115409
+ 1.48e+10Hz 0.985773 -0.116169
+ 1.49e+10Hz 0.985673 -0.11693
+ 1.5e+10Hz 0.985574 -0.11769
+ 1.51e+10Hz 0.985474 -0.11845
+ 1.52e+10Hz 0.985373 -0.119211
+ 1.53e+10Hz 0.985273 -0.119971
+ 1.54e+10Hz 0.985172 -0.120732
+ 1.55e+10Hz 0.98507 -0.121492
+ 1.56e+10Hz 0.984968 -0.122253
+ 1.57e+10Hz 0.984866 -0.123013
+ 1.58e+10Hz 0.984763 -0.123774
+ 1.59e+10Hz 0.98466 -0.124535
+ 1.6e+10Hz 0.984557 -0.125295
+ 1.61e+10Hz 0.984453 -0.126056
+ 1.62e+10Hz 0.984349 -0.126817
+ 1.63e+10Hz 0.984244 -0.127578
+ 1.64e+10Hz 0.984139 -0.128339
+ 1.65e+10Hz 0.984034 -0.1291
+ 1.66e+10Hz 0.983928 -0.129861
+ 1.67e+10Hz 0.983822 -0.130623
+ 1.68e+10Hz 0.983715 -0.131384
+ 1.69e+10Hz 0.983607 -0.132145
+ 1.7e+10Hz 0.9835 -0.132907
+ 1.71e+10Hz 0.983391 -0.133669
+ 1.72e+10Hz 0.983283 -0.13443
+ 1.73e+10Hz 0.983174 -0.135192
+ 1.74e+10Hz 0.983064 -0.135954
+ 1.75e+10Hz 0.982954 -0.136716
+ 1.76e+10Hz 0.982843 -0.137478
+ 1.77e+10Hz 0.982732 -0.13824
+ 1.78e+10Hz 0.98262 -0.139002
+ 1.79e+10Hz 0.982508 -0.139765
+ 1.8e+10Hz 0.982395 -0.140527
+ 1.81e+10Hz 0.982281 -0.14129
+ 1.82e+10Hz 0.982167 -0.142052
+ 1.83e+10Hz 0.982053 -0.142815
+ 1.84e+10Hz 0.981938 -0.143578
+ 1.85e+10Hz 0.981822 -0.14434
+ 1.86e+10Hz 0.981706 -0.145103
+ 1.87e+10Hz 0.981589 -0.145866
+ 1.88e+10Hz 0.981472 -0.146629
+ 1.89e+10Hz 0.981354 -0.147393
+ 1.9e+10Hz 0.981235 -0.148156
+ 1.91e+10Hz 0.981116 -0.148919
+ 1.92e+10Hz 0.980996 -0.149682
+ 1.93e+10Hz 0.980876 -0.150446
+ 1.94e+10Hz 0.980754 -0.151209
+ 1.95e+10Hz 0.980633 -0.151973
+ 1.96e+10Hz 0.98051 -0.152736
+ 1.97e+10Hz 0.980387 -0.1535
+ 1.98e+10Hz 0.980264 -0.154264
+ 1.99e+10Hz 0.980139 -0.155027
+ 2e+10Hz 0.980014 -0.155791
+ 2.01e+10Hz 0.979889 -0.156555
+ 2.02e+10Hz 0.979762 -0.157319
+ 2.03e+10Hz 0.979635 -0.158083
+ 2.04e+10Hz 0.979508 -0.158846
+ 2.05e+10Hz 0.979379 -0.15961
+ 2.06e+10Hz 0.97925 -0.160374
+ 2.07e+10Hz 0.979121 -0.161138
+ 2.08e+10Hz 0.97899 -0.161902
+ 2.09e+10Hz 0.978859 -0.162666
+ 2.1e+10Hz 0.978727 -0.16343
+ 2.11e+10Hz 0.978595 -0.164193
+ 2.12e+10Hz 0.978461 -0.164957
+ 2.13e+10Hz 0.978327 -0.165721
+ 2.14e+10Hz 0.978193 -0.166485
+ 2.15e+10Hz 0.978057 -0.167249
+ 2.16e+10Hz 0.977921 -0.168012
+ 2.17e+10Hz 0.977785 -0.168776
+ 2.18e+10Hz 0.977647 -0.169539
+ 2.19e+10Hz 0.977509 -0.170303
+ 2.2e+10Hz 0.97737 -0.171066
+ 2.21e+10Hz 0.97723 -0.17183
+ 2.22e+10Hz 0.97709 -0.172593
+ 2.23e+10Hz 0.976948 -0.173356
+ 2.24e+10Hz 0.976807 -0.174119
+ 2.25e+10Hz 0.976664 -0.174882
+ 2.26e+10Hz 0.976521 -0.175645
+ 2.27e+10Hz 0.976377 -0.176408
+ 2.28e+10Hz 0.976232 -0.17717
+ 2.29e+10Hz 0.976086 -0.177933
+ 2.3e+10Hz 0.97594 -0.178695
+ 2.31e+10Hz 0.975793 -0.179458
+ 2.32e+10Hz 0.975645 -0.18022
+ 2.33e+10Hz 0.975497 -0.180982
+ 2.34e+10Hz 0.975348 -0.181743
+ 2.35e+10Hz 0.975198 -0.182505
+ 2.36e+10Hz 0.975047 -0.183267
+ 2.37e+10Hz 0.974896 -0.184028
+ 2.38e+10Hz 0.974744 -0.184789
+ 2.39e+10Hz 0.974591 -0.18555
+ 2.4e+10Hz 0.974438 -0.186311
+ 2.41e+10Hz 0.974284 -0.187072
+ 2.42e+10Hz 0.974129 -0.187832
+ 2.43e+10Hz 0.973973 -0.188592
+ 2.44e+10Hz 0.973817 -0.189352
+ 2.45e+10Hz 0.97366 -0.190112
+ 2.46e+10Hz 0.973502 -0.190872
+ 2.47e+10Hz 0.973344 -0.191631
+ 2.48e+10Hz 0.973185 -0.19239
+ 2.49e+10Hz 0.973025 -0.193149
+ 2.5e+10Hz 0.972864 -0.193908
+ 2.51e+10Hz 0.972703 -0.194667
+ 2.52e+10Hz 0.972541 -0.195425
+ 2.53e+10Hz 0.972379 -0.196183
+ 2.54e+10Hz 0.972216 -0.196941
+ 2.55e+10Hz 0.972052 -0.197698
+ 2.56e+10Hz 0.971887 -0.198455
+ 2.57e+10Hz 0.971722 -0.199212
+ 2.58e+10Hz 0.971556 -0.199969
+ 2.59e+10Hz 0.97139 -0.200726
+ 2.6e+10Hz 0.971223 -0.201482
+ 2.61e+10Hz 0.971055 -0.202238
+ 2.62e+10Hz 0.970886 -0.202994
+ 2.63e+10Hz 0.970717 -0.203749
+ 2.64e+10Hz 0.970548 -0.204504
+ 2.65e+10Hz 0.970377 -0.205259
+ 2.66e+10Hz 0.970206 -0.206014
+ 2.67e+10Hz 0.970035 -0.206768
+ 2.68e+10Hz 0.969863 -0.207522
+ 2.69e+10Hz 0.96969 -0.208276
+ 2.7e+10Hz 0.969516 -0.209029
+ 2.71e+10Hz 0.969342 -0.209782
+ 2.72e+10Hz 0.969168 -0.210535
+ 2.73e+10Hz 0.968993 -0.211288
+ 2.74e+10Hz 0.968817 -0.21204
+ 2.75e+10Hz 0.968641 -0.212792
+ 2.76e+10Hz 0.968464 -0.213544
+ 2.77e+10Hz 0.968286 -0.214296
+ 2.78e+10Hz 0.968108 -0.215047
+ 2.79e+10Hz 0.96793 -0.215798
+ 2.8e+10Hz 0.96775 -0.216548
+ 2.81e+10Hz 0.967571 -0.217298
+ 2.82e+10Hz 0.96739 -0.218048
+ 2.83e+10Hz 0.96721 -0.218798
+ 2.84e+10Hz 0.967028 -0.219548
+ 2.85e+10Hz 0.966846 -0.220297
+ 2.86e+10Hz 0.966664 -0.221046
+ 2.87e+10Hz 0.966481 -0.221794
+ 2.88e+10Hz 0.966298 -0.222542
+ 2.89e+10Hz 0.966114 -0.22329
+ 2.9e+10Hz 0.965929 -0.224038
+ 2.91e+10Hz 0.965744 -0.224785
+ 2.92e+10Hz 0.965559 -0.225533
+ 2.93e+10Hz 0.965373 -0.22628
+ 2.94e+10Hz 0.965186 -0.227026
+ 2.95e+10Hz 0.964999 -0.227772
+ 2.96e+10Hz 0.964812 -0.228519
+ 2.97e+10Hz 0.964624 -0.229264
+ 2.98e+10Hz 0.964435 -0.23001
+ 2.99e+10Hz 0.964246 -0.230755
+ 3e+10Hz 0.964057 -0.2315
+ 3.01e+10Hz 0.963867 -0.232245
+ 3.02e+10Hz 0.963677 -0.232989
+ 3.03e+10Hz 0.963486 -0.233734
+ 3.04e+10Hz 0.963295 -0.234478
+ 3.05e+10Hz 0.963103 -0.235221
+ 3.06e+10Hz 0.962911 -0.235965
+ 3.07e+10Hz 0.962718 -0.236708
+ 3.08e+10Hz 0.962525 -0.237451
+ 3.09e+10Hz 0.962332 -0.238194
+ 3.1e+10Hz 0.962138 -0.238936
+ 3.11e+10Hz 0.961943 -0.239679
+ 3.12e+10Hz 0.961748 -0.240421
+ 3.13e+10Hz 0.961553 -0.241163
+ 3.14e+10Hz 0.961357 -0.241905
+ 3.15e+10Hz 0.961161 -0.242646
+ 3.16e+10Hz 0.960964 -0.243387
+ 3.17e+10Hz 0.960767 -0.244128
+ 3.18e+10Hz 0.96057 -0.244869
+ 3.19e+10Hz 0.960372 -0.24561
+ 3.2e+10Hz 0.960174 -0.24635
+ 3.21e+10Hz 0.959975 -0.247091
+ 3.22e+10Hz 0.959775 -0.247831
+ 3.23e+10Hz 0.959576 -0.248571
+ 3.24e+10Hz 0.959376 -0.24931
+ 3.25e+10Hz 0.959175 -0.25005
+ 3.26e+10Hz 0.958974 -0.250789
+ 3.27e+10Hz 0.958773 -0.251528
+ 3.28e+10Hz 0.958571 -0.252267
+ 3.29e+10Hz 0.958369 -0.253006
+ 3.3e+10Hz 0.958166 -0.253745
+ 3.31e+10Hz 0.957963 -0.254484
+ 3.32e+10Hz 0.95776 -0.255222
+ 3.33e+10Hz 0.957556 -0.25596
+ 3.34e+10Hz 0.957351 -0.256698
+ 3.35e+10Hz 0.957146 -0.257436
+ 3.36e+10Hz 0.956941 -0.258174
+ 3.37e+10Hz 0.956735 -0.258912
+ 3.38e+10Hz 0.956529 -0.25965
+ 3.39e+10Hz 0.956323 -0.260387
+ 3.4e+10Hz 0.956116 -0.261125
+ 3.41e+10Hz 0.955908 -0.261862
+ 3.42e+10Hz 0.9557 -0.262599
+ 3.43e+10Hz 0.955492 -0.263336
+ 3.44e+10Hz 0.955283 -0.264073
+ 3.45e+10Hz 0.955074 -0.26481
+ 3.46e+10Hz 0.954864 -0.265546
+ 3.47e+10Hz 0.954654 -0.266283
+ 3.48e+10Hz 0.954443 -0.26702
+ 3.49e+10Hz 0.954232 -0.267756
+ 3.5e+10Hz 0.954021 -0.268492
+ 3.51e+10Hz 0.953809 -0.269228
+ 3.52e+10Hz 0.953596 -0.269965
+ 3.53e+10Hz 0.953383 -0.270701
+ 3.54e+10Hz 0.95317 -0.271437
+ 3.55e+10Hz 0.952956 -0.272173
+ 3.56e+10Hz 0.952742 -0.272908
+ 3.57e+10Hz 0.952527 -0.273644
+ 3.58e+10Hz 0.952312 -0.27438
+ 3.59e+10Hz 0.952096 -0.275115
+ 3.6e+10Hz 0.951879 -0.275851
+ 3.61e+10Hz 0.951663 -0.276586
+ 3.62e+10Hz 0.951445 -0.277322
+ 3.63e+10Hz 0.951227 -0.278057
+ 3.64e+10Hz 0.951009 -0.278792
+ 3.65e+10Hz 0.95079 -0.279528
+ 3.66e+10Hz 0.950571 -0.280263
+ 3.67e+10Hz 0.950351 -0.280998
+ 3.68e+10Hz 0.950131 -0.281733
+ 3.69e+10Hz 0.94991 -0.282468
+ 3.7e+10Hz 0.949689 -0.283203
+ 3.71e+10Hz 0.949467 -0.283938
+ 3.72e+10Hz 0.949244 -0.284672
+ 3.73e+10Hz 0.949021 -0.285407
+ 3.74e+10Hz 0.948798 -0.286142
+ 3.75e+10Hz 0.948574 -0.286876
+ 3.76e+10Hz 0.948349 -0.287611
+ 3.77e+10Hz 0.948124 -0.288345
+ 3.78e+10Hz 0.947898 -0.28908
+ 3.79e+10Hz 0.947672 -0.289814
+ 3.8e+10Hz 0.947445 -0.290549
+ 3.81e+10Hz 0.947218 -0.291283
+ 3.82e+10Hz 0.94699 -0.292017
+ 3.83e+10Hz 0.946761 -0.292751
+ 3.84e+10Hz 0.946532 -0.293485
+ 3.85e+10Hz 0.946302 -0.294219
+ 3.86e+10Hz 0.946072 -0.294953
+ 3.87e+10Hz 0.945841 -0.295687
+ 3.88e+10Hz 0.94561 -0.296421
+ 3.89e+10Hz 0.945377 -0.297154
+ 3.9e+10Hz 0.945145 -0.297888
+ 3.91e+10Hz 0.944912 -0.298622
+ 3.92e+10Hz 0.944678 -0.299355
+ 3.93e+10Hz 0.944443 -0.300088
+ 3.94e+10Hz 0.944208 -0.300822
+ 3.95e+10Hz 0.943972 -0.301555
+ 3.96e+10Hz 0.943736 -0.302288
+ 3.97e+10Hz 0.943499 -0.303021
+ 3.98e+10Hz 0.943262 -0.303754
+ 3.99e+10Hz 0.943023 -0.304487
+ 4e+10Hz 0.942785 -0.30522
+ 4.01e+10Hz 0.942545 -0.305953
+ 4.02e+10Hz 0.942305 -0.306685
+ 4.03e+10Hz 0.942065 -0.307418
+ 4.04e+10Hz 0.941823 -0.30815
+ 4.05e+10Hz 0.941581 -0.308882
+ 4.06e+10Hz 0.941339 -0.309615
+ 4.07e+10Hz 0.941095 -0.310347
+ 4.08e+10Hz 0.940851 -0.311079
+ 4.09e+10Hz 0.940607 -0.31181
+ 4.1e+10Hz 0.940362 -0.312542
+ 4.11e+10Hz 0.940116 -0.313274
+ 4.12e+10Hz 0.939869 -0.314005
+ 4.13e+10Hz 0.939622 -0.314736
+ 4.14e+10Hz 0.939374 -0.315468
+ 4.15e+10Hz 0.939126 -0.316199
+ 4.16e+10Hz 0.938877 -0.316929
+ 4.17e+10Hz 0.938627 -0.31766
+ 4.18e+10Hz 0.938377 -0.318391
+ 4.19e+10Hz 0.938126 -0.319121
+ 4.2e+10Hz 0.937874 -0.319851
+ 4.21e+10Hz 0.937621 -0.320581
+ 4.22e+10Hz 0.937368 -0.321311
+ 4.23e+10Hz 0.937114 -0.322041
+ 4.24e+10Hz 0.93686 -0.322771
+ 4.25e+10Hz 0.936605 -0.3235
+ 4.26e+10Hz 0.936349 -0.324229
+ 4.27e+10Hz 0.936093 -0.324958
+ 4.28e+10Hz 0.935836 -0.325687
+ 4.29e+10Hz 0.935578 -0.326416
+ 4.3e+10Hz 0.935319 -0.327144
+ 4.31e+10Hz 0.93506 -0.327872
+ 4.32e+10Hz 0.934801 -0.328601
+ 4.33e+10Hz 0.93454 -0.329328
+ 4.34e+10Hz 0.934279 -0.330056
+ 4.35e+10Hz 0.934017 -0.330783
+ 4.36e+10Hz 0.933755 -0.331511
+ 4.37e+10Hz 0.933492 -0.332238
+ 4.38e+10Hz 0.933228 -0.332964
+ 4.39e+10Hz 0.932964 -0.333691
+ 4.4e+10Hz 0.932698 -0.334417
+ 4.41e+10Hz 0.932433 -0.335143
+ 4.42e+10Hz 0.932166 -0.335869
+ 4.43e+10Hz 0.931899 -0.336594
+ 4.44e+10Hz 0.931632 -0.33732
+ 4.45e+10Hz 0.931363 -0.338045
+ 4.46e+10Hz 0.931094 -0.338769
+ 4.47e+10Hz 0.930825 -0.339494
+ 4.48e+10Hz 0.930554 -0.340218
+ 4.49e+10Hz 0.930283 -0.340942
+ 4.5e+10Hz 0.930012 -0.341666
+ 4.51e+10Hz 0.929739 -0.342389
+ 4.52e+10Hz 0.929467 -0.343113
+ 4.53e+10Hz 0.929193 -0.343836
+ 4.54e+10Hz 0.928919 -0.344558
+ 4.55e+10Hz 0.928644 -0.345281
+ 4.56e+10Hz 0.928369 -0.346003
+ 4.57e+10Hz 0.928093 -0.346724
+ 4.58e+10Hz 0.927816 -0.347446
+ 4.59e+10Hz 0.927539 -0.348167
+ 4.6e+10Hz 0.927261 -0.348888
+ 4.61e+10Hz 0.926982 -0.349609
+ 4.62e+10Hz 0.926703 -0.350329
+ 4.63e+10Hz 0.926423 -0.351049
+ 4.64e+10Hz 0.926143 -0.351769
+ 4.65e+10Hz 0.925862 -0.352488
+ 4.66e+10Hz 0.92558 -0.353207
+ 4.67e+10Hz 0.925298 -0.353926
+ 4.68e+10Hz 0.925015 -0.354644
+ 4.69e+10Hz 0.924732 -0.355362
+ 4.7e+10Hz 0.924448 -0.35608
+ 4.71e+10Hz 0.924163 -0.356798
+ 4.72e+10Hz 0.923878 -0.357515
+ 4.73e+10Hz 0.923592 -0.358232
+ 4.74e+10Hz 0.923306 -0.358949
+ 4.75e+10Hz 0.923019 -0.359665
+ 4.76e+10Hz 0.922732 -0.360381
+ 4.77e+10Hz 0.922444 -0.361096
+ 4.78e+10Hz 0.922155 -0.361812
+ 4.79e+10Hz 0.921866 -0.362527
+ 4.8e+10Hz 0.921576 -0.363241
+ 4.81e+10Hz 0.921286 -0.363955
+ 4.82e+10Hz 0.920995 -0.364669
+ 4.83e+10Hz 0.920704 -0.365383
+ 4.84e+10Hz 0.920412 -0.366096
+ 4.85e+10Hz 0.920119 -0.366809
+ 4.86e+10Hz 0.919826 -0.367522
+ 4.87e+10Hz 0.919532 -0.368234
+ 4.88e+10Hz 0.919238 -0.368946
+ 4.89e+10Hz 0.918944 -0.369658
+ 4.9e+10Hz 0.918649 -0.37037
+ 4.91e+10Hz 0.918353 -0.371081
+ 4.92e+10Hz 0.918057 -0.371791
+ 4.93e+10Hz 0.91776 -0.372502
+ 4.94e+10Hz 0.917463 -0.373212
+ 4.95e+10Hz 0.917165 -0.373922
+ 4.96e+10Hz 0.916866 -0.374631
+ 4.97e+10Hz 0.916568 -0.37534
+ 4.98e+10Hz 0.916268 -0.376049
+ 4.99e+10Hz 0.915969 -0.376757
+ 5e+10Hz 0.915668 -0.377465
+ 5.01e+10Hz 0.915367 -0.378173
+ 5.02e+10Hz 0.915066 -0.378881
+ 5.03e+10Hz 0.914764 -0.379588
+ 5.04e+10Hz 0.914462 -0.380295
+ 5.05e+10Hz 0.914159 -0.381002
+ 5.06e+10Hz 0.913856 -0.381708
+ 5.07e+10Hz 0.913552 -0.382414
+ 5.08e+10Hz 0.913248 -0.383119
+ 5.09e+10Hz 0.912943 -0.383825
+ 5.1e+10Hz 0.912638 -0.38453
+ 5.11e+10Hz 0.912332 -0.385234
+ 5.12e+10Hz 0.912026 -0.385939
+ 5.13e+10Hz 0.91172 -0.386643
+ 5.14e+10Hz 0.911412 -0.387347
+ 5.15e+10Hz 0.911105 -0.38805
+ 5.16e+10Hz 0.910797 -0.388754
+ 5.17e+10Hz 0.910488 -0.389457
+ 5.18e+10Hz 0.910179 -0.390159
+ 5.19e+10Hz 0.90987 -0.390862
+ 5.2e+10Hz 0.90956 -0.391564
+ 5.21e+10Hz 0.90925 -0.392266
+ 5.22e+10Hz 0.908939 -0.392967
+ 5.23e+10Hz 0.908628 -0.393668
+ 5.24e+10Hz 0.908316 -0.394369
+ 5.25e+10Hz 0.908004 -0.39507
+ 5.26e+10Hz 0.907691 -0.395771
+ 5.27e+10Hz 0.907378 -0.396471
+ 5.28e+10Hz 0.907065 -0.397171
+ 5.29e+10Hz 0.906751 -0.39787
+ 5.3e+10Hz 0.906436 -0.39857
+ 5.31e+10Hz 0.906121 -0.399269
+ 5.32e+10Hz 0.905806 -0.399968
+ 5.33e+10Hz 0.90549 -0.400666
+ 5.34e+10Hz 0.905174 -0.401365
+ 5.35e+10Hz 0.904857 -0.402063
+ 5.36e+10Hz 0.90454 -0.402761
+ 5.37e+10Hz 0.904223 -0.403458
+ 5.38e+10Hz 0.903905 -0.404156
+ 5.39e+10Hz 0.903586 -0.404853
+ 5.4e+10Hz 0.903267 -0.40555
+ 5.41e+10Hz 0.902948 -0.406246
+ 5.42e+10Hz 0.902628 -0.406943
+ 5.43e+10Hz 0.902308 -0.407639
+ 5.44e+10Hz 0.901987 -0.408335
+ 5.45e+10Hz 0.901666 -0.409031
+ 5.46e+10Hz 0.901344 -0.409726
+ 5.47e+10Hz 0.901022 -0.410421
+ 5.48e+10Hz 0.9007 -0.411116
+ 5.49e+10Hz 0.900377 -0.411811
+ 5.5e+10Hz 0.900053 -0.412506
+ 5.51e+10Hz 0.899729 -0.4132
+ 5.52e+10Hz 0.899405 -0.413894
+ 5.53e+10Hz 0.89908 -0.414588
+ 5.54e+10Hz 0.898755 -0.415282
+ 5.55e+10Hz 0.898429 -0.415976
+ 5.56e+10Hz 0.898103 -0.416669
+ 5.57e+10Hz 0.897776 -0.417362
+ 5.58e+10Hz 0.897449 -0.418055
+ 5.59e+10Hz 0.897121 -0.418748
+ 5.6e+10Hz 0.896793 -0.41944
+ 5.61e+10Hz 0.896465 -0.420133
+ 5.62e+10Hz 0.896135 -0.420825
+ 5.63e+10Hz 0.895806 -0.421517
+ 5.64e+10Hz 0.895476 -0.422209
+ 5.65e+10Hz 0.895145 -0.4229
+ 5.66e+10Hz 0.894814 -0.423592
+ 5.67e+10Hz 0.894483 -0.424283
+ 5.68e+10Hz 0.894151 -0.424974
+ 5.69e+10Hz 0.893819 -0.425665
+ 5.7e+10Hz 0.893486 -0.426355
+ 5.71e+10Hz 0.893152 -0.427046
+ 5.72e+10Hz 0.892818 -0.427736
+ 5.73e+10Hz 0.892484 -0.428426
+ 5.74e+10Hz 0.892149 -0.429116
+ 5.75e+10Hz 0.891814 -0.429805
+ 5.76e+10Hz 0.891478 -0.430495
+ 5.77e+10Hz 0.891141 -0.431184
+ 5.78e+10Hz 0.890805 -0.431873
+ 5.79e+10Hz 0.890467 -0.432562
+ 5.8e+10Hz 0.890129 -0.433251
+ 5.81e+10Hz 0.889791 -0.433939
+ 5.82e+10Hz 0.889452 -0.434628
+ 5.83e+10Hz 0.889112 -0.435316
+ 5.84e+10Hz 0.888772 -0.436004
+ 5.85e+10Hz 0.888432 -0.436692
+ 5.86e+10Hz 0.888091 -0.43738
+ 5.87e+10Hz 0.887749 -0.438067
+ 5.88e+10Hz 0.887407 -0.438754
+ 5.89e+10Hz 0.887064 -0.439441
+ 5.9e+10Hz 0.886721 -0.440128
+ 5.91e+10Hz 0.886378 -0.440815
+ 5.92e+10Hz 0.886033 -0.441501
+ 5.93e+10Hz 0.885689 -0.442188
+ 5.94e+10Hz 0.885343 -0.442874
+ 5.95e+10Hz 0.884997 -0.44356
+ 5.96e+10Hz 0.884651 -0.444246
+ 5.97e+10Hz 0.884304 -0.444931
+ 5.98e+10Hz 0.883956 -0.445617
+ 5.99e+10Hz 0.883608 -0.446302
+ 6e+10Hz 0.88326 -0.446987
+ 6.01e+10Hz 0.882911 -0.447671
+ 6.02e+10Hz 0.882561 -0.448356
+ 6.03e+10Hz 0.88221 -0.44904
+ 6.04e+10Hz 0.88186 -0.449725
+ 6.05e+10Hz 0.881508 -0.450409
+ 6.06e+10Hz 0.881156 -0.451092
+ 6.07e+10Hz 0.880804 -0.451776
+ 6.08e+10Hz 0.88045 -0.452459
+ 6.09e+10Hz 0.880097 -0.453142
+ 6.1e+10Hz 0.879742 -0.453825
+ 6.11e+10Hz 0.879388 -0.454508
+ 6.12e+10Hz 0.879032 -0.45519
+ 6.13e+10Hz 0.878676 -0.455873
+ 6.14e+10Hz 0.87832 -0.456555
+ 6.15e+10Hz 0.877962 -0.457237
+ 6.16e+10Hz 0.877605 -0.457918
+ 6.17e+10Hz 0.877246 -0.458599
+ 6.18e+10Hz 0.876887 -0.459281
+ 6.19e+10Hz 0.876528 -0.459962
+ 6.2e+10Hz 0.876168 -0.460642
+ 6.21e+10Hz 0.875807 -0.461323
+ 6.22e+10Hz 0.875446 -0.462003
+ 6.23e+10Hz 0.875084 -0.462683
+ 6.24e+10Hz 0.874721 -0.463362
+ 6.25e+10Hz 0.874358 -0.464042
+ 6.26e+10Hz 0.873995 -0.464721
+ 6.27e+10Hz 0.87363 -0.4654
+ 6.28e+10Hz 0.873265 -0.466079
+ 6.29e+10Hz 0.8729 -0.466757
+ 6.3e+10Hz 0.872534 -0.467435
+ 6.31e+10Hz 0.872167 -0.468113
+ 6.32e+10Hz 0.8718 -0.468791
+ 6.33e+10Hz 0.871432 -0.469468
+ 6.34e+10Hz 0.871064 -0.470146
+ 6.35e+10Hz 0.870695 -0.470822
+ 6.36e+10Hz 0.870325 -0.471499
+ 6.37e+10Hz 0.869955 -0.472175
+ 6.38e+10Hz 0.869584 -0.472851
+ 6.39e+10Hz 0.869213 -0.473527
+ 6.4e+10Hz 0.868841 -0.474202
+ 6.41e+10Hz 0.868468 -0.474878
+ 6.42e+10Hz 0.868095 -0.475552
+ 6.43e+10Hz 0.867721 -0.476227
+ 6.44e+10Hz 0.867347 -0.476901
+ 6.45e+10Hz 0.866972 -0.477575
+ 6.46e+10Hz 0.866596 -0.478249
+ 6.47e+10Hz 0.86622 -0.478922
+ 6.48e+10Hz 0.865843 -0.479595
+ 6.49e+10Hz 0.865466 -0.480268
+ 6.5e+10Hz 0.865088 -0.480941
+ 6.51e+10Hz 0.864709 -0.481613
+ 6.52e+10Hz 0.86433 -0.482284
+ 6.53e+10Hz 0.863951 -0.482956
+ 6.54e+10Hz 0.86357 -0.483627
+ 6.55e+10Hz 0.863189 -0.484298
+ 6.56e+10Hz 0.862808 -0.484969
+ 6.57e+10Hz 0.862426 -0.485639
+ 6.58e+10Hz 0.862043 -0.486309
+ 6.59e+10Hz 0.86166 -0.486978
+ 6.6e+10Hz 0.861276 -0.487647
+ 6.61e+10Hz 0.860892 -0.488316
+ 6.62e+10Hz 0.860507 -0.488985
+ 6.63e+10Hz 0.860121 -0.489653
+ 6.64e+10Hz 0.859735 -0.490321
+ 6.65e+10Hz 0.859349 -0.490988
+ 6.66e+10Hz 0.858961 -0.491655
+ 6.67e+10Hz 0.858573 -0.492322
+ 6.68e+10Hz 0.858185 -0.492988
+ 6.69e+10Hz 0.857796 -0.493655
+ 6.7e+10Hz 0.857407 -0.49432
+ 6.71e+10Hz 0.857017 -0.494986
+ 6.72e+10Hz 0.856626 -0.495651
+ 6.73e+10Hz 0.856235 -0.496315
+ 6.74e+10Hz 0.855843 -0.49698
+ 6.75e+10Hz 0.855451 -0.497643
+ 6.76e+10Hz 0.855058 -0.498307
+ 6.77e+10Hz 0.854665 -0.49897
+ 6.78e+10Hz 0.854271 -0.499633
+ 6.79e+10Hz 0.853876 -0.500295
+ 6.8e+10Hz 0.853481 -0.500958
+ 6.81e+10Hz 0.853085 -0.501619
+ 6.82e+10Hz 0.852689 -0.502281
+ 6.83e+10Hz 0.852293 -0.502942
+ 6.84e+10Hz 0.851896 -0.503602
+ 6.85e+10Hz 0.851498 -0.504262
+ 6.86e+10Hz 0.8511 -0.504922
+ 6.87e+10Hz 0.850701 -0.505582
+ 6.88e+10Hz 0.850302 -0.506241
+ 6.89e+10Hz 0.849902 -0.506899
+ 6.9e+10Hz 0.849501 -0.507558
+ 6.91e+10Hz 0.849101 -0.508216
+ 6.92e+10Hz 0.848699 -0.508873
+ 6.93e+10Hz 0.848297 -0.509531
+ 6.94e+10Hz 0.847895 -0.510187
+ 6.95e+10Hz 0.847492 -0.510844
+ 6.96e+10Hz 0.847089 -0.5115
+ 6.97e+10Hz 0.846685 -0.512156
+ 6.98e+10Hz 0.84628 -0.512811
+ 6.99e+10Hz 0.845875 -0.513466
+ 7e+10Hz 0.84547 -0.51412
+ 7.01e+10Hz 0.845064 -0.514774
+ 7.02e+10Hz 0.844658 -0.515428
+ 7.03e+10Hz 0.844251 -0.516082
+ 7.04e+10Hz 0.843843 -0.516735
+ 7.05e+10Hz 0.843436 -0.517387
+ 7.06e+10Hz 0.843027 -0.518039
+ 7.07e+10Hz 0.842618 -0.518691
+ 7.08e+10Hz 0.842209 -0.519343
+ 7.09e+10Hz 0.841799 -0.519994
+ 7.1e+10Hz 0.841389 -0.520645
+ 7.11e+10Hz 0.840978 -0.521295
+ 7.12e+10Hz 0.840567 -0.521945
+ 7.13e+10Hz 0.840155 -0.522595
+ 7.14e+10Hz 0.839743 -0.523244
+ 7.15e+10Hz 0.839331 -0.523893
+ 7.16e+10Hz 0.838918 -0.524541
+ 7.17e+10Hz 0.838504 -0.525189
+ 7.18e+10Hz 0.83809 -0.525837
+ 7.19e+10Hz 0.837676 -0.526484
+ 7.2e+10Hz 0.837261 -0.527131
+ 7.21e+10Hz 0.836845 -0.527778
+ 7.22e+10Hz 0.836429 -0.528424
+ 7.23e+10Hz 0.836013 -0.52907
+ 7.24e+10Hz 0.835596 -0.529716
+ 7.25e+10Hz 0.835179 -0.530361
+ 7.26e+10Hz 0.834762 -0.531005
+ 7.27e+10Hz 0.834343 -0.53165
+ 7.28e+10Hz 0.833925 -0.532294
+ 7.29e+10Hz 0.833506 -0.532938
+ 7.3e+10Hz 0.833087 -0.533581
+ 7.31e+10Hz 0.832667 -0.534224
+ 7.32e+10Hz 0.832246 -0.534867
+ 7.33e+10Hz 0.831826 -0.535509
+ 7.34e+10Hz 0.831404 -0.536151
+ 7.35e+10Hz 0.830983 -0.536792
+ 7.36e+10Hz 0.830561 -0.537434
+ 7.37e+10Hz 0.830138 -0.538075
+ 7.38e+10Hz 0.829715 -0.538715
+ 7.39e+10Hz 0.829292 -0.539355
+ 7.4e+10Hz 0.828868 -0.539995
+ 7.41e+10Hz 0.828444 -0.540635
+ 7.42e+10Hz 0.828019 -0.541274
+ 7.43e+10Hz 0.827594 -0.541913
+ 7.44e+10Hz 0.827168 -0.542551
+ 7.45e+10Hz 0.826742 -0.543189
+ 7.46e+10Hz 0.826316 -0.543827
+ 7.47e+10Hz 0.825889 -0.544465
+ 7.48e+10Hz 0.825462 -0.545102
+ 7.49e+10Hz 0.825034 -0.545739
+ 7.5e+10Hz 0.824606 -0.546375
+ 7.51e+10Hz 0.824177 -0.547011
+ 7.52e+10Hz 0.823748 -0.547647
+ 7.53e+10Hz 0.823318 -0.548283
+ 7.54e+10Hz 0.822888 -0.548918
+ 7.55e+10Hz 0.822458 -0.549553
+ 7.56e+10Hz 0.822027 -0.550187
+ 7.57e+10Hz 0.821596 -0.550821
+ 7.58e+10Hz 0.821164 -0.551455
+ 7.59e+10Hz 0.820732 -0.552089
+ 7.6e+10Hz 0.8203 -0.552722
+ 7.61e+10Hz 0.819867 -0.553355
+ 7.62e+10Hz 0.819433 -0.553988
+ 7.63e+10Hz 0.819 -0.55462
+ 7.64e+10Hz 0.818565 -0.555252
+ 7.65e+10Hz 0.818131 -0.555884
+ 7.66e+10Hz 0.817695 -0.556515
+ 7.67e+10Hz 0.81726 -0.557146
+ 7.68e+10Hz 0.816824 -0.557777
+ 7.69e+10Hz 0.816387 -0.558408
+ 7.7e+10Hz 0.81595 -0.559038
+ 7.71e+10Hz 0.815513 -0.559668
+ 7.72e+10Hz 0.815075 -0.560297
+ 7.73e+10Hz 0.814637 -0.560926
+ 7.74e+10Hz 0.814198 -0.561555
+ 7.75e+10Hz 0.813759 -0.562184
+ 7.76e+10Hz 0.813319 -0.562812
+ 7.77e+10Hz 0.812879 -0.563441
+ 7.78e+10Hz 0.812439 -0.564068
+ 7.79e+10Hz 0.811998 -0.564696
+ 7.8e+10Hz 0.811556 -0.565323
+ 7.81e+10Hz 0.811114 -0.56595
+ 7.82e+10Hz 0.810672 -0.566576
+ 7.83e+10Hz 0.810229 -0.567203
+ 7.84e+10Hz 0.809786 -0.567829
+ 7.85e+10Hz 0.809342 -0.568454
+ 7.86e+10Hz 0.808898 -0.56908
+ 7.87e+10Hz 0.808453 -0.569705
+ 7.88e+10Hz 0.808008 -0.57033
+ 7.89e+10Hz 0.807563 -0.570954
+ 7.9e+10Hz 0.807117 -0.571579
+ 7.91e+10Hz 0.80667 -0.572202
+ 7.92e+10Hz 0.806223 -0.572826
+ 7.93e+10Hz 0.805776 -0.573449
+ 7.94e+10Hz 0.805328 -0.574072
+ 7.95e+10Hz 0.804879 -0.574695
+ 7.96e+10Hz 0.804431 -0.575318
+ 7.97e+10Hz 0.803981 -0.57594
+ 7.98e+10Hz 0.803531 -0.576562
+ 7.99e+10Hz 0.803081 -0.577183
+ 8e+10Hz 0.80263 -0.577805
+ 8.01e+10Hz 0.802179 -0.578426
+ 8.02e+10Hz 0.801727 -0.579046
+ 8.03e+10Hz 0.801275 -0.579667
+ 8.04e+10Hz 0.800822 -0.580287
+ 8.05e+10Hz 0.800369 -0.580907
+ 8.06e+10Hz 0.799915 -0.581526
+ 8.07e+10Hz 0.799461 -0.582145
+ 8.08e+10Hz 0.799006 -0.582764
+ 8.09e+10Hz 0.798551 -0.583383
+ 8.1e+10Hz 0.798095 -0.584001
+ 8.11e+10Hz 0.797639 -0.584619
+ 8.12e+10Hz 0.797182 -0.585237
+ 8.13e+10Hz 0.796725 -0.585854
+ 8.14e+10Hz 0.796267 -0.586471
+ 8.15e+10Hz 0.795809 -0.587088
+ 8.16e+10Hz 0.795351 -0.587704
+ 8.17e+10Hz 0.794891 -0.58832
+ 8.18e+10Hz 0.794432 -0.588936
+ 8.19e+10Hz 0.793971 -0.589552
+ 8.2e+10Hz 0.793511 -0.590167
+ 8.21e+10Hz 0.793049 -0.590782
+ 8.22e+10Hz 0.792588 -0.591396
+ 8.23e+10Hz 0.792125 -0.592011
+ 8.24e+10Hz 0.791663 -0.592625
+ 8.25e+10Hz 0.791199 -0.593238
+ 8.26e+10Hz 0.790736 -0.593852
+ 8.27e+10Hz 0.790271 -0.594464
+ 8.28e+10Hz 0.789806 -0.595077
+ 8.29e+10Hz 0.789341 -0.595689
+ 8.3e+10Hz 0.788875 -0.596301
+ 8.31e+10Hz 0.788409 -0.596913
+ 8.32e+10Hz 0.787942 -0.597524
+ 8.33e+10Hz 0.787475 -0.598135
+ 8.34e+10Hz 0.787007 -0.598746
+ 8.35e+10Hz 0.786538 -0.599356
+ 8.36e+10Hz 0.786069 -0.599966
+ 8.37e+10Hz 0.7856 -0.600576
+ 8.38e+10Hz 0.78513 -0.601185
+ 8.39e+10Hz 0.784659 -0.601794
+ 8.4e+10Hz 0.784188 -0.602403
+ 8.41e+10Hz 0.783716 -0.603011
+ 8.42e+10Hz 0.783244 -0.603619
+ 8.43e+10Hz 0.782772 -0.604226
+ 8.44e+10Hz 0.782299 -0.604833
+ 8.45e+10Hz 0.781825 -0.60544
+ 8.46e+10Hz 0.781351 -0.606047
+ 8.47e+10Hz 0.780876 -0.606653
+ 8.48e+10Hz 0.780401 -0.607259
+ 8.49e+10Hz 0.779925 -0.607864
+ 8.5e+10Hz 0.779449 -0.608469
+ 8.51e+10Hz 0.778972 -0.609074
+ 8.52e+10Hz 0.778495 -0.609678
+ 8.53e+10Hz 0.778017 -0.610282
+ 8.54e+10Hz 0.777539 -0.610885
+ 8.55e+10Hz 0.77706 -0.611488
+ 8.56e+10Hz 0.77658 -0.612091
+ 8.57e+10Hz 0.7761 -0.612693
+ 8.58e+10Hz 0.77562 -0.613295
+ 8.59e+10Hz 0.775139 -0.613897
+ 8.6e+10Hz 0.774657 -0.614498
+ 8.61e+10Hz 0.774176 -0.615099
+ 8.62e+10Hz 0.773693 -0.6157
+ 8.63e+10Hz 0.77321 -0.6163
+ 8.64e+10Hz 0.772726 -0.616899
+ 8.65e+10Hz 0.772242 -0.617499
+ 8.66e+10Hz 0.771758 -0.618098
+ 8.67e+10Hz 0.771273 -0.618696
+ 8.68e+10Hz 0.770787 -0.619294
+ 8.69e+10Hz 0.770301 -0.619892
+ 8.7e+10Hz 0.769815 -0.620489
+ 8.71e+10Hz 0.769327 -0.621086
+ 8.72e+10Hz 0.76884 -0.621682
+ 8.73e+10Hz 0.768352 -0.622278
+ 8.74e+10Hz 0.767863 -0.622874
+ 8.75e+10Hz 0.767374 -0.623469
+ 8.76e+10Hz 0.766884 -0.624064
+ 8.77e+10Hz 0.766394 -0.624659
+ 8.78e+10Hz 0.765904 -0.625253
+ 8.79e+10Hz 0.765413 -0.625846
+ 8.8e+10Hz 0.764921 -0.626439
+ 8.81e+10Hz 0.764429 -0.627032
+ 8.82e+10Hz 0.763936 -0.627624
+ 8.83e+10Hz 0.763443 -0.628216
+ 8.84e+10Hz 0.76295 -0.628808
+ 8.85e+10Hz 0.762456 -0.629399
+ 8.86e+10Hz 0.761961 -0.629989
+ 8.87e+10Hz 0.761466 -0.63058
+ 8.88e+10Hz 0.760971 -0.631169
+ 8.89e+10Hz 0.760475 -0.631759
+ 8.9e+10Hz 0.759978 -0.632348
+ 8.91e+10Hz 0.759481 -0.632936
+ 8.92e+10Hz 0.758984 -0.633524
+ 8.93e+10Hz 0.758486 -0.634112
+ 8.94e+10Hz 0.757987 -0.634699
+ 8.95e+10Hz 0.757489 -0.635286
+ 8.96e+10Hz 0.756989 -0.635872
+ 8.97e+10Hz 0.756489 -0.636458
+ 8.98e+10Hz 0.755989 -0.637043
+ 8.99e+10Hz 0.755489 -0.637628
+ 9e+10Hz 0.754987 -0.638213
+ 9.01e+10Hz 0.754486 -0.638797
+ 9.02e+10Hz 0.753984 -0.639381
+ 9.03e+10Hz 0.753481 -0.639964
+ 9.04e+10Hz 0.752978 -0.640547
+ 9.05e+10Hz 0.752475 -0.641129
+ 9.06e+10Hz 0.751971 -0.641711
+ 9.07e+10Hz 0.751466 -0.642292
+ 9.08e+10Hz 0.750961 -0.642873
+ 9.09e+10Hz 0.750456 -0.643454
+ 9.1e+10Hz 0.749951 -0.644034
+ 9.11e+10Hz 0.749444 -0.644614
+ 9.12e+10Hz 0.748938 -0.645193
+ 9.13e+10Hz 0.748431 -0.645772
+ 9.14e+10Hz 0.747923 -0.646351
+ 9.15e+10Hz 0.747415 -0.646928
+ 9.16e+10Hz 0.746907 -0.647506
+ 9.17e+10Hz 0.746398 -0.648083
+ 9.18e+10Hz 0.745889 -0.64866
+ 9.19e+10Hz 0.745379 -0.649236
+ 9.2e+10Hz 0.744869 -0.649812
+ 9.21e+10Hz 0.744359 -0.650387
+ 9.22e+10Hz 0.743848 -0.650962
+ 9.23e+10Hz 0.743337 -0.651536
+ 9.24e+10Hz 0.742825 -0.65211
+ 9.25e+10Hz 0.742313 -0.652684
+ 9.26e+10Hz 0.7418 -0.653257
+ 9.27e+10Hz 0.741287 -0.65383
+ 9.28e+10Hz 0.740774 -0.654402
+ 9.29e+10Hz 0.74026 -0.654974
+ 9.3e+10Hz 0.739745 -0.655545
+ 9.31e+10Hz 0.739231 -0.656116
+ 9.32e+10Hz 0.738716 -0.656687
+ 9.33e+10Hz 0.7382 -0.657257
+ 9.34e+10Hz 0.737684 -0.657827
+ 9.35e+10Hz 0.737168 -0.658396
+ 9.36e+10Hz 0.736651 -0.658965
+ 9.37e+10Hz 0.736134 -0.659533
+ 9.38e+10Hz 0.735617 -0.660101
+ 9.39e+10Hz 0.735099 -0.660668
+ 9.4e+10Hz 0.73458 -0.661235
+ 9.41e+10Hz 0.734062 -0.661802
+ 9.42e+10Hz 0.733542 -0.662368
+ 9.43e+10Hz 0.733023 -0.662934
+ 9.44e+10Hz 0.732503 -0.6635
+ 9.45e+10Hz 0.731983 -0.664065
+ 9.46e+10Hz 0.731462 -0.664629
+ 9.47e+10Hz 0.730941 -0.665193
+ 9.48e+10Hz 0.730419 -0.665757
+ 9.49e+10Hz 0.729897 -0.66632
+ 9.5e+10Hz 0.729375 -0.666883
+ 9.51e+10Hz 0.728852 -0.667446
+ 9.52e+10Hz 0.728329 -0.668008
+ 9.53e+10Hz 0.727806 -0.668569
+ 9.54e+10Hz 0.727282 -0.669131
+ 9.55e+10Hz 0.726758 -0.669691
+ 9.56e+10Hz 0.726233 -0.670252
+ 9.57e+10Hz 0.725708 -0.670812
+ 9.58e+10Hz 0.725182 -0.671371
+ 9.59e+10Hz 0.724657 -0.671931
+ 9.6e+10Hz 0.72413 -0.672489
+ 9.61e+10Hz 0.723604 -0.673048
+ 9.62e+10Hz 0.723077 -0.673606
+ 9.63e+10Hz 0.722549 -0.674163
+ 9.64e+10Hz 0.722022 -0.67472
+ 9.65e+10Hz 0.721493 -0.675277
+ 9.66e+10Hz 0.720965 -0.675833
+ 9.67e+10Hz 0.720436 -0.676389
+ 9.68e+10Hz 0.719906 -0.676945
+ 9.69e+10Hz 0.719377 -0.6775
+ 9.7e+10Hz 0.718847 -0.678055
+ 9.71e+10Hz 0.718316 -0.678609
+ 9.72e+10Hz 0.717785 -0.679163
+ 9.73e+10Hz 0.717254 -0.679717
+ 9.74e+10Hz 0.716722 -0.68027
+ 9.75e+10Hz 0.71619 -0.680823
+ 9.76e+10Hz 0.715658 -0.681375
+ 9.77e+10Hz 0.715125 -0.681927
+ 9.78e+10Hz 0.714591 -0.682479
+ 9.79e+10Hz 0.714058 -0.68303
+ 9.8e+10Hz 0.713524 -0.683581
+ 9.81e+10Hz 0.712989 -0.684132
+ 9.82e+10Hz 0.712454 -0.684682
+ 9.83e+10Hz 0.711919 -0.685231
+ 9.84e+10Hz 0.711383 -0.685781
+ 9.85e+10Hz 0.710847 -0.68633
+ 9.86e+10Hz 0.710311 -0.686878
+ 9.87e+10Hz 0.709774 -0.687426
+ 9.88e+10Hz 0.709237 -0.687974
+ 9.89e+10Hz 0.708699 -0.688521
+ 9.9e+10Hz 0.708161 -0.689068
+ 9.91e+10Hz 0.707623 -0.689615
+ 9.92e+10Hz 0.707084 -0.690161
+ 9.93e+10Hz 0.706545 -0.690707
+ 9.94e+10Hz 0.706005 -0.691253
+ 9.95e+10Hz 0.705465 -0.691798
+ 9.96e+10Hz 0.704924 -0.692343
+ 9.97e+10Hz 0.704383 -0.692887
+ 9.98e+10Hz 0.703842 -0.693431
+ 9.99e+10Hz 0.7033 -0.693975
+ 1e+11Hz 0.702758 -0.694518
+ 1.001e+11Hz 0.702216 -0.695061
+ 1.002e+11Hz 0.701673 -0.695603
+ 1.003e+11Hz 0.70113 -0.696145
+ 1.004e+11Hz 0.700586 -0.696687
+ 1.005e+11Hz 0.700042 -0.697228
+ 1.006e+11Hz 0.699497 -0.697769
+ 1.007e+11Hz 0.698952 -0.69831
+ 1.008e+11Hz 0.698407 -0.69885
+ 1.009e+11Hz 0.697861 -0.69939
+ 1.01e+11Hz 0.697314 -0.699929
+ 1.011e+11Hz 0.696768 -0.700468
+ 1.012e+11Hz 0.696221 -0.701007
+ 1.013e+11Hz 0.695673 -0.701545
+ 1.014e+11Hz 0.695125 -0.702083
+ 1.015e+11Hz 0.694577 -0.702621
+ 1.016e+11Hz 0.694028 -0.703158
+ 1.017e+11Hz 0.693479 -0.703694
+ 1.018e+11Hz 0.692929 -0.704231
+ 1.019e+11Hz 0.692379 -0.704767
+ 1.02e+11Hz 0.691828 -0.705302
+ 1.021e+11Hz 0.691277 -0.705838
+ 1.022e+11Hz 0.690726 -0.706373
+ 1.023e+11Hz 0.690174 -0.706907
+ 1.024e+11Hz 0.689622 -0.707441
+ 1.025e+11Hz 0.689069 -0.707975
+ 1.026e+11Hz 0.688516 -0.708508
+ 1.027e+11Hz 0.687962 -0.709041
+ 1.028e+11Hz 0.687408 -0.709573
+ 1.029e+11Hz 0.686854 -0.710106
+ 1.03e+11Hz 0.686299 -0.710637
+ 1.031e+11Hz 0.685743 -0.711169
+ 1.032e+11Hz 0.685188 -0.711699
+ 1.033e+11Hz 0.684631 -0.71223
+ 1.034e+11Hz 0.684075 -0.71276
+ 1.035e+11Hz 0.683518 -0.71329
+ 1.036e+11Hz 0.68296 -0.713819
+ 1.037e+11Hz 0.682402 -0.714348
+ 1.038e+11Hz 0.681844 -0.714877
+ 1.039e+11Hz 0.681285 -0.715405
+ 1.04e+11Hz 0.680725 -0.715932
+ 1.041e+11Hz 0.680165 -0.71646
+ 1.042e+11Hz 0.679605 -0.716987
+ 1.043e+11Hz 0.679044 -0.717513
+ 1.044e+11Hz 0.678483 -0.718039
+ 1.045e+11Hz 0.677922 -0.718565
+ 1.046e+11Hz 0.67736 -0.71909
+ 1.047e+11Hz 0.676797 -0.719615
+ 1.048e+11Hz 0.676234 -0.720139
+ 1.049e+11Hz 0.675671 -0.720663
+ 1.05e+11Hz 0.675107 -0.721187
+ 1.051e+11Hz 0.674543 -0.72171
+ 1.052e+11Hz 0.673978 -0.722233
+ 1.053e+11Hz 0.673413 -0.722755
+ 1.054e+11Hz 0.672847 -0.723277
+ 1.055e+11Hz 0.672281 -0.723799
+ 1.056e+11Hz 0.671714 -0.72432
+ 1.057e+11Hz 0.671147 -0.72484
+ 1.058e+11Hz 0.67058 -0.72536
+ 1.059e+11Hz 0.670012 -0.72588
+ 1.06e+11Hz 0.669444 -0.7264
+ 1.061e+11Hz 0.668875 -0.726918
+ 1.062e+11Hz 0.668305 -0.727437
+ 1.063e+11Hz 0.667736 -0.727955
+ 1.064e+11Hz 0.667166 -0.728472
+ 1.065e+11Hz 0.666595 -0.728989
+ 1.066e+11Hz 0.666024 -0.729506
+ 1.067e+11Hz 0.665452 -0.730022
+ 1.068e+11Hz 0.66488 -0.730538
+ 1.069e+11Hz 0.664308 -0.731053
+ 1.07e+11Hz 0.663735 -0.731568
+ 1.071e+11Hz 0.663162 -0.732083
+ 1.072e+11Hz 0.662588 -0.732597
+ 1.073e+11Hz 0.662014 -0.73311
+ 1.074e+11Hz 0.661439 -0.733623
+ 1.075e+11Hz 0.660864 -0.734136
+ 1.076e+11Hz 0.660288 -0.734648
+ 1.077e+11Hz 0.659712 -0.73516
+ 1.078e+11Hz 0.659136 -0.735671
+ 1.079e+11Hz 0.658559 -0.736182
+ 1.08e+11Hz 0.657982 -0.736692
+ 1.081e+11Hz 0.657404 -0.737202
+ 1.082e+11Hz 0.656826 -0.737711
+ 1.083e+11Hz 0.656247 -0.73822
+ 1.084e+11Hz 0.655668 -0.738728
+ 1.085e+11Hz 0.655088 -0.739236
+ 1.086e+11Hz 0.654508 -0.739744
+ 1.087e+11Hz 0.653928 -0.740251
+ 1.088e+11Hz 0.653347 -0.740757
+ 1.089e+11Hz 0.652766 -0.741263
+ 1.09e+11Hz 0.652184 -0.741769
+ 1.091e+11Hz 0.651602 -0.742274
+ 1.092e+11Hz 0.65102 -0.742778
+ 1.093e+11Hz 0.650437 -0.743282
+ 1.094e+11Hz 0.649853 -0.743786
+ 1.095e+11Hz 0.649269 -0.744289
+ 1.096e+11Hz 0.648685 -0.744792
+ 1.097e+11Hz 0.6481 -0.745294
+ 1.098e+11Hz 0.647515 -0.745796
+ 1.099e+11Hz 0.64693 -0.746297
+ 1.1e+11Hz 0.646344 -0.746797
+ 1.101e+11Hz 0.645757 -0.747298
+ 1.102e+11Hz 0.645171 -0.747797
+ 1.103e+11Hz 0.644583 -0.748297
+ 1.104e+11Hz 0.643996 -0.748795
+ 1.105e+11Hz 0.643408 -0.749293
+ 1.106e+11Hz 0.642819 -0.749791
+ 1.107e+11Hz 0.642231 -0.750288
+ 1.108e+11Hz 0.641641 -0.750785
+ 1.109e+11Hz 0.641052 -0.751281
+ 1.11e+11Hz 0.640462 -0.751777
+ 1.111e+11Hz 0.639871 -0.752272
+ 1.112e+11Hz 0.63928 -0.752767
+ 1.113e+11Hz 0.638689 -0.753261
+ 1.114e+11Hz 0.638097 -0.753755
+ 1.115e+11Hz 0.637505 -0.754248
+ 1.116e+11Hz 0.636913 -0.754741
+ 1.117e+11Hz 0.63632 -0.755233
+ 1.118e+11Hz 0.635727 -0.755725
+ 1.119e+11Hz 0.635133 -0.756216
+ 1.12e+11Hz 0.634539 -0.756707
+ 1.121e+11Hz 0.633944 -0.757197
+ 1.122e+11Hz 0.63335 -0.757687
+ 1.123e+11Hz 0.632754 -0.758176
+ 1.124e+11Hz 0.632159 -0.758665
+ 1.125e+11Hz 0.631563 -0.759153
+ 1.126e+11Hz 0.630966 -0.75964
+ 1.127e+11Hz 0.63037 -0.760128
+ 1.128e+11Hz 0.629773 -0.760614
+ 1.129e+11Hz 0.629175 -0.761101
+ 1.13e+11Hz 0.628577 -0.761586
+ 1.131e+11Hz 0.627979 -0.762071
+ 1.132e+11Hz 0.62738 -0.762556
+ 1.133e+11Hz 0.626781 -0.76304
+ 1.134e+11Hz 0.626182 -0.763524
+ 1.135e+11Hz 0.625582 -0.764007
+ 1.136e+11Hz 0.624982 -0.76449
+ 1.137e+11Hz 0.624382 -0.764972
+ 1.138e+11Hz 0.623781 -0.765453
+ 1.139e+11Hz 0.62318 -0.765935
+ 1.14e+11Hz 0.622578 -0.766415
+ 1.141e+11Hz 0.621976 -0.766895
+ 1.142e+11Hz 0.621374 -0.767375
+ 1.143e+11Hz 0.620771 -0.767854
+ 1.144e+11Hz 0.620168 -0.768333
+ 1.145e+11Hz 0.619565 -0.768811
+ 1.146e+11Hz 0.618961 -0.769288
+ 1.147e+11Hz 0.618357 -0.769766
+ 1.148e+11Hz 0.617753 -0.770242
+ 1.149e+11Hz 0.617148 -0.770718
+ 1.15e+11Hz 0.616543 -0.771194
+ 1.151e+11Hz 0.615938 -0.771669
+ 1.152e+11Hz 0.615332 -0.772144
+ 1.153e+11Hz 0.614726 -0.772618
+ 1.154e+11Hz 0.614119 -0.773091
+ 1.155e+11Hz 0.613512 -0.773565
+ 1.156e+11Hz 0.612905 -0.774037
+ 1.157e+11Hz 0.612298 -0.774509
+ 1.158e+11Hz 0.61169 -0.774981
+ 1.159e+11Hz 0.611081 -0.775452
+ 1.16e+11Hz 0.610473 -0.775923
+ 1.161e+11Hz 0.609864 -0.776393
+ 1.162e+11Hz 0.609255 -0.776863
+ 1.163e+11Hz 0.608645 -0.777332
+ 1.164e+11Hz 0.608035 -0.777801
+ 1.165e+11Hz 0.607425 -0.778269
+ 1.166e+11Hz 0.606814 -0.778737
+ 1.167e+11Hz 0.606203 -0.779204
+ 1.168e+11Hz 0.605592 -0.779671
+ 1.169e+11Hz 0.60498 -0.780137
+ 1.17e+11Hz 0.604368 -0.780603
+ 1.171e+11Hz 0.603756 -0.781068
+ 1.172e+11Hz 0.603144 -0.781533
+ 1.173e+11Hz 0.602531 -0.781997
+ 1.174e+11Hz 0.601917 -0.782461
+ 1.175e+11Hz 0.601304 -0.782925
+ 1.176e+11Hz 0.60069 -0.783388
+ 1.177e+11Hz 0.600075 -0.78385
+ 1.178e+11Hz 0.599461 -0.784312
+ 1.179e+11Hz 0.598846 -0.784774
+ 1.18e+11Hz 0.59823 -0.785235
+ 1.181e+11Hz 0.597615 -0.785695
+ 1.182e+11Hz 0.596999 -0.786155
+ 1.183e+11Hz 0.596382 -0.786615
+ 1.184e+11Hz 0.595766 -0.787074
+ 1.185e+11Hz 0.595149 -0.787533
+ 1.186e+11Hz 0.594531 -0.787991
+ 1.187e+11Hz 0.593914 -0.788448
+ 1.188e+11Hz 0.593296 -0.788906
+ 1.189e+11Hz 0.592677 -0.789362
+ 1.19e+11Hz 0.592059 -0.789819
+ 1.191e+11Hz 0.59144 -0.790274
+ 1.192e+11Hz 0.59082 -0.79073
+ 1.193e+11Hz 0.590201 -0.791185
+ 1.194e+11Hz 0.589581 -0.791639
+ 1.195e+11Hz 0.58896 -0.792093
+ 1.196e+11Hz 0.58834 -0.792547
+ 1.197e+11Hz 0.587719 -0.793
+ 1.198e+11Hz 0.587097 -0.793452
+ 1.199e+11Hz 0.586475 -0.793904
+ 1.2e+11Hz 0.585853 -0.794356
+ 1.201e+11Hz 0.585231 -0.794807
+ 1.202e+11Hz 0.584608 -0.795258
+ 1.203e+11Hz 0.583985 -0.795708
+ 1.204e+11Hz 0.583362 -0.796158
+ 1.205e+11Hz 0.582738 -0.796607
+ 1.206e+11Hz 0.582114 -0.797056
+ 1.207e+11Hz 0.58149 -0.797504
+ 1.208e+11Hz 0.580865 -0.797952
+ 1.209e+11Hz 0.58024 -0.798399
+ 1.21e+11Hz 0.579614 -0.798846
+ 1.211e+11Hz 0.578988 -0.799293
+ 1.212e+11Hz 0.578362 -0.799739
+ 1.213e+11Hz 0.577736 -0.800185
+ 1.214e+11Hz 0.577109 -0.80063
+ 1.215e+11Hz 0.576482 -0.801074
+ 1.216e+11Hz 0.575854 -0.801519
+ 1.217e+11Hz 0.575226 -0.801962
+ 1.218e+11Hz 0.574598 -0.802406
+ 1.219e+11Hz 0.573969 -0.802848
+ 1.22e+11Hz 0.57334 -0.803291
+ 1.221e+11Hz 0.572711 -0.803733
+ 1.222e+11Hz 0.572081 -0.804174
+ 1.223e+11Hz 0.571451 -0.804615
+ 1.224e+11Hz 0.570821 -0.805055
+ 1.225e+11Hz 0.57019 -0.805495
+ 1.226e+11Hz 0.569559 -0.805935
+ 1.227e+11Hz 0.568928 -0.806374
+ 1.228e+11Hz 0.568296 -0.806813
+ 1.229e+11Hz 0.567664 -0.807251
+ 1.23e+11Hz 0.567032 -0.807689
+ 1.231e+11Hz 0.566399 -0.808126
+ 1.232e+11Hz 0.565765 -0.808563
+ 1.233e+11Hz 0.565132 -0.808999
+ 1.234e+11Hz 0.564498 -0.809435
+ 1.235e+11Hz 0.563864 -0.80987
+ 1.236e+11Hz 0.563229 -0.810305
+ 1.237e+11Hz 0.562594 -0.810739
+ 1.238e+11Hz 0.561959 -0.811173
+ 1.239e+11Hz 0.561323 -0.811607
+ 1.24e+11Hz 0.560687 -0.81204
+ 1.241e+11Hz 0.56005 -0.812472
+ 1.242e+11Hz 0.559413 -0.812904
+ 1.243e+11Hz 0.558776 -0.813336
+ 1.244e+11Hz 0.558139 -0.813767
+ 1.245e+11Hz 0.557501 -0.814198
+ 1.246e+11Hz 0.556862 -0.814628
+ 1.247e+11Hz 0.556224 -0.815057
+ 1.248e+11Hz 0.555585 -0.815487
+ 1.249e+11Hz 0.554945 -0.815915
+ 1.25e+11Hz 0.554305 -0.816343
+ 1.251e+11Hz 0.553665 -0.816771
+ 1.252e+11Hz 0.553025 -0.817198
+ 1.253e+11Hz 0.552384 -0.817625
+ 1.254e+11Hz 0.551743 -0.818051
+ 1.255e+11Hz 0.551101 -0.818477
+ 1.256e+11Hz 0.550459 -0.818902
+ 1.257e+11Hz 0.549817 -0.819327
+ 1.258e+11Hz 0.549174 -0.819752
+ 1.259e+11Hz 0.548531 -0.820175
+ 1.26e+11Hz 0.547887 -0.820599
+ 1.261e+11Hz 0.547243 -0.821021
+ 1.262e+11Hz 0.546599 -0.821444
+ 1.263e+11Hz 0.545954 -0.821866
+ 1.264e+11Hz 0.54531 -0.822287
+ 1.265e+11Hz 0.544664 -0.822708
+ 1.266e+11Hz 0.544018 -0.823128
+ 1.267e+11Hz 0.543372 -0.823548
+ 1.268e+11Hz 0.542726 -0.823967
+ 1.269e+11Hz 0.542079 -0.824386
+ 1.27e+11Hz 0.541432 -0.824804
+ 1.271e+11Hz 0.540784 -0.825222
+ 1.272e+11Hz 0.540136 -0.825639
+ 1.273e+11Hz 0.539488 -0.826056
+ 1.274e+11Hz 0.538839 -0.826472
+ 1.275e+11Hz 0.53819 -0.826888
+ 1.276e+11Hz 0.537541 -0.827303
+ 1.277e+11Hz 0.536891 -0.827718
+ 1.278e+11Hz 0.536241 -0.828132
+ 1.279e+11Hz 0.53559 -0.828546
+ 1.28e+11Hz 0.534939 -0.828959
+ 1.281e+11Hz 0.534288 -0.829372
+ 1.282e+11Hz 0.533636 -0.829784
+ 1.283e+11Hz 0.532984 -0.830195
+ 1.284e+11Hz 0.532332 -0.830606
+ 1.285e+11Hz 0.531679 -0.831017
+ 1.286e+11Hz 0.531026 -0.831427
+ 1.287e+11Hz 0.530373 -0.831836
+ 1.288e+11Hz 0.529719 -0.832245
+ 1.289e+11Hz 0.529065 -0.832654
+ 1.29e+11Hz 0.52841 -0.833062
+ 1.291e+11Hz 0.527755 -0.833469
+ 1.292e+11Hz 0.5271 -0.833876
+ 1.293e+11Hz 0.526444 -0.834282
+ 1.294e+11Hz 0.525788 -0.834688
+ 1.295e+11Hz 0.525132 -0.835093
+ 1.296e+11Hz 0.524475 -0.835498
+ 1.297e+11Hz 0.523818 -0.835902
+ 1.298e+11Hz 0.52316 -0.836305
+ 1.299e+11Hz 0.522503 -0.836708
+ 1.3e+11Hz 0.521844 -0.837111
+ 1.301e+11Hz 0.521186 -0.837513
+ 1.302e+11Hz 0.520527 -0.837914
+ 1.303e+11Hz 0.519868 -0.838315
+ 1.304e+11Hz 0.519208 -0.838715
+ 1.305e+11Hz 0.518548 -0.839115
+ 1.306e+11Hz 0.517888 -0.839514
+ 1.307e+11Hz 0.517228 -0.839912
+ 1.308e+11Hz 0.516567 -0.84031
+ 1.309e+11Hz 0.515905 -0.840708
+ 1.31e+11Hz 0.515244 -0.841105
+ 1.311e+11Hz 0.514582 -0.841501
+ 1.312e+11Hz 0.513919 -0.841897
+ 1.313e+11Hz 0.513257 -0.842292
+ 1.314e+11Hz 0.512594 -0.842687
+ 1.315e+11Hz 0.51193 -0.843081
+ 1.316e+11Hz 0.511267 -0.843475
+ 1.317e+11Hz 0.510603 -0.843868
+ 1.318e+11Hz 0.509938 -0.84426
+ 1.319e+11Hz 0.509274 -0.844652
+ 1.32e+11Hz 0.508609 -0.845043
+ 1.321e+11Hz 0.507943 -0.845434
+ 1.322e+11Hz 0.507278 -0.845824
+ 1.323e+11Hz 0.506612 -0.846214
+ 1.324e+11Hz 0.505945 -0.846603
+ 1.325e+11Hz 0.505279 -0.846992
+ 1.326e+11Hz 0.504612 -0.847379
+ 1.327e+11Hz 0.503944 -0.847767
+ 1.328e+11Hz 0.503277 -0.848154
+ 1.329e+11Hz 0.502609 -0.84854
+ 1.33e+11Hz 0.501941 -0.848925
+ 1.331e+11Hz 0.501272 -0.84931
+ 1.332e+11Hz 0.500603 -0.849695
+ 1.333e+11Hz 0.499934 -0.850079
+ 1.334e+11Hz 0.499265 -0.850462
+ 1.335e+11Hz 0.498595 -0.850845
+ 1.336e+11Hz 0.497925 -0.851227
+ 1.337e+11Hz 0.497254 -0.851609
+ 1.338e+11Hz 0.496584 -0.85199
+ 1.339e+11Hz 0.495913 -0.85237
+ 1.34e+11Hz 0.495241 -0.85275
+ 1.341e+11Hz 0.49457 -0.85313
+ 1.342e+11Hz 0.493898 -0.853509
+ 1.343e+11Hz 0.493225 -0.853887
+ 1.344e+11Hz 0.492553 -0.854264
+ 1.345e+11Hz 0.49188 -0.854641
+ 1.346e+11Hz 0.491207 -0.855018
+ 1.347e+11Hz 0.490534 -0.855394
+ 1.348e+11Hz 0.48986 -0.855769
+ 1.349e+11Hz 0.489186 -0.856144
+ 1.35e+11Hz 0.488512 -0.856518
+ 1.351e+11Hz 0.487837 -0.856892
+ 1.352e+11Hz 0.487162 -0.857265
+ 1.353e+11Hz 0.486487 -0.857637
+ 1.354e+11Hz 0.485812 -0.858009
+ 1.355e+11Hz 0.485136 -0.858381
+ 1.356e+11Hz 0.48446 -0.858751
+ 1.357e+11Hz 0.483784 -0.859122
+ 1.358e+11Hz 0.483107 -0.859491
+ 1.359e+11Hz 0.48243 -0.85986
+ 1.36e+11Hz 0.481753 -0.860229
+ 1.361e+11Hz 0.481076 -0.860597
+ 1.362e+11Hz 0.480398 -0.860964
+ 1.363e+11Hz 0.47972 -0.861331
+ 1.364e+11Hz 0.479042 -0.861697
+ 1.365e+11Hz 0.478363 -0.862063
+ 1.366e+11Hz 0.477684 -0.862428
+ 1.367e+11Hz 0.477005 -0.862792
+ 1.368e+11Hz 0.476326 -0.863156
+ 1.369e+11Hz 0.475646 -0.86352
+ 1.37e+11Hz 0.474967 -0.863882
+ 1.371e+11Hz 0.474286 -0.864245
+ 1.372e+11Hz 0.473606 -0.864606
+ 1.373e+11Hz 0.472925 -0.864967
+ 1.374e+11Hz 0.472244 -0.865328
+ 1.375e+11Hz 0.471563 -0.865688
+ 1.376e+11Hz 0.470882 -0.866047
+ 1.377e+11Hz 0.4702 -0.866406
+ 1.378e+11Hz 0.469518 -0.866765
+ 1.379e+11Hz 0.468836 -0.867122
+ 1.38e+11Hz 0.468153 -0.867479
+ 1.381e+11Hz 0.46747 -0.867836
+ 1.382e+11Hz 0.466787 -0.868192
+ 1.383e+11Hz 0.466104 -0.868548
+ 1.384e+11Hz 0.46542 -0.868903
+ 1.385e+11Hz 0.464737 -0.869257
+ 1.386e+11Hz 0.464053 -0.869611
+ 1.387e+11Hz 0.463368 -0.869964
+ 1.388e+11Hz 0.462684 -0.870317
+ 1.389e+11Hz 0.461999 -0.870669
+ 1.39e+11Hz 0.461314 -0.871021
+ 1.391e+11Hz 0.460628 -0.871372
+ 1.392e+11Hz 0.459942 -0.871722
+ 1.393e+11Hz 0.459257 -0.872072
+ 1.394e+11Hz 0.45857 -0.872422
+ 1.395e+11Hz 0.457884 -0.87277
+ 1.396e+11Hz 0.457197 -0.873119
+ 1.397e+11Hz 0.45651 -0.873466
+ 1.398e+11Hz 0.455823 -0.873814
+ 1.399e+11Hz 0.455136 -0.87416
+ 1.4e+11Hz 0.454448 -0.874506
+ 1.401e+11Hz 0.45376 -0.874852
+ 1.402e+11Hz 0.453072 -0.875197
+ 1.403e+11Hz 0.452383 -0.875541
+ 1.404e+11Hz 0.451694 -0.875885
+ 1.405e+11Hz 0.451005 -0.876229
+ 1.406e+11Hz 0.450316 -0.876571
+ 1.407e+11Hz 0.449627 -0.876914
+ 1.408e+11Hz 0.448937 -0.877255
+ 1.409e+11Hz 0.448247 -0.877597
+ 1.41e+11Hz 0.447556 -0.877937
+ 1.411e+11Hz 0.446866 -0.878277
+ 1.412e+11Hz 0.446175 -0.878617
+ 1.413e+11Hz 0.445484 -0.878956
+ 1.414e+11Hz 0.444793 -0.879294
+ 1.415e+11Hz 0.444101 -0.879632
+ 1.416e+11Hz 0.443409 -0.879969
+ 1.417e+11Hz 0.442717 -0.880306
+ 1.418e+11Hz 0.442025 -0.880642
+ 1.419e+11Hz 0.441332 -0.880978
+ 1.42e+11Hz 0.440639 -0.881313
+ 1.421e+11Hz 0.439946 -0.881648
+ 1.422e+11Hz 0.439252 -0.881982
+ 1.423e+11Hz 0.438559 -0.882316
+ 1.424e+11Hz 0.437865 -0.882649
+ 1.425e+11Hz 0.437171 -0.882981
+ 1.426e+11Hz 0.436476 -0.883313
+ 1.427e+11Hz 0.435781 -0.883644
+ 1.428e+11Hz 0.435086 -0.883975
+ 1.429e+11Hz 0.434391 -0.884305
+ 1.43e+11Hz 0.433695 -0.884635
+ 1.431e+11Hz 0.433 -0.884964
+ 1.432e+11Hz 0.432304 -0.885293
+ 1.433e+11Hz 0.431607 -0.885621
+ 1.434e+11Hz 0.430911 -0.885948
+ 1.435e+11Hz 0.430214 -0.886275
+ 1.436e+11Hz 0.429517 -0.886602
+ 1.437e+11Hz 0.428819 -0.886927
+ 1.438e+11Hz 0.428121 -0.887253
+ 1.439e+11Hz 0.427423 -0.887578
+ 1.44e+11Hz 0.426725 -0.887902
+ 1.441e+11Hz 0.426027 -0.888225
+ 1.442e+11Hz 0.425328 -0.888548
+ 1.443e+11Hz 0.424629 -0.888871
+ 1.444e+11Hz 0.42393 -0.889193
+ 1.445e+11Hz 0.42323 -0.889514
+ 1.446e+11Hz 0.42253 -0.889835
+ 1.447e+11Hz 0.42183 -0.890156
+ 1.448e+11Hz 0.42113 -0.890476
+ 1.449e+11Hz 0.420429 -0.890795
+ 1.45e+11Hz 0.419728 -0.891113
+ 1.451e+11Hz 0.419027 -0.891432
+ 1.452e+11Hz 0.418325 -0.891749
+ 1.453e+11Hz 0.417623 -0.892066
+ 1.454e+11Hz 0.416921 -0.892382
+ 1.455e+11Hz 0.416219 -0.892698
+ 1.456e+11Hz 0.415517 -0.893014
+ 1.457e+11Hz 0.414814 -0.893328
+ 1.458e+11Hz 0.41411 -0.893643
+ 1.459e+11Hz 0.413407 -0.893956
+ 1.46e+11Hz 0.412703 -0.894269
+ 1.461e+11Hz 0.411999 -0.894582
+ 1.462e+11Hz 0.411295 -0.894894
+ 1.463e+11Hz 0.410591 -0.895205
+ 1.464e+11Hz 0.409886 -0.895516
+ 1.465e+11Hz 0.409181 -0.895826
+ 1.466e+11Hz 0.408475 -0.896136
+ 1.467e+11Hz 0.40777 -0.896445
+ 1.468e+11Hz 0.407064 -0.896753
+ 1.469e+11Hz 0.406358 -0.897061
+ 1.47e+11Hz 0.405651 -0.897368
+ 1.471e+11Hz 0.404944 -0.897675
+ 1.472e+11Hz 0.404237 -0.897981
+ 1.473e+11Hz 0.40353 -0.898287
+ 1.474e+11Hz 0.402823 -0.898592
+ 1.475e+11Hz 0.402115 -0.898896
+ 1.476e+11Hz 0.401407 -0.8992
+ 1.477e+11Hz 0.400698 -0.899503
+ 1.478e+11Hz 0.39999 -0.899806
+ 1.479e+11Hz 0.399281 -0.900108
+ 1.48e+11Hz 0.398572 -0.900409
+ 1.481e+11Hz 0.397862 -0.90071
+ 1.482e+11Hz 0.397152 -0.90101
+ 1.483e+11Hz 0.396442 -0.90131
+ 1.484e+11Hz 0.395732 -0.901609
+ 1.485e+11Hz 0.395021 -0.901908
+ 1.486e+11Hz 0.394311 -0.902205
+ 1.487e+11Hz 0.393599 -0.902503
+ 1.488e+11Hz 0.392888 -0.902799
+ 1.489e+11Hz 0.392176 -0.903095
+ 1.49e+11Hz 0.391465 -0.903391
+ 1.491e+11Hz 0.390752 -0.903686
+ 1.492e+11Hz 0.39004 -0.90398
+ 1.493e+11Hz 0.389327 -0.904274
+ 1.494e+11Hz 0.388614 -0.904567
+ 1.495e+11Hz 0.387901 -0.904859
+ 1.496e+11Hz 0.387187 -0.905151
+ 1.497e+11Hz 0.386474 -0.905442
+ 1.498e+11Hz 0.38576 -0.905733
+ 1.499e+11Hz 0.385045 -0.906023
+ 1.5e+11Hz 0.384331 -0.906312
+ 1.501e+11Hz 0.383616 -0.906601
+ 1.502e+11Hz 0.382901 -0.906889
+ 1.503e+11Hz 0.382186 -0.907176
+ 1.504e+11Hz 0.38147 -0.907463
+ 1.505e+11Hz 0.380754 -0.907749
+ 1.506e+11Hz 0.380038 -0.908035
+ 1.507e+11Hz 0.379322 -0.90832
+ 1.508e+11Hz 0.378605 -0.908604
+ 1.509e+11Hz 0.377888 -0.908888
+ 1.51e+11Hz 0.377171 -0.909171
+ 1.511e+11Hz 0.376454 -0.909453
+ 1.512e+11Hz 0.375736 -0.909735
+ 1.513e+11Hz 0.375018 -0.910016
+ 1.514e+11Hz 0.3743 -0.910297
+ 1.515e+11Hz 0.373582 -0.910577
+ 1.516e+11Hz 0.372863 -0.910856
+ 1.517e+11Hz 0.372145 -0.911135
+ 1.518e+11Hz 0.371426 -0.911413
+ 1.519e+11Hz 0.370706 -0.91169
+ 1.52e+11Hz 0.369987 -0.911967
+ 1.521e+11Hz 0.369267 -0.912243
+ 1.522e+11Hz 0.368547 -0.912518
+ 1.523e+11Hz 0.367827 -0.912793
+ 1.524e+11Hz 0.367107 -0.913067
+ 1.525e+11Hz 0.366386 -0.91334
+ 1.526e+11Hz 0.365665 -0.913613
+ 1.527e+11Hz 0.364944 -0.913885
+ 1.528e+11Hz 0.364223 -0.914157
+ 1.529e+11Hz 0.363501 -0.914428
+ 1.53e+11Hz 0.362779 -0.914698
+ 1.531e+11Hz 0.362057 -0.914967
+ 1.532e+11Hz 0.361335 -0.915236
+ 1.533e+11Hz 0.360613 -0.915504
+ 1.534e+11Hz 0.35989 -0.915772
+ 1.535e+11Hz 0.359167 -0.916039
+ 1.536e+11Hz 0.358444 -0.916305
+ 1.537e+11Hz 0.357721 -0.916571
+ 1.538e+11Hz 0.356997 -0.916836
+ 1.539e+11Hz 0.356274 -0.9171
+ 1.54e+11Hz 0.35555 -0.917364
+ 1.541e+11Hz 0.354826 -0.917627
+ 1.542e+11Hz 0.354102 -0.917889
+ 1.543e+11Hz 0.353377 -0.91815
+ 1.544e+11Hz 0.352652 -0.918411
+ 1.545e+11Hz 0.351928 -0.918672
+ 1.546e+11Hz 0.351203 -0.918931
+ 1.547e+11Hz 0.350477 -0.91919
+ 1.548e+11Hz 0.349752 -0.919449
+ 1.549e+11Hz 0.349026 -0.919706
+ 1.55e+11Hz 0.348301 -0.919963
+ 1.551e+11Hz 0.347575 -0.92022
+ 1.552e+11Hz 0.346849 -0.920475
+ 1.553e+11Hz 0.346122 -0.920731
+ 1.554e+11Hz 0.345396 -0.920985
+ 1.555e+11Hz 0.344669 -0.921239
+ 1.556e+11Hz 0.343942 -0.921492
+ 1.557e+11Hz 0.343215 -0.921744
+ 1.558e+11Hz 0.342488 -0.921996
+ 1.559e+11Hz 0.341761 -0.922247
+ 1.56e+11Hz 0.341033 -0.922497
+ 1.561e+11Hz 0.340306 -0.922747
+ 1.562e+11Hz 0.339578 -0.922996
+ 1.563e+11Hz 0.33885 -0.923244
+ 1.564e+11Hz 0.338122 -0.923492
+ 1.565e+11Hz 0.337393 -0.923739
+ 1.566e+11Hz 0.336665 -0.923985
+ 1.567e+11Hz 0.335936 -0.924231
+ 1.568e+11Hz 0.335207 -0.924476
+ 1.569e+11Hz 0.334479 -0.924721
+ 1.57e+11Hz 0.33375 -0.924964
+ 1.571e+11Hz 0.33302 -0.925207
+ 1.572e+11Hz 0.332291 -0.92545
+ 1.573e+11Hz 0.331561 -0.925692
+ 1.574e+11Hz 0.330832 -0.925933
+ 1.575e+11Hz 0.330102 -0.926173
+ 1.576e+11Hz 0.329372 -0.926413
+ 1.577e+11Hz 0.328642 -0.926652
+ 1.578e+11Hz 0.327912 -0.92689
+ 1.579e+11Hz 0.327182 -0.927128
+ 1.58e+11Hz 0.326451 -0.927365
+ 1.581e+11Hz 0.325721 -0.927602
+ 1.582e+11Hz 0.32499 -0.927838
+ 1.583e+11Hz 0.324259 -0.928073
+ 1.584e+11Hz 0.323528 -0.928307
+ 1.585e+11Hz 0.322797 -0.928541
+ 1.586e+11Hz 0.322066 -0.928774
+ 1.587e+11Hz 0.321335 -0.929007
+ 1.588e+11Hz 0.320603 -0.929239
+ 1.589e+11Hz 0.319872 -0.92947
+ 1.59e+11Hz 0.31914 -0.929701
+ 1.591e+11Hz 0.318408 -0.929931
+ 1.592e+11Hz 0.317676 -0.93016
+ 1.593e+11Hz 0.316944 -0.930389
+ 1.594e+11Hz 0.316212 -0.930617
+ 1.595e+11Hz 0.31548 -0.930844
+ 1.596e+11Hz 0.314747 -0.931071
+ 1.597e+11Hz 0.314015 -0.931297
+ 1.598e+11Hz 0.313282 -0.931522
+ 1.599e+11Hz 0.31255 -0.931747
+ 1.6e+11Hz 0.311817 -0.931971
+ 1.601e+11Hz 0.311084 -0.932194
+ 1.602e+11Hz 0.310351 -0.932417
+ 1.603e+11Hz 0.309618 -0.932639
+ 1.604e+11Hz 0.308885 -0.932861
+ 1.605e+11Hz 0.308152 -0.933082
+ 1.606e+11Hz 0.307418 -0.933302
+ 1.607e+11Hz 0.306685 -0.933522
+ 1.608e+11Hz 0.305951 -0.933741
+ 1.609e+11Hz 0.305217 -0.933959
+ 1.61e+11Hz 0.304484 -0.934177
+ 1.611e+11Hz 0.30375 -0.934394
+ 1.612e+11Hz 0.303016 -0.93461
+ 1.613e+11Hz 0.302282 -0.934826
+ 1.614e+11Hz 0.301548 -0.935041
+ 1.615e+11Hz 0.300813 -0.935256
+ 1.616e+11Hz 0.300079 -0.935469
+ 1.617e+11Hz 0.299345 -0.935683
+ 1.618e+11Hz 0.29861 -0.935895
+ 1.619e+11Hz 0.297876 -0.936107
+ 1.62e+11Hz 0.297141 -0.936319
+ 1.621e+11Hz 0.296406 -0.936529
+ 1.622e+11Hz 0.295671 -0.936739
+ 1.623e+11Hz 0.294937 -0.936949
+ 1.624e+11Hz 0.294202 -0.937158
+ 1.625e+11Hz 0.293466 -0.937366
+ 1.626e+11Hz 0.292731 -0.937574
+ 1.627e+11Hz 0.291996 -0.93778
+ 1.628e+11Hz 0.291261 -0.937987
+ 1.629e+11Hz 0.290525 -0.938193
+ 1.63e+11Hz 0.28979 -0.938398
+ 1.631e+11Hz 0.289054 -0.938602
+ 1.632e+11Hz 0.288319 -0.938806
+ 1.633e+11Hz 0.287583 -0.939009
+ 1.634e+11Hz 0.286847 -0.939212
+ 1.635e+11Hz 0.286111 -0.939414
+ 1.636e+11Hz 0.285375 -0.939615
+ 1.637e+11Hz 0.284639 -0.939816
+ 1.638e+11Hz 0.283903 -0.940016
+ 1.639e+11Hz 0.283167 -0.940215
+ 1.64e+11Hz 0.282431 -0.940414
+ 1.641e+11Hz 0.281694 -0.940612
+ 1.642e+11Hz 0.280958 -0.94081
+ 1.643e+11Hz 0.280221 -0.941007
+ 1.644e+11Hz 0.279485 -0.941203
+ 1.645e+11Hz 0.278748 -0.941399
+ 1.646e+11Hz 0.278012 -0.941594
+ 1.647e+11Hz 0.277275 -0.941789
+ 1.648e+11Hz 0.276538 -0.941983
+ 1.649e+11Hz 0.275801 -0.942176
+ 1.65e+11Hz 0.275064 -0.942369
+ 1.651e+11Hz 0.274327 -0.942561
+ 1.652e+11Hz 0.27359 -0.942752
+ 1.653e+11Hz 0.272853 -0.942943
+ 1.654e+11Hz 0.272116 -0.943133
+ 1.655e+11Hz 0.271378 -0.943323
+ 1.656e+11Hz 0.270641 -0.943512
+ 1.657e+11Hz 0.269903 -0.9437
+ 1.658e+11Hz 0.269166 -0.943888
+ 1.659e+11Hz 0.268428 -0.944075
+ 1.66e+11Hz 0.267691 -0.944262
+ 1.661e+11Hz 0.266953 -0.944448
+ 1.662e+11Hz 0.266215 -0.944633
+ 1.663e+11Hz 0.265478 -0.944818
+ 1.664e+11Hz 0.26474 -0.945002
+ 1.665e+11Hz 0.264002 -0.945185
+ 1.666e+11Hz 0.263264 -0.945368
+ 1.667e+11Hz 0.262526 -0.945551
+ 1.668e+11Hz 0.261788 -0.945732
+ 1.669e+11Hz 0.261049 -0.945913
+ 1.67e+11Hz 0.260311 -0.946094
+ 1.671e+11Hz 0.259573 -0.946273
+ 1.672e+11Hz 0.258834 -0.946453
+ 1.673e+11Hz 0.258096 -0.946631
+ 1.674e+11Hz 0.257358 -0.946809
+ 1.675e+11Hz 0.256619 -0.946987
+ 1.676e+11Hz 0.255881 -0.947163
+ 1.677e+11Hz 0.255142 -0.94734
+ 1.678e+11Hz 0.254403 -0.947515
+ 1.679e+11Hz 0.253665 -0.94769
+ 1.68e+11Hz 0.252926 -0.947864
+ 1.681e+11Hz 0.252187 -0.948038
+ 1.682e+11Hz 0.251448 -0.948211
+ 1.683e+11Hz 0.250709 -0.948384
+ 1.684e+11Hz 0.24997 -0.948556
+ 1.685e+11Hz 0.249231 -0.948727
+ 1.686e+11Hz 0.248492 -0.948898
+ 1.687e+11Hz 0.247753 -0.949068
+ 1.688e+11Hz 0.247014 -0.949237
+ 1.689e+11Hz 0.246275 -0.949406
+ 1.69e+11Hz 0.245535 -0.949574
+ 1.691e+11Hz 0.244796 -0.949742
+ 1.692e+11Hz 0.244057 -0.949909
+ 1.693e+11Hz 0.243317 -0.950075
+ 1.694e+11Hz 0.242578 -0.950241
+ 1.695e+11Hz 0.241839 -0.950406
+ 1.696e+11Hz 0.241099 -0.950571
+ 1.697e+11Hz 0.24036 -0.950735
+ 1.698e+11Hz 0.23962 -0.950898
+ 1.699e+11Hz 0.23888 -0.951061
+ 1.7e+11Hz 0.238141 -0.951223
+ 1.701e+11Hz 0.237401 -0.951384
+ 1.702e+11Hz 0.236662 -0.951545
+ 1.703e+11Hz 0.235922 -0.951706
+ 1.704e+11Hz 0.235182 -0.951865
+ 1.705e+11Hz 0.234442 -0.952024
+ 1.706e+11Hz 0.233703 -0.952183
+ 1.707e+11Hz 0.232963 -0.952341
+ 1.708e+11Hz 0.232223 -0.952498
+ 1.709e+11Hz 0.231483 -0.952655
+ 1.71e+11Hz 0.230743 -0.952811
+ 1.711e+11Hz 0.230003 -0.952966
+ 1.712e+11Hz 0.229263 -0.953121
+ 1.713e+11Hz 0.228523 -0.953275
+ 1.714e+11Hz 0.227783 -0.953429
+ 1.715e+11Hz 0.227043 -0.953582
+ 1.716e+11Hz 0.226303 -0.953735
+ 1.717e+11Hz 0.225563 -0.953886
+ 1.718e+11Hz 0.224823 -0.954038
+ 1.719e+11Hz 0.224083 -0.954188
+ 1.72e+11Hz 0.223343 -0.954338
+ 1.721e+11Hz 0.222603 -0.954488
+ 1.722e+11Hz 0.221863 -0.954637
+ 1.723e+11Hz 0.221123 -0.954785
+ 1.724e+11Hz 0.220383 -0.954933
+ 1.725e+11Hz 0.219643 -0.95508
+ 1.726e+11Hz 0.218903 -0.955226
+ 1.727e+11Hz 0.218163 -0.955372
+ 1.728e+11Hz 0.217423 -0.955517
+ 1.729e+11Hz 0.216683 -0.955662
+ 1.73e+11Hz 0.215943 -0.955806
+ 1.731e+11Hz 0.215203 -0.955949
+ 1.732e+11Hz 0.214463 -0.956092
+ 1.733e+11Hz 0.213723 -0.956234
+ 1.734e+11Hz 0.212983 -0.956376
+ 1.735e+11Hz 0.212243 -0.956517
+ 1.736e+11Hz 0.211503 -0.956658
+ 1.737e+11Hz 0.210763 -0.956798
+ 1.738e+11Hz 0.210023 -0.956937
+ 1.739e+11Hz 0.209283 -0.957076
+ 1.74e+11Hz 0.208543 -0.957214
+ 1.741e+11Hz 0.207803 -0.957352
+ 1.742e+11Hz 0.207063 -0.957489
+ 1.743e+11Hz 0.206323 -0.957625
+ 1.744e+11Hz 0.205583 -0.957761
+ 1.745e+11Hz 0.204844 -0.957896
+ 1.746e+11Hz 0.204104 -0.958031
+ 1.747e+11Hz 0.203364 -0.958165
+ 1.748e+11Hz 0.202624 -0.958298
+ 1.749e+11Hz 0.201884 -0.958431
+ 1.75e+11Hz 0.201145 -0.958564
+ 1.751e+11Hz 0.200405 -0.958696
+ 1.752e+11Hz 0.199665 -0.958827
+ 1.753e+11Hz 0.198926 -0.958957
+ 1.754e+11Hz 0.198186 -0.959088
+ 1.755e+11Hz 0.197447 -0.959217
+ 1.756e+11Hz 0.196707 -0.959346
+ 1.757e+11Hz 0.195968 -0.959474
+ 1.758e+11Hz 0.195228 -0.959602
+ 1.759e+11Hz 0.194489 -0.95973
+ 1.76e+11Hz 0.19375 -0.959856
+ 1.761e+11Hz 0.19301 -0.959983
+ 1.762e+11Hz 0.192271 -0.960108
+ 1.763e+11Hz 0.191532 -0.960233
+ 1.764e+11Hz 0.190792 -0.960358
+ 1.765e+11Hz 0.190053 -0.960482
+ 1.766e+11Hz 0.189314 -0.960605
+ 1.767e+11Hz 0.188575 -0.960728
+ 1.768e+11Hz 0.187836 -0.96085
+ 1.769e+11Hz 0.187097 -0.960972
+ 1.77e+11Hz 0.186358 -0.961093
+ 1.771e+11Hz 0.185619 -0.961214
+ 1.772e+11Hz 0.18488 -0.961334
+ 1.773e+11Hz 0.184142 -0.961454
+ 1.774e+11Hz 0.183403 -0.961573
+ 1.775e+11Hz 0.182664 -0.961692
+ 1.776e+11Hz 0.181926 -0.96181
+ 1.777e+11Hz 0.181187 -0.961927
+ 1.778e+11Hz 0.180448 -0.962044
+ 1.779e+11Hz 0.17971 -0.962161
+ 1.78e+11Hz 0.178971 -0.962277
+ 1.781e+11Hz 0.178233 -0.962392
+ 1.782e+11Hz 0.177495 -0.962507
+ 1.783e+11Hz 0.176756 -0.962622
+ 1.784e+11Hz 0.176018 -0.962735
+ 1.785e+11Hz 0.17528 -0.962849
+ 1.786e+11Hz 0.174542 -0.962962
+ 1.787e+11Hz 0.173804 -0.963074
+ 1.788e+11Hz 0.173066 -0.963186
+ 1.789e+11Hz 0.172328 -0.963297
+ 1.79e+11Hz 0.17159 -0.963408
+ 1.791e+11Hz 0.170852 -0.963518
+ 1.792e+11Hz 0.170114 -0.963628
+ 1.793e+11Hz 0.169376 -0.963738
+ 1.794e+11Hz 0.168638 -0.963847
+ 1.795e+11Hz 0.167901 -0.963955
+ 1.796e+11Hz 0.167163 -0.964063
+ 1.797e+11Hz 0.166425 -0.96417
+ 1.798e+11Hz 0.165688 -0.964277
+ 1.799e+11Hz 0.16495 -0.964384
+ 1.8e+11Hz 0.164213 -0.96449
+ 1.801e+11Hz 0.163475 -0.964595
+ 1.802e+11Hz 0.162738 -0.9647
+ 1.803e+11Hz 0.162001 -0.964805
+ 1.804e+11Hz 0.161263 -0.964909
+ 1.805e+11Hz 0.160526 -0.965012
+ 1.806e+11Hz 0.159789 -0.965115
+ 1.807e+11Hz 0.159052 -0.965218
+ 1.808e+11Hz 0.158314 -0.96532
+ 1.809e+11Hz 0.157577 -0.965422
+ 1.81e+11Hz 0.15684 -0.965523
+ 1.811e+11Hz 0.156103 -0.965624
+ 1.812e+11Hz 0.155366 -0.965724
+ 1.813e+11Hz 0.154629 -0.965824
+ 1.814e+11Hz 0.153892 -0.965923
+ 1.815e+11Hz 0.153155 -0.966022
+ 1.816e+11Hz 0.152418 -0.966121
+ 1.817e+11Hz 0.151682 -0.966219
+ 1.818e+11Hz 0.150945 -0.966317
+ 1.819e+11Hz 0.150208 -0.966414
+ 1.82e+11Hz 0.149471 -0.96651
+ 1.821e+11Hz 0.148734 -0.966607
+ 1.822e+11Hz 0.147998 -0.966703
+ 1.823e+11Hz 0.147261 -0.966798
+ 1.824e+11Hz 0.146524 -0.966893
+ 1.825e+11Hz 0.145787 -0.966987
+ 1.826e+11Hz 0.145051 -0.967081
+ 1.827e+11Hz 0.144314 -0.967175
+ 1.828e+11Hz 0.143577 -0.967268
+ 1.829e+11Hz 0.142841 -0.967361
+ 1.83e+11Hz 0.142104 -0.967453
+ 1.831e+11Hz 0.141367 -0.967545
+ 1.832e+11Hz 0.140631 -0.967637
+ 1.833e+11Hz 0.139894 -0.967728
+ 1.834e+11Hz 0.139158 -0.967818
+ 1.835e+11Hz 0.138421 -0.967908
+ 1.836e+11Hz 0.137684 -0.967998
+ 1.837e+11Hz 0.136948 -0.968088
+ 1.838e+11Hz 0.136211 -0.968176
+ 1.839e+11Hz 0.135474 -0.968265
+ 1.84e+11Hz 0.134738 -0.968353
+ 1.841e+11Hz 0.134001 -0.968441
+ 1.842e+11Hz 0.133264 -0.968528
+ 1.843e+11Hz 0.132527 -0.968615
+ 1.844e+11Hz 0.131791 -0.968701
+ 1.845e+11Hz 0.131054 -0.968787
+ 1.846e+11Hz 0.130317 -0.968872
+ 1.847e+11Hz 0.12958 -0.968957
+ 1.848e+11Hz 0.128843 -0.969042
+ 1.849e+11Hz 0.128106 -0.969126
+ 1.85e+11Hz 0.127369 -0.96921
+ 1.851e+11Hz 0.126632 -0.969293
+ 1.852e+11Hz 0.125895 -0.969376
+ 1.853e+11Hz 0.125158 -0.969459
+ 1.854e+11Hz 0.124421 -0.969541
+ 1.855e+11Hz 0.123684 -0.969623
+ 1.856e+11Hz 0.122947 -0.969704
+ 1.857e+11Hz 0.12221 -0.969785
+ 1.858e+11Hz 0.121472 -0.969866
+ 1.859e+11Hz 0.120735 -0.969946
+ 1.86e+11Hz 0.119998 -0.970025
+ 1.861e+11Hz 0.11926 -0.970104
+ 1.862e+11Hz 0.118523 -0.970183
+ 1.863e+11Hz 0.117785 -0.970261
+ 1.864e+11Hz 0.117047 -0.970339
+ 1.865e+11Hz 0.11631 -0.970417
+ 1.866e+11Hz 0.115572 -0.970494
+ 1.867e+11Hz 0.114834 -0.970571
+ 1.868e+11Hz 0.114096 -0.970647
+ 1.869e+11Hz 0.113358 -0.970723
+ 1.87e+11Hz 0.11262 -0.970798
+ 1.871e+11Hz 0.111882 -0.970873
+ 1.872e+11Hz 0.111144 -0.970947
+ 1.873e+11Hz 0.110405 -0.971021
+ 1.874e+11Hz 0.109667 -0.971095
+ 1.875e+11Hz 0.108928 -0.971168
+ 1.876e+11Hz 0.10819 -0.971241
+ 1.877e+11Hz 0.107451 -0.971313
+ 1.878e+11Hz 0.106712 -0.971385
+ 1.879e+11Hz 0.105973 -0.971457
+ 1.88e+11Hz 0.105234 -0.971528
+ 1.881e+11Hz 0.104495 -0.971598
+ 1.882e+11Hz 0.103756 -0.971668
+ 1.883e+11Hz 0.103017 -0.971738
+ 1.884e+11Hz 0.102277 -0.971807
+ 1.885e+11Hz 0.101538 -0.971876
+ 1.886e+11Hz 0.100798 -0.971944
+ 1.887e+11Hz 0.100059 -0.972012
+ 1.888e+11Hz 0.0993189 -0.972079
+ 1.889e+11Hz 0.098579 -0.972146
+ 1.89e+11Hz 0.097839 -0.972213
+ 1.891e+11Hz 0.0970988 -0.972279
+ 1.892e+11Hz 0.0963586 -0.972344
+ 1.893e+11Hz 0.0956182 -0.97241
+ 1.894e+11Hz 0.0948777 -0.972474
+ 1.895e+11Hz 0.0941371 -0.972538
+ 1.896e+11Hz 0.0933963 -0.972602
+ 1.897e+11Hz 0.0926555 -0.972665
+ 1.898e+11Hz 0.0919145 -0.972728
+ 1.899e+11Hz 0.0911734 -0.97279
+ 1.9e+11Hz 0.0904321 -0.972852
+ 1.901e+11Hz 0.0896908 -0.972914
+ 1.902e+11Hz 0.0889493 -0.972974
+ 1.903e+11Hz 0.0882077 -0.973035
+ 1.904e+11Hz 0.0874659 -0.973095
+ 1.905e+11Hz 0.0867241 -0.973154
+ 1.906e+11Hz 0.0859821 -0.973213
+ 1.907e+11Hz 0.0852399 -0.973271
+ 1.908e+11Hz 0.0844977 -0.973329
+ 1.909e+11Hz 0.0837553 -0.973387
+ 1.91e+11Hz 0.0830128 -0.973444
+ 1.911e+11Hz 0.0822701 -0.9735
+ 1.912e+11Hz 0.0815273 -0.973556
+ 1.913e+11Hz 0.0807844 -0.973611
+ 1.914e+11Hz 0.0800413 -0.973666
+ 1.915e+11Hz 0.0792981 -0.97372
+ 1.916e+11Hz 0.0785548 -0.973774
+ 1.917e+11Hz 0.0778114 -0.973828
+ 1.918e+11Hz 0.0770678 -0.97388
+ 1.919e+11Hz 0.076324 -0.973933
+ 1.92e+11Hz 0.0755802 -0.973985
+ 1.921e+11Hz 0.0748362 -0.974036
+ 1.922e+11Hz 0.074092 -0.974086
+ 1.923e+11Hz 0.0733478 -0.974137
+ 1.924e+11Hz 0.0726034 -0.974186
+ 1.925e+11Hz 0.0718589 -0.974235
+ 1.926e+11Hz 0.0711142 -0.974284
+ 1.927e+11Hz 0.0703694 -0.974332
+ 1.928e+11Hz 0.0696245 -0.974379
+ 1.929e+11Hz 0.0688794 -0.974426
+ 1.93e+11Hz 0.0681342 -0.974473
+ 1.931e+11Hz 0.0673889 -0.974519
+ 1.932e+11Hz 0.0666435 -0.974564
+ 1.933e+11Hz 0.0658979 -0.974609
+ 1.934e+11Hz 0.0651522 -0.974653
+ 1.935e+11Hz 0.0644063 -0.974696
+ 1.936e+11Hz 0.0636604 -0.974739
+ 1.937e+11Hz 0.0629143 -0.974782
+ 1.938e+11Hz 0.0621681 -0.974824
+ 1.939e+11Hz 0.0614217 -0.974865
+ 1.94e+11Hz 0.0606753 -0.974906
+ 1.941e+11Hz 0.0599287 -0.974946
+ 1.942e+11Hz 0.059182 -0.974985
+ 1.943e+11Hz 0.0584352 -0.975025
+ 1.944e+11Hz 0.0576883 -0.975063
+ 1.945e+11Hz 0.0569412 -0.975101
+ 1.946e+11Hz 0.056194 -0.975138
+ 1.947e+11Hz 0.0554468 -0.975175
+ 1.948e+11Hz 0.0546994 -0.975211
+ 1.949e+11Hz 0.0539519 -0.975246
+ 1.95e+11Hz 0.0532043 -0.975281
+ 1.951e+11Hz 0.0524565 -0.975316
+ 1.952e+11Hz 0.0517087 -0.975349
+ 1.953e+11Hz 0.0509608 -0.975382
+ 1.954e+11Hz 0.0502128 -0.975415
+ 1.955e+11Hz 0.0494646 -0.975447
+ 1.956e+11Hz 0.0487164 -0.975478
+ 1.957e+11Hz 0.0479681 -0.975509
+ 1.958e+11Hz 0.0472196 -0.975539
+ 1.959e+11Hz 0.0464711 -0.975568
+ 1.96e+11Hz 0.0457225 -0.975597
+ 1.961e+11Hz 0.0449738 -0.975625
+ 1.962e+11Hz 0.044225 -0.975653
+ 1.963e+11Hz 0.0434761 -0.97568
+ 1.964e+11Hz 0.0427272 -0.975706
+ 1.965e+11Hz 0.0419781 -0.975732
+ 1.966e+11Hz 0.041229 -0.975757
+ 1.967e+11Hz 0.0404798 -0.975782
+ 1.968e+11Hz 0.0397305 -0.975806
+ 1.969e+11Hz 0.0389812 -0.975829
+ 1.97e+11Hz 0.0382317 -0.975852
+ 1.971e+11Hz 0.0374822 -0.975874
+ 1.972e+11Hz 0.0367327 -0.975895
+ 1.973e+11Hz 0.035983 -0.975916
+ 1.974e+11Hz 0.0352333 -0.975936
+ 1.975e+11Hz 0.0344836 -0.975955
+ 1.976e+11Hz 0.0337338 -0.975974
+ 1.977e+11Hz 0.0329839 -0.975992
+ 1.978e+11Hz 0.032234 -0.97601
+ 1.979e+11Hz 0.031484 -0.976027
+ 1.98e+11Hz 0.0307339 -0.976043
+ 1.981e+11Hz 0.0299839 -0.976059
+ 1.982e+11Hz 0.0292337 -0.976074
+ 1.983e+11Hz 0.0284836 -0.976088
+ 1.984e+11Hz 0.0277334 -0.976102
+ 1.985e+11Hz 0.0269831 -0.976115
+ 1.986e+11Hz 0.0262328 -0.976128
+ 1.987e+11Hz 0.0254825 -0.97614
+ 1.988e+11Hz 0.0247321 -0.976151
+ 1.989e+11Hz 0.0239817 -0.976161
+ 1.99e+11Hz 0.0232313 -0.976171
+ 1.991e+11Hz 0.0224809 -0.976181
+ 1.992e+11Hz 0.0217304 -0.976189
+ 1.993e+11Hz 0.0209799 -0.976197
+ 1.994e+11Hz 0.0202294 -0.976205
+ 1.995e+11Hz 0.0194789 -0.976211
+ 1.996e+11Hz 0.0187284 -0.976217
+ 1.997e+11Hz 0.0179778 -0.976223
+ 1.998e+11Hz 0.0172273 -0.976227
+ 1.999e+11Hz 0.0164767 -0.976232
+ 2e+11Hz 0.0157261 -0.976235
+ 2.001e+11Hz 0.0149755 -0.976238
+ 2.002e+11Hz 0.014225 -0.97624
+ 2.003e+11Hz 0.0134744 -0.976242
+ 2.004e+11Hz 0.0127238 -0.976242
+ 2.005e+11Hz 0.0119732 -0.976243
+ 2.006e+11Hz 0.0112227 -0.976242
+ 2.007e+11Hz 0.0104721 -0.976241
+ 2.008e+11Hz 0.00972156 -0.97624
+ 2.009e+11Hz 0.00897103 -0.976237
+ 2.01e+11Hz 0.00822051 -0.976234
+ 2.011e+11Hz 0.00747001 -0.976231
+ 2.012e+11Hz 0.00671953 -0.976226
+ 2.013e+11Hz 0.00596907 -0.976222
+ 2.014e+11Hz 0.00521864 -0.976216
+ 2.015e+11Hz 0.00446823 -0.97621
+ 2.016e+11Hz 0.00371784 -0.976203
+ 2.017e+11Hz 0.00296749 -0.976196
+ 2.018e+11Hz 0.00221717 -0.976187
+ 2.019e+11Hz 0.00146688 -0.976179
+ 2.02e+11Hz 0.00071662 -0.976169
+ 2.021e+11Hz -3.35995e-05 -0.976159
+ 2.022e+11Hz -0.00078378 -0.976149
+ 2.023e+11Hz -0.00153392 -0.976137
+ 2.024e+11Hz -0.00228402 -0.976125
+ 2.025e+11Hz -0.00303408 -0.976113
+ 2.026e+11Hz -0.00378409 -0.9761
+ 2.027e+11Hz -0.00453405 -0.976086
+ 2.028e+11Hz -0.00528396 -0.976071
+ 2.029e+11Hz -0.00603383 -0.976056
+ 2.03e+11Hz -0.00678364 -0.97604
+ 2.031e+11Hz -0.0075334 -0.976024
+ 2.032e+11Hz -0.0082831 -0.976007
+ 2.033e+11Hz -0.00903275 -0.975989
+ 2.034e+11Hz -0.00978234 -0.975971
+ 2.035e+11Hz -0.0105319 -0.975952
+ 2.036e+11Hz -0.0112813 -0.975933
+ 2.037e+11Hz -0.0120307 -0.975913
+ 2.038e+11Hz -0.0127801 -0.975892
+ 2.039e+11Hz -0.0135294 -0.97587
+ 2.04e+11Hz -0.0142786 -0.975848
+ 2.041e+11Hz -0.0150277 -0.975826
+ 2.042e+11Hz -0.0157768 -0.975802
+ 2.043e+11Hz -0.0165258 -0.975779
+ 2.044e+11Hz -0.0172747 -0.975754
+ 2.045e+11Hz -0.0180236 -0.975729
+ 2.046e+11Hz -0.0187723 -0.975703
+ 2.047e+11Hz -0.019521 -0.975677
+ 2.048e+11Hz -0.0202697 -0.97565
+ 2.049e+11Hz -0.0210182 -0.975622
+ 2.05e+11Hz -0.0217667 -0.975594
+ 2.051e+11Hz -0.0225151 -0.975565
+ 2.052e+11Hz -0.0232634 -0.975536
+ 2.053e+11Hz -0.0240116 -0.975506
+ 2.054e+11Hz -0.0247597 -0.975475
+ 2.055e+11Hz -0.0255078 -0.975444
+ 2.056e+11Hz -0.0262557 -0.975412
+ 2.057e+11Hz -0.0270036 -0.975379
+ 2.058e+11Hz -0.0277514 -0.975346
+ 2.059e+11Hz -0.0284991 -0.975312
+ 2.06e+11Hz -0.0292467 -0.975278
+ 2.061e+11Hz -0.0299942 -0.975243
+ 2.062e+11Hz -0.0307416 -0.975208
+ 2.063e+11Hz -0.0314889 -0.975171
+ 2.064e+11Hz -0.0322361 -0.975135
+ 2.065e+11Hz -0.0329833 -0.975097
+ 2.066e+11Hz -0.0337303 -0.975059
+ 2.067e+11Hz -0.0344772 -0.975021
+ 2.068e+11Hz -0.0352241 -0.974982
+ 2.069e+11Hz -0.0359708 -0.974942
+ 2.07e+11Hz -0.0367175 -0.974901
+ 2.071e+11Hz -0.037464 -0.97486
+ 2.072e+11Hz -0.0382104 -0.974819
+ 2.073e+11Hz -0.0389567 -0.974777
+ 2.074e+11Hz -0.039703 -0.974734
+ 2.075e+11Hz -0.0404491 -0.974691
+ 2.076e+11Hz -0.0411951 -0.974647
+ 2.077e+11Hz -0.041941 -0.974602
+ 2.078e+11Hz -0.0426868 -0.974557
+ 2.079e+11Hz -0.0434324 -0.974511
+ 2.08e+11Hz -0.044178 -0.974465
+ 2.081e+11Hz -0.0449235 -0.974418
+ 2.082e+11Hz -0.0456688 -0.97437
+ 2.083e+11Hz -0.046414 -0.974322
+ 2.084e+11Hz -0.0471591 -0.974274
+ 2.085e+11Hz -0.0479041 -0.974224
+ 2.086e+11Hz -0.048649 -0.974174
+ 2.087e+11Hz -0.0493938 -0.974124
+ 2.088e+11Hz -0.0501384 -0.974073
+ 2.089e+11Hz -0.050883 -0.974021
+ 2.09e+11Hz -0.0516274 -0.973969
+ 2.091e+11Hz -0.0523716 -0.973916
+ 2.092e+11Hz -0.0531158 -0.973863
+ 2.093e+11Hz -0.0538598 -0.973809
+ 2.094e+11Hz -0.0546038 -0.973754
+ 2.095e+11Hz -0.0553475 -0.973699
+ 2.096e+11Hz -0.0560912 -0.973644
+ 2.097e+11Hz -0.0568347 -0.973587
+ 2.098e+11Hz -0.0575781 -0.97353
+ 2.099e+11Hz -0.0583214 -0.973473
+ 2.1e+11Hz -0.0590646 -0.973415
+ 2.101e+11Hz -0.0598076 -0.973356
+ 2.102e+11Hz -0.0605504 -0.973297
+ 2.103e+11Hz -0.0612932 -0.973237
+ 2.104e+11Hz -0.0620358 -0.973177
+ 2.105e+11Hz -0.0627783 -0.973116
+ 2.106e+11Hz -0.0635206 -0.973055
+ 2.107e+11Hz -0.0642628 -0.972992
+ 2.108e+11Hz -0.0650049 -0.97293
+ 2.109e+11Hz -0.0657468 -0.972867
+ 2.11e+11Hz -0.0664885 -0.972803
+ 2.111e+11Hz -0.0672302 -0.972739
+ 2.112e+11Hz -0.0679717 -0.972674
+ 2.113e+11Hz -0.068713 -0.972608
+ 2.114e+11Hz -0.0694542 -0.972542
+ 2.115e+11Hz -0.0701952 -0.972475
+ 2.116e+11Hz -0.0709361 -0.972408
+ 2.117e+11Hz -0.0716769 -0.97234
+ 2.118e+11Hz -0.0724175 -0.972272
+ 2.119e+11Hz -0.0731579 -0.972203
+ 2.12e+11Hz -0.0738982 -0.972134
+ 2.121e+11Hz -0.0746383 -0.972064
+ 2.122e+11Hz -0.0753783 -0.971993
+ 2.123e+11Hz -0.0761181 -0.971922
+ 2.124e+11Hz -0.0768577 -0.97185
+ 2.125e+11Hz -0.0775972 -0.971778
+ 2.126e+11Hz -0.0783366 -0.971705
+ 2.127e+11Hz -0.0790757 -0.971632
+ 2.128e+11Hz -0.0798147 -0.971558
+ 2.129e+11Hz -0.0805536 -0.971484
+ 2.13e+11Hz -0.0812922 -0.971409
+ 2.131e+11Hz -0.0820307 -0.971333
+ 2.132e+11Hz -0.0827691 -0.971257
+ 2.133e+11Hz -0.0835072 -0.97118
+ 2.134e+11Hz -0.0842452 -0.971103
+ 2.135e+11Hz -0.084983 -0.971026
+ 2.136e+11Hz -0.0857206 -0.970947
+ 2.137e+11Hz -0.0864581 -0.970868
+ 2.138e+11Hz -0.0871954 -0.970789
+ 2.139e+11Hz -0.0879325 -0.970709
+ 2.14e+11Hz -0.0886694 -0.970629
+ 2.141e+11Hz -0.0894061 -0.970548
+ 2.142e+11Hz -0.0901427 -0.970466
+ 2.143e+11Hz -0.090879 -0.970384
+ 2.144e+11Hz -0.0916152 -0.970302
+ 2.145e+11Hz -0.0923512 -0.970219
+ 2.146e+11Hz -0.093087 -0.970135
+ 2.147e+11Hz -0.0938226 -0.970051
+ 2.148e+11Hz -0.0945581 -0.969966
+ 2.149e+11Hz -0.0952933 -0.969881
+ 2.15e+11Hz -0.0960283 -0.969795
+ 2.151e+11Hz -0.0967632 -0.969709
+ 2.152e+11Hz -0.0974978 -0.969622
+ 2.153e+11Hz -0.0982323 -0.969535
+ 2.154e+11Hz -0.0989665 -0.969447
+ 2.155e+11Hz -0.0997006 -0.969359
+ 2.156e+11Hz -0.100434 -0.96927
+ 2.157e+11Hz -0.101168 -0.969181
+ 2.158e+11Hz -0.101902 -0.969091
+ 2.159e+11Hz -0.102635 -0.969001
+ 2.16e+11Hz -0.103368 -0.96891
+ 2.161e+11Hz -0.104101 -0.968819
+ 2.162e+11Hz -0.104833 -0.968727
+ 2.163e+11Hz -0.105566 -0.968635
+ 2.164e+11Hz -0.106298 -0.968542
+ 2.165e+11Hz -0.10703 -0.968449
+ 2.166e+11Hz -0.107762 -0.968355
+ 2.167e+11Hz -0.108493 -0.968261
+ 2.168e+11Hz -0.109225 -0.968166
+ 2.169e+11Hz -0.109956 -0.968071
+ 2.17e+11Hz -0.110687 -0.967976
+ 2.171e+11Hz -0.111418 -0.96788
+ 2.172e+11Hz -0.112148 -0.967783
+ 2.173e+11Hz -0.112878 -0.967686
+ 2.174e+11Hz -0.113608 -0.967589
+ 2.175e+11Hz -0.114338 -0.967491
+ 2.176e+11Hz -0.115068 -0.967392
+ 2.177e+11Hz -0.115797 -0.967294
+ 2.178e+11Hz -0.116527 -0.967194
+ 2.179e+11Hz -0.117256 -0.967095
+ 2.18e+11Hz -0.117984 -0.966995
+ 2.181e+11Hz -0.118713 -0.966894
+ 2.182e+11Hz -0.119441 -0.966793
+ 2.183e+11Hz -0.12017 -0.966691
+ 2.184e+11Hz -0.120898 -0.96659
+ 2.185e+11Hz -0.121625 -0.966487
+ 2.186e+11Hz -0.122353 -0.966385
+ 2.187e+11Hz -0.12308 -0.966281
+ 2.188e+11Hz -0.123807 -0.966178
+ 2.189e+11Hz -0.124534 -0.966074
+ 2.19e+11Hz -0.125261 -0.96597
+ 2.191e+11Hz -0.125987 -0.965865
+ 2.192e+11Hz -0.126713 -0.96576
+ 2.193e+11Hz -0.127439 -0.965654
+ 2.194e+11Hz -0.128165 -0.965548
+ 2.195e+11Hz -0.128891 -0.965442
+ 2.196e+11Hz -0.129616 -0.965335
+ 2.197e+11Hz -0.130341 -0.965228
+ 2.198e+11Hz -0.131066 -0.96512
+ 2.199e+11Hz -0.131791 -0.965012
+ 2.2e+11Hz -0.132516 -0.964904
+ 2.201e+11Hz -0.13324 -0.964795
+ 2.202e+11Hz -0.133964 -0.964686
+ 2.203e+11Hz -0.134688 -0.964577
+ 2.204e+11Hz -0.135412 -0.964467
+ 2.205e+11Hz -0.136136 -0.964357
+ 2.206e+11Hz -0.136859 -0.964247
+ 2.207e+11Hz -0.137582 -0.964136
+ 2.208e+11Hz -0.138305 -0.964025
+ 2.209e+11Hz -0.139028 -0.963913
+ 2.21e+11Hz -0.139751 -0.963801
+ 2.211e+11Hz -0.140473 -0.963689
+ 2.212e+11Hz -0.141195 -0.963576
+ 2.213e+11Hz -0.141917 -0.963464
+ 2.214e+11Hz -0.142639 -0.96335
+ 2.215e+11Hz -0.143361 -0.963237
+ 2.216e+11Hz -0.144083 -0.963123
+ 2.217e+11Hz -0.144804 -0.963009
+ 2.218e+11Hz -0.145525 -0.962894
+ 2.219e+11Hz -0.146246 -0.96278
+ 2.22e+11Hz -0.146967 -0.962665
+ 2.221e+11Hz -0.147688 -0.962549
+ 2.222e+11Hz -0.148409 -0.962433
+ 2.223e+11Hz -0.149129 -0.962317
+ 2.224e+11Hz -0.149849 -0.962201
+ 2.225e+11Hz -0.15057 -0.962085
+ 2.226e+11Hz -0.15129 -0.961968
+ 2.227e+11Hz -0.152009 -0.96185
+ 2.228e+11Hz -0.152729 -0.961733
+ 2.229e+11Hz -0.153449 -0.961615
+ 2.23e+11Hz -0.154168 -0.961497
+ 2.231e+11Hz -0.154888 -0.961379
+ 2.232e+11Hz -0.155607 -0.96126
+ 2.233e+11Hz -0.156326 -0.961141
+ 2.234e+11Hz -0.157045 -0.961022
+ 2.235e+11Hz -0.157764 -0.960903
+ 2.236e+11Hz -0.158483 -0.960783
+ 2.237e+11Hz -0.159202 -0.960663
+ 2.238e+11Hz -0.15992 -0.960543
+ 2.239e+11Hz -0.160639 -0.960422
+ 2.24e+11Hz -0.161357 -0.960302
+ 2.241e+11Hz -0.162076 -0.960181
+ 2.242e+11Hz -0.162794 -0.960059
+ 2.243e+11Hz -0.163512 -0.959938
+ 2.244e+11Hz -0.16423 -0.959816
+ 2.245e+11Hz -0.164948 -0.959694
+ 2.246e+11Hz -0.165667 -0.959572
+ 2.247e+11Hz -0.166385 -0.959449
+ 2.248e+11Hz -0.167102 -0.959326
+ 2.249e+11Hz -0.16782 -0.959203
+ 2.25e+11Hz -0.168538 -0.95908
+ 2.251e+11Hz -0.169256 -0.958956
+ 2.252e+11Hz -0.169974 -0.958832
+ 2.253e+11Hz -0.170692 -0.958708
+ 2.254e+11Hz -0.17141 -0.958584
+ 2.255e+11Hz -0.172127 -0.958459
+ 2.256e+11Hz -0.172845 -0.958335
+ 2.257e+11Hz -0.173563 -0.95821
+ 2.258e+11Hz -0.174281 -0.958084
+ 2.259e+11Hz -0.174999 -0.957959
+ 2.26e+11Hz -0.175716 -0.957833
+ 2.261e+11Hz -0.176434 -0.957707
+ 2.262e+11Hz -0.177152 -0.95758
+ 2.263e+11Hz -0.17787 -0.957454
+ 2.264e+11Hz -0.178588 -0.957327
+ 2.265e+11Hz -0.179306 -0.9572
+ 2.266e+11Hz -0.180024 -0.957073
+ 2.267e+11Hz -0.180742 -0.956945
+ 2.268e+11Hz -0.18146 -0.956817
+ 2.269e+11Hz -0.182178 -0.956689
+ 2.27e+11Hz -0.182897 -0.956561
+ 2.271e+11Hz -0.183615 -0.956432
+ 2.272e+11Hz -0.184333 -0.956303
+ 2.273e+11Hz -0.185052 -0.956174
+ 2.274e+11Hz -0.18577 -0.956044
+ 2.275e+11Hz -0.186489 -0.955915
+ 2.276e+11Hz -0.187208 -0.955785
+ 2.277e+11Hz -0.187927 -0.955655
+ 2.278e+11Hz -0.188646 -0.955524
+ 2.279e+11Hz -0.189365 -0.955393
+ 2.28e+11Hz -0.190084 -0.955262
+ 2.281e+11Hz -0.190804 -0.955131
+ 2.282e+11Hz -0.191523 -0.954999
+ 2.283e+11Hz -0.192243 -0.954867
+ 2.284e+11Hz -0.192963 -0.954735
+ 2.285e+11Hz -0.193683 -0.954602
+ 2.286e+11Hz -0.194403 -0.954469
+ 2.287e+11Hz -0.195123 -0.954336
+ 2.288e+11Hz -0.195844 -0.954203
+ 2.289e+11Hz -0.196564 -0.954069
+ 2.29e+11Hz -0.197285 -0.953935
+ 2.291e+11Hz -0.198006 -0.9538
+ 2.292e+11Hz -0.198727 -0.953665
+ 2.293e+11Hz -0.199449 -0.95353
+ 2.294e+11Hz -0.20017 -0.953395
+ 2.295e+11Hz -0.200892 -0.953259
+ 2.296e+11Hz -0.201614 -0.953123
+ 2.297e+11Hz -0.202336 -0.952986
+ 2.298e+11Hz -0.203058 -0.952849
+ 2.299e+11Hz -0.203781 -0.952712
+ 2.3e+11Hz -0.204504 -0.952575
+ 2.301e+11Hz -0.205227 -0.952437
+ 2.302e+11Hz -0.20595 -0.952298
+ 2.303e+11Hz -0.206673 -0.952159
+ 2.304e+11Hz -0.207397 -0.95202
+ 2.305e+11Hz -0.208121 -0.951881
+ 2.306e+11Hz -0.208845 -0.951741
+ 2.307e+11Hz -0.209569 -0.951601
+ 2.308e+11Hz -0.210294 -0.95146
+ 2.309e+11Hz -0.211019 -0.951319
+ 2.31e+11Hz -0.211744 -0.951177
+ 2.311e+11Hz -0.212469 -0.951035
+ 2.312e+11Hz -0.213195 -0.950893
+ 2.313e+11Hz -0.213921 -0.95075
+ 2.314e+11Hz -0.214647 -0.950606
+ 2.315e+11Hz -0.215374 -0.950462
+ 2.316e+11Hz -0.2161 -0.950318
+ 2.317e+11Hz -0.216827 -0.950173
+ 2.318e+11Hz -0.217554 -0.950028
+ 2.319e+11Hz -0.218282 -0.949883
+ 2.32e+11Hz -0.21901 -0.949736
+ 2.321e+11Hz -0.219738 -0.94959
+ 2.322e+11Hz -0.220466 -0.949442
+ 2.323e+11Hz -0.221195 -0.949295
+ 2.324e+11Hz -0.221923 -0.949146
+ 2.325e+11Hz -0.222653 -0.948998
+ 2.326e+11Hz -0.223382 -0.948848
+ 2.327e+11Hz -0.224112 -0.948699
+ 2.328e+11Hz -0.224842 -0.948548
+ 2.329e+11Hz -0.225572 -0.948397
+ 2.33e+11Hz -0.226302 -0.948246
+ 2.331e+11Hz -0.227033 -0.948094
+ 2.332e+11Hz -0.227764 -0.947941
+ 2.333e+11Hz -0.228495 -0.947788
+ 2.334e+11Hz -0.229227 -0.947634
+ 2.335e+11Hz -0.229959 -0.947479
+ 2.336e+11Hz -0.230691 -0.947324
+ 2.337e+11Hz -0.231424 -0.947169
+ 2.338e+11Hz -0.232156 -0.947012
+ 2.339e+11Hz -0.232889 -0.946855
+ 2.34e+11Hz -0.233623 -0.946698
+ 2.341e+11Hz -0.234356 -0.94654
+ 2.342e+11Hz -0.23509 -0.946381
+ 2.343e+11Hz -0.235824 -0.946221
+ 2.344e+11Hz -0.236558 -0.946061
+ 2.345e+11Hz -0.237293 -0.9459
+ 2.346e+11Hz -0.238028 -0.945739
+ 2.347e+11Hz -0.238763 -0.945577
+ 2.348e+11Hz -0.239498 -0.945414
+ 2.349e+11Hz -0.240234 -0.94525
+ 2.35e+11Hz -0.240969 -0.945086
+ 2.351e+11Hz -0.241706 -0.944921
+ 2.352e+11Hz -0.242442 -0.944755
+ 2.353e+11Hz -0.243178 -0.944589
+ 2.354e+11Hz -0.243915 -0.944421
+ 2.355e+11Hz -0.244652 -0.944253
+ 2.356e+11Hz -0.245389 -0.944085
+ 2.357e+11Hz -0.246127 -0.943915
+ 2.358e+11Hz -0.246865 -0.943745
+ 2.359e+11Hz -0.247602 -0.943574
+ 2.36e+11Hz -0.248341 -0.943402
+ 2.361e+11Hz -0.249079 -0.94323
+ 2.362e+11Hz -0.249817 -0.943057
+ 2.363e+11Hz -0.250556 -0.942882
+ 2.364e+11Hz -0.251295 -0.942708
+ 2.365e+11Hz -0.252034 -0.942532
+ 2.366e+11Hz -0.252773 -0.942355
+ 2.367e+11Hz -0.253513 -0.942178
+ 2.368e+11Hz -0.254252 -0.942
+ 2.369e+11Hz -0.254992 -0.941821
+ 2.37e+11Hz -0.255732 -0.941641
+ 2.371e+11Hz -0.256472 -0.94146
+ 2.372e+11Hz -0.257212 -0.941279
+ 2.373e+11Hz -0.257952 -0.941096
+ 2.374e+11Hz -0.258693 -0.940913
+ 2.375e+11Hz -0.259433 -0.940729
+ 2.376e+11Hz -0.260174 -0.940544
+ 2.377e+11Hz -0.260915 -0.940359
+ 2.378e+11Hz -0.261656 -0.940172
+ 2.379e+11Hz -0.262397 -0.939984
+ 2.38e+11Hz -0.263138 -0.939796
+ 2.381e+11Hz -0.263879 -0.939607
+ 2.382e+11Hz -0.26462 -0.939417
+ 2.383e+11Hz -0.265362 -0.939225
+ 2.384e+11Hz -0.266103 -0.939034
+ 2.385e+11Hz -0.266845 -0.938841
+ 2.386e+11Hz -0.267586 -0.938647
+ 2.387e+11Hz -0.268328 -0.938452
+ 2.388e+11Hz -0.269069 -0.938257
+ 2.389e+11Hz -0.269811 -0.93806
+ 2.39e+11Hz -0.270553 -0.937863
+ 2.391e+11Hz -0.271294 -0.937665
+ 2.392e+11Hz -0.272036 -0.937465
+ 2.393e+11Hz -0.272778 -0.937265
+ 2.394e+11Hz -0.273519 -0.937064
+ 2.395e+11Hz -0.274261 -0.936862
+ 2.396e+11Hz -0.275003 -0.936659
+ 2.397e+11Hz -0.275744 -0.936456
+ 2.398e+11Hz -0.276486 -0.936251
+ 2.399e+11Hz -0.277227 -0.936045
+ 2.4e+11Hz -0.277969 -0.935839
+ 2.401e+11Hz -0.27871 -0.935631
+ 2.402e+11Hz -0.279451 -0.935423
+ 2.403e+11Hz -0.280193 -0.935213
+ 2.404e+11Hz -0.280934 -0.935003
+ 2.405e+11Hz -0.281675 -0.934792
+ 2.406e+11Hz -0.282416 -0.93458
+ 2.407e+11Hz -0.283157 -0.934367
+ 2.408e+11Hz -0.283898 -0.934153
+ 2.409e+11Hz -0.284638 -0.933938
+ 2.41e+11Hz -0.285379 -0.933722
+ 2.411e+11Hz -0.286119 -0.933505
+ 2.412e+11Hz -0.286859 -0.933287
+ 2.413e+11Hz -0.287599 -0.933069
+ 2.414e+11Hz -0.288339 -0.932849
+ 2.415e+11Hz -0.289079 -0.932629
+ 2.416e+11Hz -0.289819 -0.932407
+ 2.417e+11Hz -0.290558 -0.932185
+ 2.418e+11Hz -0.291297 -0.931962
+ 2.419e+11Hz -0.292036 -0.931737
+ 2.42e+11Hz -0.292775 -0.931512
+ 2.421e+11Hz -0.293514 -0.931286
+ 2.422e+11Hz -0.294252 -0.931059
+ 2.423e+11Hz -0.29499 -0.930832
+ 2.424e+11Hz -0.295728 -0.930603
+ 2.425e+11Hz -0.296466 -0.930373
+ 2.426e+11Hz -0.297203 -0.930143
+ 2.427e+11Hz -0.29794 -0.929911
+ 2.428e+11Hz -0.298677 -0.929679
+ 2.429e+11Hz -0.299414 -0.929446
+ 2.43e+11Hz -0.30015 -0.929212
+ 2.431e+11Hz -0.300887 -0.928977
+ 2.432e+11Hz -0.301622 -0.928741
+ 2.433e+11Hz -0.302358 -0.928504
+ 2.434e+11Hz -0.303093 -0.928267
+ 2.435e+11Hz -0.303828 -0.928028
+ 2.436e+11Hz -0.304563 -0.927789
+ 2.437e+11Hz -0.305297 -0.927549
+ 2.438e+11Hz -0.306031 -0.927308
+ 2.439e+11Hz -0.306765 -0.927066
+ 2.44e+11Hz -0.307498 -0.926823
+ 2.441e+11Hz -0.308231 -0.926579
+ 2.442e+11Hz -0.308964 -0.926335
+ 2.443e+11Hz -0.309697 -0.92609
+ 2.444e+11Hz -0.310429 -0.925844
+ 2.445e+11Hz -0.31116 -0.925597
+ 2.446e+11Hz -0.311892 -0.925349
+ 2.447e+11Hz -0.312623 -0.925101
+ 2.448e+11Hz -0.313353 -0.924851
+ 2.449e+11Hz -0.314083 -0.924601
+ 2.45e+11Hz -0.314813 -0.92435
+ 2.451e+11Hz -0.315543 -0.924099
+ 2.452e+11Hz -0.316272 -0.923846
+ 2.453e+11Hz -0.317001 -0.923593
+ 2.454e+11Hz -0.317729 -0.923339
+ 2.455e+11Hz -0.318457 -0.923084
+ 2.456e+11Hz -0.319185 -0.922828
+ 2.457e+11Hz -0.319912 -0.922572
+ 2.458e+11Hz -0.320639 -0.922315
+ 2.459e+11Hz -0.321365 -0.922057
+ 2.46e+11Hz -0.322091 -0.921798
+ 2.461e+11Hz -0.322817 -0.921539
+ 2.462e+11Hz -0.323542 -0.921279
+ 2.463e+11Hz -0.324267 -0.921018
+ 2.464e+11Hz -0.324991 -0.920756
+ 2.465e+11Hz -0.325715 -0.920494
+ 2.466e+11Hz -0.326439 -0.920231
+ 2.467e+11Hz -0.327162 -0.919968
+ 2.468e+11Hz -0.327884 -0.919703
+ 2.469e+11Hz -0.328607 -0.919438
+ 2.47e+11Hz -0.329329 -0.919172
+ 2.471e+11Hz -0.33005 -0.918906
+ 2.472e+11Hz -0.330771 -0.918639
+ 2.473e+11Hz -0.331492 -0.918371
+ 2.474e+11Hz -0.332212 -0.918103
+ 2.475e+11Hz -0.332932 -0.917833
+ 2.476e+11Hz -0.333651 -0.917564
+ 2.477e+11Hz -0.33437 -0.917293
+ 2.478e+11Hz -0.335089 -0.917022
+ 2.479e+11Hz -0.335807 -0.91675
+ 2.48e+11Hz -0.336524 -0.916478
+ 2.481e+11Hz -0.337242 -0.916205
+ 2.482e+11Hz -0.337958 -0.915931
+ 2.483e+11Hz -0.338675 -0.915657
+ 2.484e+11Hz -0.339391 -0.915382
+ 2.485e+11Hz -0.340106 -0.915107
+ 2.486e+11Hz -0.340821 -0.914831
+ 2.487e+11Hz -0.341536 -0.914554
+ 2.488e+11Hz -0.342251 -0.914277
+ 2.489e+11Hz -0.342964 -0.913999
+ 2.49e+11Hz -0.343678 -0.91372
+ 2.491e+11Hz -0.344391 -0.913441
+ 2.492e+11Hz -0.345104 -0.913162
+ 2.493e+11Hz -0.345816 -0.912881
+ 2.494e+11Hz -0.346528 -0.912601
+ 2.495e+11Hz -0.347239 -0.912319
+ 2.496e+11Hz -0.34795 -0.912037
+ 2.497e+11Hz -0.348661 -0.911755
+ 2.498e+11Hz -0.349371 -0.911472
+ 2.499e+11Hz -0.350081 -0.911188
+ 2.5e+11Hz -0.35079 -0.910904
+ 2.501e+11Hz -0.351499 -0.910619
+ 2.502e+11Hz -0.352208 -0.910334
+ 2.503e+11Hz -0.352916 -0.910048
+ 2.504e+11Hz -0.353624 -0.909762
+ 2.505e+11Hz -0.354332 -0.909475
+ 2.506e+11Hz -0.355039 -0.909187
+ 2.507e+11Hz -0.355745 -0.908899
+ 2.508e+11Hz -0.356452 -0.908611
+ 2.509e+11Hz -0.357158 -0.908322
+ 2.51e+11Hz -0.357863 -0.908032
+ 2.511e+11Hz -0.358568 -0.907742
+ 2.512e+11Hz -0.359273 -0.907452
+ 2.513e+11Hz -0.359978 -0.907161
+ 2.514e+11Hz -0.360682 -0.906869
+ 2.515e+11Hz -0.361386 -0.906577
+ 2.516e+11Hz -0.362089 -0.906284
+ 2.517e+11Hz -0.362792 -0.905991
+ 2.518e+11Hz -0.363495 -0.905697
+ 2.519e+11Hz -0.364197 -0.905403
+ 2.52e+11Hz -0.364899 -0.905108
+ 2.521e+11Hz -0.3656 -0.904813
+ 2.522e+11Hz -0.366302 -0.904517
+ 2.523e+11Hz -0.367003 -0.904221
+ 2.524e+11Hz -0.367703 -0.903924
+ 2.525e+11Hz -0.368404 -0.903627
+ 2.526e+11Hz -0.369103 -0.903329
+ 2.527e+11Hz -0.369803 -0.903031
+ 2.528e+11Hz -0.370502 -0.902732
+ 2.529e+11Hz -0.371201 -0.902433
+ 2.53e+11Hz -0.3719 -0.902133
+ 2.531e+11Hz -0.372598 -0.901833
+ 2.532e+11Hz -0.373296 -0.901532
+ 2.533e+11Hz -0.373994 -0.901231
+ 2.534e+11Hz -0.374691 -0.900929
+ 2.535e+11Hz -0.375388 -0.900627
+ 2.536e+11Hz -0.376085 -0.900324
+ 2.537e+11Hz -0.376781 -0.90002
+ 2.538e+11Hz -0.377477 -0.899717
+ 2.539e+11Hz -0.378173 -0.899412
+ 2.54e+11Hz -0.378868 -0.899107
+ 2.541e+11Hz -0.379564 -0.898802
+ 2.542e+11Hz -0.380258 -0.898496
+ 2.543e+11Hz -0.380953 -0.89819
+ 2.544e+11Hz -0.381647 -0.897883
+ 2.545e+11Hz -0.382341 -0.897575
+ 2.546e+11Hz -0.383035 -0.897267
+ 2.547e+11Hz -0.383728 -0.896959
+ 2.548e+11Hz -0.384421 -0.89665
+ 2.549e+11Hz -0.385114 -0.89634
+ 2.55e+11Hz -0.385806 -0.89603
+ 2.551e+11Hz -0.386498 -0.89572
+ 2.552e+11Hz -0.38719 -0.895409
+ 2.553e+11Hz -0.387882 -0.895097
+ 2.554e+11Hz -0.388573 -0.894785
+ 2.555e+11Hz -0.389264 -0.894472
+ 2.556e+11Hz -0.389955 -0.894159
+ 2.557e+11Hz -0.390645 -0.893845
+ 2.558e+11Hz -0.391335 -0.893531
+ 2.559e+11Hz -0.392025 -0.893216
+ 2.56e+11Hz -0.392715 -0.892901
+ 2.561e+11Hz -0.393404 -0.892585
+ 2.562e+11Hz -0.394093 -0.892269
+ 2.563e+11Hz -0.394782 -0.891952
+ 2.564e+11Hz -0.39547 -0.891634
+ 2.565e+11Hz -0.396158 -0.891316
+ 2.566e+11Hz -0.396846 -0.890997
+ 2.567e+11Hz -0.397533 -0.890678
+ 2.568e+11Hz -0.39822 -0.890359
+ 2.569e+11Hz -0.398907 -0.890038
+ 2.57e+11Hz -0.399594 -0.889717
+ 2.571e+11Hz -0.40028 -0.889396
+ 2.572e+11Hz -0.400966 -0.889074
+ 2.573e+11Hz -0.401652 -0.888751
+ 2.574e+11Hz -0.402337 -0.888428
+ 2.575e+11Hz -0.403022 -0.888105
+ 2.576e+11Hz -0.403707 -0.88778
+ 2.577e+11Hz -0.404391 -0.887456
+ 2.578e+11Hz -0.405075 -0.88713
+ 2.579e+11Hz -0.405759 -0.886804
+ 2.58e+11Hz -0.406442 -0.886478
+ 2.581e+11Hz -0.407125 -0.886151
+ 2.582e+11Hz -0.407808 -0.885823
+ 2.583e+11Hz -0.408491 -0.885495
+ 2.584e+11Hz -0.409173 -0.885166
+ 2.585e+11Hz -0.409855 -0.884837
+ 2.586e+11Hz -0.410536 -0.884507
+ 2.587e+11Hz -0.411217 -0.884176
+ 2.588e+11Hz -0.411898 -0.883845
+ 2.589e+11Hz -0.412578 -0.883513
+ 2.59e+11Hz -0.413258 -0.883181
+ 2.591e+11Hz -0.413938 -0.882848
+ 2.592e+11Hz -0.414617 -0.882515
+ 2.593e+11Hz -0.415296 -0.882181
+ 2.594e+11Hz -0.415975 -0.881846
+ 2.595e+11Hz -0.416653 -0.881511
+ 2.596e+11Hz -0.417331 -0.881175
+ 2.597e+11Hz -0.418009 -0.880839
+ 2.598e+11Hz -0.418686 -0.880502
+ 2.599e+11Hz -0.419363 -0.880164
+ 2.6e+11Hz -0.420039 -0.879826
+ 2.601e+11Hz -0.420715 -0.879487
+ 2.602e+11Hz -0.42139 -0.879148
+ 2.603e+11Hz -0.422066 -0.878808
+ 2.604e+11Hz -0.42274 -0.878468
+ 2.605e+11Hz -0.423415 -0.878127
+ 2.606e+11Hz -0.424089 -0.877785
+ 2.607e+11Hz -0.424762 -0.877443
+ 2.608e+11Hz -0.425435 -0.8771
+ 2.609e+11Hz -0.426108 -0.876757
+ 2.61e+11Hz -0.42678 -0.876413
+ 2.611e+11Hz -0.427452 -0.876069
+ 2.612e+11Hz -0.428124 -0.875724
+ 2.613e+11Hz -0.428794 -0.875378
+ 2.614e+11Hz -0.429465 -0.875032
+ 2.615e+11Hz -0.430135 -0.874686
+ 2.616e+11Hz -0.430805 -0.874338
+ 2.617e+11Hz -0.431474 -0.873991
+ 2.618e+11Hz -0.432143 -0.873642
+ 2.619e+11Hz -0.432811 -0.873293
+ 2.62e+11Hz -0.433479 -0.872944
+ 2.621e+11Hz -0.434146 -0.872594
+ 2.622e+11Hz -0.434813 -0.872244
+ 2.623e+11Hz -0.435479 -0.871893
+ 2.624e+11Hz -0.436145 -0.871541
+ 2.625e+11Hz -0.43681 -0.871189
+ 2.626e+11Hz -0.437475 -0.870837
+ 2.627e+11Hz -0.43814 -0.870484
+ 2.628e+11Hz -0.438803 -0.87013
+ 2.629e+11Hz -0.439467 -0.869776
+ 2.63e+11Hz -0.44013 -0.869422
+ 2.631e+11Hz -0.440792 -0.869067
+ 2.632e+11Hz -0.441454 -0.868711
+ 2.633e+11Hz -0.442115 -0.868355
+ 2.634e+11Hz -0.442776 -0.867999
+ 2.635e+11Hz -0.443437 -0.867642
+ 2.636e+11Hz -0.444096 -0.867284
+ 2.637e+11Hz -0.444756 -0.866926
+ 2.638e+11Hz -0.445415 -0.866568
+ 2.639e+11Hz -0.446073 -0.866209
+ 2.64e+11Hz -0.44673 -0.86585
+ 2.641e+11Hz -0.447388 -0.86549
+ 2.642e+11Hz -0.448044 -0.86513
+ 2.643e+11Hz -0.4487 -0.86477
+ 2.644e+11Hz -0.449356 -0.864409
+ 2.645e+11Hz -0.450011 -0.864048
+ 2.646e+11Hz -0.450666 -0.863686
+ 2.647e+11Hz -0.45132 -0.863324
+ 2.648e+11Hz -0.451973 -0.862961
+ 2.649e+11Hz -0.452626 -0.862598
+ 2.65e+11Hz -0.453278 -0.862235
+ 2.651e+11Hz -0.45393 -0.861871
+ 2.652e+11Hz -0.454581 -0.861507
+ 2.653e+11Hz -0.455232 -0.861143
+ 2.654e+11Hz -0.455882 -0.860778
+ 2.655e+11Hz -0.456532 -0.860413
+ 2.656e+11Hz -0.457181 -0.860048
+ 2.657e+11Hz -0.45783 -0.859682
+ 2.658e+11Hz -0.458478 -0.859316
+ 2.659e+11Hz -0.459125 -0.858949
+ 2.66e+11Hz -0.459772 -0.858583
+ 2.661e+11Hz -0.460419 -0.858216
+ 2.662e+11Hz -0.461065 -0.857848
+ 2.663e+11Hz -0.46171 -0.857481
+ 2.664e+11Hz -0.462355 -0.857113
+ 2.665e+11Hz -0.462999 -0.856745
+ 2.666e+11Hz -0.463643 -0.856377
+ 2.667e+11Hz -0.464286 -0.856008
+ 2.668e+11Hz -0.464929 -0.855639
+ 2.669e+11Hz -0.465571 -0.85527
+ 2.67e+11Hz -0.466213 -0.854901
+ 2.671e+11Hz -0.466854 -0.854531
+ 2.672e+11Hz -0.467495 -0.854161
+ 2.673e+11Hz -0.468135 -0.853791
+ 2.674e+11Hz -0.468775 -0.853421
+ 2.675e+11Hz -0.469414 -0.85305
+ 2.676e+11Hz -0.470053 -0.85268
+ 2.677e+11Hz -0.470691 -0.852309
+ 2.678e+11Hz -0.471329 -0.851938
+ 2.679e+11Hz -0.471966 -0.851567
+ 2.68e+11Hz -0.472603 -0.851196
+ 2.681e+11Hz -0.473239 -0.850824
+ 2.682e+11Hz -0.473875 -0.850452
+ 2.683e+11Hz -0.47451 -0.850081
+ 2.684e+11Hz -0.475145 -0.849709
+ 2.685e+11Hz -0.47578 -0.849337
+ 2.686e+11Hz -0.476414 -0.848964
+ 2.687e+11Hz -0.477048 -0.848592
+ 2.688e+11Hz -0.477681 -0.84822
+ 2.689e+11Hz -0.478314 -0.847847
+ 2.69e+11Hz -0.478946 -0.847475
+ 2.691e+11Hz -0.479578 -0.847102
+ 2.692e+11Hz -0.48021 -0.846729
+ 2.693e+11Hz -0.480841 -0.846356
+ 2.694e+11Hz -0.481472 -0.845983
+ 2.695e+11Hz -0.482102 -0.84561
+ 2.696e+11Hz -0.482732 -0.845237
+ 2.697e+11Hz -0.483362 -0.844864
+ 2.698e+11Hz -0.483992 -0.84449
+ 2.699e+11Hz -0.484621 -0.844117
+ 2.7e+11Hz -0.48525 -0.843743
+ 2.701e+11Hz -0.485878 -0.84337
+ 2.702e+11Hz -0.486506 -0.842996
+ 2.703e+11Hz -0.487134 -0.842623
+ 2.704e+11Hz -0.487761 -0.842249
+ 2.705e+11Hz -0.488389 -0.841875
+ 2.706e+11Hz -0.489016 -0.841502
+ 2.707e+11Hz -0.489642 -0.841128
+ 2.708e+11Hz -0.490269 -0.840754
+ 2.709e+11Hz -0.490895 -0.84038
+ 2.71e+11Hz -0.491521 -0.840006
+ 2.711e+11Hz -0.492147 -0.839633
+ 2.712e+11Hz -0.492772 -0.839259
+ 2.713e+11Hz -0.493398 -0.838885
+ 2.714e+11Hz -0.494023 -0.838511
+ 2.715e+11Hz -0.494648 -0.838137
+ 2.716e+11Hz -0.495272 -0.837763
+ 2.717e+11Hz -0.495897 -0.837388
+ 2.718e+11Hz -0.496522 -0.837014
+ 2.719e+11Hz -0.497146 -0.83664
+ 2.72e+11Hz -0.49777 -0.836266
+ 2.721e+11Hz -0.498394 -0.835892
+ 2.722e+11Hz -0.499018 -0.835517
+ 2.723e+11Hz -0.499642 -0.835143
+ 2.724e+11Hz -0.500265 -0.834769
+ 2.725e+11Hz -0.500889 -0.834394
+ 2.726e+11Hz -0.501513 -0.83402
+ 2.727e+11Hz -0.502136 -0.833646
+ 2.728e+11Hz -0.502759 -0.833271
+ 2.729e+11Hz -0.503383 -0.832897
+ 2.73e+11Hz -0.504006 -0.832522
+ 2.731e+11Hz -0.50463 -0.832147
+ 2.732e+11Hz -0.505253 -0.831772
+ 2.733e+11Hz -0.505876 -0.831398
+ 2.734e+11Hz -0.506499 -0.831023
+ 2.735e+11Hz -0.507123 -0.830648
+ 2.736e+11Hz -0.507746 -0.830273
+ 2.737e+11Hz -0.50837 -0.829898
+ 2.738e+11Hz -0.508993 -0.829522
+ 2.739e+11Hz -0.509616 -0.829147
+ 2.74e+11Hz -0.51024 -0.828772
+ 2.741e+11Hz -0.510864 -0.828396
+ 2.742e+11Hz -0.511487 -0.828021
+ 2.743e+11Hz -0.512111 -0.827645
+ 2.744e+11Hz -0.512735 -0.827269
+ 2.745e+11Hz -0.513359 -0.826893
+ 2.746e+11Hz -0.513983 -0.826517
+ 2.747e+11Hz -0.514607 -0.82614
+ 2.748e+11Hz -0.515232 -0.825764
+ 2.749e+11Hz -0.515856 -0.825387
+ 2.75e+11Hz -0.516481 -0.82501
+ 2.751e+11Hz -0.517106 -0.824633
+ 2.752e+11Hz -0.517731 -0.824256
+ 2.753e+11Hz -0.518356 -0.823879
+ 2.754e+11Hz -0.518981 -0.823501
+ 2.755e+11Hz -0.519607 -0.823123
+ 2.756e+11Hz -0.520232 -0.822745
+ 2.757e+11Hz -0.520858 -0.822367
+ 2.758e+11Hz -0.521484 -0.821988
+ 2.759e+11Hz -0.522111 -0.821609
+ 2.76e+11Hz -0.522737 -0.82123
+ 2.761e+11Hz -0.523364 -0.820851
+ 2.762e+11Hz -0.523991 -0.820471
+ 2.763e+11Hz -0.524618 -0.820091
+ 2.764e+11Hz -0.525246 -0.819711
+ 2.765e+11Hz -0.525873 -0.81933
+ 2.766e+11Hz -0.526501 -0.818949
+ 2.767e+11Hz -0.527129 -0.818568
+ 2.768e+11Hz -0.527758 -0.818186
+ 2.769e+11Hz -0.528386 -0.817804
+ 2.77e+11Hz -0.529015 -0.817422
+ 2.771e+11Hz -0.529645 -0.817039
+ 2.772e+11Hz -0.530274 -0.816655
+ 2.773e+11Hz -0.530904 -0.816272
+ 2.774e+11Hz -0.531534 -0.815888
+ 2.775e+11Hz -0.532164 -0.815503
+ 2.776e+11Hz -0.532795 -0.815118
+ 2.777e+11Hz -0.533426 -0.814733
+ 2.778e+11Hz -0.534057 -0.814347
+ 2.779e+11Hz -0.534688 -0.81396
+ 2.78e+11Hz -0.53532 -0.813573
+ 2.781e+11Hz -0.535952 -0.813186
+ 2.782e+11Hz -0.536584 -0.812798
+ 2.783e+11Hz -0.537217 -0.812409
+ 2.784e+11Hz -0.537849 -0.81202
+ 2.785e+11Hz -0.538482 -0.81163
+ 2.786e+11Hz -0.539116 -0.81124
+ 2.787e+11Hz -0.539749 -0.810849
+ 2.788e+11Hz -0.540383 -0.810457
+ 2.789e+11Hz -0.541017 -0.810065
+ 2.79e+11Hz -0.541652 -0.809673
+ 2.791e+11Hz -0.542287 -0.809279
+ 2.792e+11Hz -0.542921 -0.808885
+ 2.793e+11Hz -0.543557 -0.80849
+ 2.794e+11Hz -0.544192 -0.808095
+ 2.795e+11Hz -0.544828 -0.807699
+ 2.796e+11Hz -0.545464 -0.807302
+ 2.797e+11Hz -0.5461 -0.806904
+ 2.798e+11Hz -0.546736 -0.806506
+ 2.799e+11Hz -0.547373 -0.806107
+ 2.8e+11Hz -0.54801 -0.805707
+ 2.801e+11Hz -0.548647 -0.805307
+ 2.802e+11Hz -0.549284 -0.804905
+ 2.803e+11Hz -0.549921 -0.804503
+ 2.804e+11Hz -0.550559 -0.8041
+ 2.805e+11Hz -0.551197 -0.803697
+ 2.806e+11Hz -0.551835 -0.803292
+ 2.807e+11Hz -0.552473 -0.802887
+ 2.808e+11Hz -0.553111 -0.80248
+ 2.809e+11Hz -0.55375 -0.802073
+ 2.81e+11Hz -0.554389 -0.801665
+ 2.811e+11Hz -0.555027 -0.801256
+ 2.812e+11Hz -0.555666 -0.800847
+ 2.813e+11Hz -0.556305 -0.800436
+ 2.814e+11Hz -0.556945 -0.800024
+ 2.815e+11Hz -0.557584 -0.799612
+ 2.816e+11Hz -0.558223 -0.799198
+ 2.817e+11Hz -0.558863 -0.798784
+ 2.818e+11Hz -0.559502 -0.798369
+ 2.819e+11Hz -0.560142 -0.797953
+ 2.82e+11Hz -0.560781 -0.797535
+ 2.821e+11Hz -0.561421 -0.797117
+ 2.822e+11Hz -0.562061 -0.796698
+ 2.823e+11Hz -0.5627 -0.796278
+ 2.824e+11Hz -0.56334 -0.795857
+ 2.825e+11Hz -0.56398 -0.795435
+ 2.826e+11Hz -0.564619 -0.795012
+ 2.827e+11Hz -0.565259 -0.794588
+ 2.828e+11Hz -0.565899 -0.794162
+ 2.829e+11Hz -0.566538 -0.793736
+ 2.83e+11Hz -0.567178 -0.793309
+ 2.831e+11Hz -0.567817 -0.792881
+ 2.832e+11Hz -0.568456 -0.792452
+ 2.833e+11Hz -0.569096 -0.792021
+ 2.834e+11Hz -0.569735 -0.79159
+ 2.835e+11Hz -0.570374 -0.791158
+ 2.836e+11Hz -0.571012 -0.790724
+ 2.837e+11Hz -0.571651 -0.79029
+ 2.838e+11Hz -0.572289 -0.789854
+ 2.839e+11Hz -0.572928 -0.789418
+ 2.84e+11Hz -0.573566 -0.78898
+ 2.841e+11Hz -0.574204 -0.788541
+ 2.842e+11Hz -0.574841 -0.788102
+ 2.843e+11Hz -0.575479 -0.787661
+ 2.844e+11Hz -0.576116 -0.787219
+ 2.845e+11Hz -0.576753 -0.786776
+ 2.846e+11Hz -0.577389 -0.786332
+ 2.847e+11Hz -0.578026 -0.785887
+ 2.848e+11Hz -0.578662 -0.78544
+ 2.849e+11Hz -0.579297 -0.784993
+ 2.85e+11Hz -0.579933 -0.784545
+ 2.851e+11Hz -0.580568 -0.784095
+ 2.852e+11Hz -0.581202 -0.783645
+ 2.853e+11Hz -0.581836 -0.783193
+ 2.854e+11Hz -0.58247 -0.782741
+ 2.855e+11Hz -0.583104 -0.782287
+ 2.856e+11Hz -0.583737 -0.781833
+ 2.857e+11Hz -0.58437 -0.781377
+ 2.858e+11Hz -0.585002 -0.78092
+ 2.859e+11Hz -0.585633 -0.780462
+ 2.86e+11Hz -0.586265 -0.780003
+ 2.861e+11Hz -0.586896 -0.779544
+ 2.862e+11Hz -0.587526 -0.779083
+ 2.863e+11Hz -0.588156 -0.778621
+ 2.864e+11Hz -0.588785 -0.778158
+ 2.865e+11Hz -0.589414 -0.777694
+ 2.866e+11Hz -0.590042 -0.777229
+ 2.867e+11Hz -0.59067 -0.776763
+ 2.868e+11Hz -0.591297 -0.776296
+ 2.869e+11Hz -0.591923 -0.775828
+ 2.87e+11Hz -0.592549 -0.775359
+ 2.871e+11Hz -0.593175 -0.774889
+ 2.872e+11Hz -0.593799 -0.774418
+ 2.873e+11Hz -0.594423 -0.773946
+ 2.874e+11Hz -0.595047 -0.773473
+ 2.875e+11Hz -0.59567 -0.773
+ 2.876e+11Hz -0.596292 -0.772525
+ 2.877e+11Hz -0.596914 -0.772049
+ 2.878e+11Hz -0.597535 -0.771573
+ 2.879e+11Hz -0.598155 -0.771095
+ 2.88e+11Hz -0.598774 -0.770617
+ 2.881e+11Hz -0.599393 -0.770138
+ 2.882e+11Hz -0.600011 -0.769658
+ 2.883e+11Hz -0.600629 -0.769177
+ 2.884e+11Hz -0.601246 -0.768695
+ 2.885e+11Hz -0.601862 -0.768212
+ 2.886e+11Hz -0.602477 -0.767729
+ 2.887e+11Hz -0.603091 -0.767245
+ 2.888e+11Hz -0.603705 -0.766759
+ 2.889e+11Hz -0.604318 -0.766273
+ 2.89e+11Hz -0.604931 -0.765787
+ 2.891e+11Hz -0.605542 -0.765299
+ 2.892e+11Hz -0.606153 -0.764811
+ 2.893e+11Hz -0.606763 -0.764322
+ 2.894e+11Hz -0.607372 -0.763832
+ 2.895e+11Hz -0.607981 -0.763341
+ 2.896e+11Hz -0.608588 -0.76285
+ 2.897e+11Hz -0.609195 -0.762358
+ 2.898e+11Hz -0.609801 -0.761865
+ 2.899e+11Hz -0.610407 -0.761372
+ 2.9e+11Hz -0.611011 -0.760878
+ 2.901e+11Hz -0.611615 -0.760383
+ 2.902e+11Hz -0.612218 -0.759888
+ 2.903e+11Hz -0.61282 -0.759392
+ 2.904e+11Hz -0.613421 -0.758895
+ 2.905e+11Hz -0.614021 -0.758398
+ 2.906e+11Hz -0.614621 -0.7579
+ 2.907e+11Hz -0.61522 -0.757401
+ 2.908e+11Hz -0.615818 -0.756902
+ 2.909e+11Hz -0.616415 -0.756402
+ 2.91e+11Hz -0.617011 -0.755902
+ 2.911e+11Hz -0.617607 -0.755401
+ 2.912e+11Hz -0.618202 -0.7549
+ 2.913e+11Hz -0.618796 -0.754398
+ 2.914e+11Hz -0.619389 -0.753896
+ 2.915e+11Hz -0.619981 -0.753393
+ 2.916e+11Hz -0.620573 -0.752889
+ 2.917e+11Hz -0.621163 -0.752385
+ 2.918e+11Hz -0.621753 -0.751881
+ 2.919e+11Hz -0.622342 -0.751376
+ 2.92e+11Hz -0.622931 -0.750871
+ 2.921e+11Hz -0.623518 -0.750365
+ 2.922e+11Hz -0.624105 -0.749859
+ 2.923e+11Hz -0.624691 -0.749352
+ 2.924e+11Hz -0.625276 -0.748845
+ 2.925e+11Hz -0.625861 -0.748338
+ 2.926e+11Hz -0.626444 -0.74783
+ 2.927e+11Hz -0.627027 -0.747322
+ 2.928e+11Hz -0.627609 -0.746813
+ 2.929e+11Hz -0.628191 -0.746304
+ 2.93e+11Hz -0.628771 -0.745795
+ 2.931e+11Hz -0.629351 -0.745285
+ 2.932e+11Hz -0.62993 -0.744775
+ 2.933e+11Hz -0.630509 -0.744264
+ 2.934e+11Hz -0.631086 -0.743754
+ 2.935e+11Hz -0.631663 -0.743243
+ 2.936e+11Hz -0.63224 -0.742731
+ 2.937e+11Hz -0.632815 -0.74222
+ 2.938e+11Hz -0.63339 -0.741708
+ 2.939e+11Hz -0.633964 -0.741195
+ 2.94e+11Hz -0.634538 -0.740683
+ 2.941e+11Hz -0.63511 -0.74017
+ 2.942e+11Hz -0.635683 -0.739657
+ 2.943e+11Hz -0.636254 -0.739143
+ 2.944e+11Hz -0.636825 -0.73863
+ 2.945e+11Hz -0.637395 -0.738116
+ 2.946e+11Hz -0.637965 -0.737602
+ 2.947e+11Hz -0.638533 -0.737087
+ 2.948e+11Hz -0.639102 -0.736573
+ 2.949e+11Hz -0.639669 -0.736058
+ 2.95e+11Hz -0.640237 -0.735543
+ 2.951e+11Hz -0.640803 -0.735027
+ 2.952e+11Hz -0.641369 -0.734512
+ 2.953e+11Hz -0.641934 -0.733996
+ 2.954e+11Hz -0.642499 -0.73348
+ 2.955e+11Hz -0.643063 -0.732963
+ 2.956e+11Hz -0.643627 -0.732447
+ 2.957e+11Hz -0.64419 -0.73193
+ 2.958e+11Hz -0.644752 -0.731413
+ 2.959e+11Hz -0.645314 -0.730896
+ 2.96e+11Hz -0.645876 -0.730378
+ 2.961e+11Hz -0.646437 -0.729861
+ 2.962e+11Hz -0.646997 -0.729343
+ 2.963e+11Hz -0.647557 -0.728825
+ 2.964e+11Hz -0.648117 -0.728307
+ 2.965e+11Hz -0.648676 -0.727788
+ 2.966e+11Hz -0.649235 -0.727269
+ 2.967e+11Hz -0.649793 -0.72675
+ 2.968e+11Hz -0.65035 -0.726231
+ 2.969e+11Hz -0.650908 -0.725712
+ 2.97e+11Hz -0.651464 -0.725192
+ 2.971e+11Hz -0.652021 -0.724672
+ 2.972e+11Hz -0.652577 -0.724152
+ 2.973e+11Hz -0.653132 -0.723631
+ 2.974e+11Hz -0.653687 -0.723111
+ 2.975e+11Hz -0.654242 -0.72259
+ 2.976e+11Hz -0.654797 -0.722069
+ 2.977e+11Hz -0.655351 -0.721547
+ 2.978e+11Hz -0.655904 -0.721026
+ 2.979e+11Hz -0.656457 -0.720504
+ 2.98e+11Hz -0.65701 -0.719981
+ 2.981e+11Hz -0.657563 -0.719459
+ 2.982e+11Hz -0.658115 -0.718936
+ 2.983e+11Hz -0.658667 -0.718413
+ 2.984e+11Hz -0.659218 -0.71789
+ 2.985e+11Hz -0.659769 -0.717366
+ 2.986e+11Hz -0.66032 -0.716842
+ 2.987e+11Hz -0.66087 -0.716318
+ 2.988e+11Hz -0.66142 -0.715793
+ 2.989e+11Hz -0.66197 -0.715268
+ 2.99e+11Hz -0.66252 -0.714743
+ 2.991e+11Hz -0.663069 -0.714218
+ 2.992e+11Hz -0.663618 -0.713692
+ 2.993e+11Hz -0.664166 -0.713165
+ 2.994e+11Hz -0.664715 -0.712639
+ 2.995e+11Hz -0.665262 -0.712112
+ 2.996e+11Hz -0.66581 -0.711584
+ 2.997e+11Hz -0.666357 -0.711057
+ 2.998e+11Hz -0.666905 -0.710528
+ 2.999e+11Hz -0.667451 -0.71
+ 3e+11Hz -0.667998 -0.709471
+ ]

A21 %vd(10 3) %vd(21, 22) xfer3
.model xfer3 xfer R_I=true table=[
+ 0Hz 0.995382 0
+ 1e+08Hz 0.995382 -0.000812217
+ 2e+08Hz 0.99538 -0.00162442
+ 3e+08Hz 0.995377 -0.0024366
+ 4e+08Hz 0.995372 -0.00324873
+ 5e+08Hz 0.995367 -0.00406082
+ 6e+08Hz 0.99536 -0.00487284
+ 7e+08Hz 0.995352 -0.00568478
+ 8e+08Hz 0.995343 -0.00649662
+ 9e+08Hz 0.995333 -0.00730836
+ 1e+09Hz 0.995321 -0.00811999
+ 1.1e+09Hz 0.995308 -0.00893148
+ 1.2e+09Hz 0.995294 -0.00974282
+ 1.3e+09Hz 0.995279 -0.010554
+ 1.4e+09Hz 0.995263 -0.011365
+ 1.5e+09Hz 0.995245 -0.0121759
+ 1.6e+09Hz 0.995226 -0.0129865
+ 1.7e+09Hz 0.995206 -0.013797
+ 1.8e+09Hz 0.995185 -0.0146072
+ 1.9e+09Hz 0.995163 -0.0154172
+ 2e+09Hz 0.995139 -0.0162269
+ 2.1e+09Hz 0.995115 -0.0170364
+ 2.2e+09Hz 0.995089 -0.0178456
+ 2.3e+09Hz 0.995062 -0.0186546
+ 2.4e+09Hz 0.995034 -0.0194632
+ 2.5e+09Hz 0.995005 -0.0202716
+ 2.6e+09Hz 0.994974 -0.0210796
+ 2.7e+09Hz 0.994943 -0.0218873
+ 2.8e+09Hz 0.99491 -0.0226947
+ 2.9e+09Hz 0.994876 -0.0235018
+ 3e+09Hz 0.994841 -0.0243085
+ 3.1e+09Hz 0.994806 -0.0251148
+ 3.2e+09Hz 0.994768 -0.0259208
+ 3.3e+09Hz 0.99473 -0.0267263
+ 3.4e+09Hz 0.994691 -0.0275315
+ 3.5e+09Hz 0.994651 -0.0283363
+ 3.6e+09Hz 0.99461 -0.0291407
+ 3.7e+09Hz 0.994567 -0.0299446
+ 3.8e+09Hz 0.994524 -0.0307482
+ 3.9e+09Hz 0.99448 -0.0315512
+ 4e+09Hz 0.994434 -0.0323539
+ 4.1e+09Hz 0.994388 -0.0331561
+ 4.2e+09Hz 0.99434 -0.0339578
+ 4.3e+09Hz 0.994292 -0.0347591
+ 4.4e+09Hz 0.994243 -0.0355599
+ 4.5e+09Hz 0.994192 -0.0363602
+ 4.6e+09Hz 0.994141 -0.0371601
+ 4.7e+09Hz 0.994089 -0.0379594
+ 4.8e+09Hz 0.994036 -0.0387583
+ 4.9e+09Hz 0.993982 -0.0395566
+ 5e+09Hz 0.993927 -0.0403545
+ 5.1e+09Hz 0.993871 -0.0411518
+ 5.2e+09Hz 0.993814 -0.0419486
+ 5.3e+09Hz 0.993757 -0.0427449
+ 5.4e+09Hz 0.993698 -0.0435407
+ 5.5e+09Hz 0.993639 -0.0443359
+ 5.6e+09Hz 0.993579 -0.0451306
+ 5.7e+09Hz 0.993518 -0.0459248
+ 5.8e+09Hz 0.993456 -0.0467184
+ 5.9e+09Hz 0.993394 -0.0475115
+ 6e+09Hz 0.99333 -0.048304
+ 6.1e+09Hz 0.993266 -0.049096
+ 6.2e+09Hz 0.993201 -0.0498875
+ 6.3e+09Hz 0.993135 -0.0506783
+ 6.4e+09Hz 0.993069 -0.0514687
+ 6.5e+09Hz 0.993002 -0.0522585
+ 6.6e+09Hz 0.992934 -0.0530477
+ 6.7e+09Hz 0.992865 -0.0538364
+ 6.8e+09Hz 0.992796 -0.0546245
+ 6.9e+09Hz 0.992726 -0.0554121
+ 7e+09Hz 0.992655 -0.0561991
+ 7.1e+09Hz 0.992584 -0.0569855
+ 7.2e+09Hz 0.992512 -0.0577714
+ 7.3e+09Hz 0.992439 -0.0585568
+ 7.4e+09Hz 0.992366 -0.0593416
+ 7.5e+09Hz 0.992292 -0.0601258
+ 7.6e+09Hz 0.992217 -0.0609095
+ 7.7e+09Hz 0.992142 -0.0616927
+ 7.8e+09Hz 0.992066 -0.0624753
+ 7.9e+09Hz 0.99199 -0.0632574
+ 8e+09Hz 0.991913 -0.0640389
+ 8.1e+09Hz 0.991836 -0.0648199
+ 8.2e+09Hz 0.991758 -0.0656004
+ 8.3e+09Hz 0.991679 -0.0663804
+ 8.4e+09Hz 0.9916 -0.0671598
+ 8.5e+09Hz 0.991521 -0.0679387
+ 8.6e+09Hz 0.99144 -0.0687171
+ 8.7e+09Hz 0.99136 -0.0694949
+ 8.8e+09Hz 0.991279 -0.0702723
+ 8.9e+09Hz 0.991197 -0.0710492
+ 9e+09Hz 0.991115 -0.0718255
+ 9.1e+09Hz 0.991033 -0.0726014
+ 9.2e+09Hz 0.99095 -0.0733768
+ 9.3e+09Hz 0.990866 -0.0741517
+ 9.4e+09Hz 0.990782 -0.0749261
+ 9.5e+09Hz 0.990698 -0.0757001
+ 9.6e+09Hz 0.990613 -0.0764736
+ 9.7e+09Hz 0.990528 -0.0772466
+ 9.8e+09Hz 0.990443 -0.0780192
+ 9.9e+09Hz 0.990357 -0.0787913
+ 1e+10Hz 0.99027 -0.079563
+ 1.01e+10Hz 0.990184 -0.0803343
+ 1.02e+10Hz 0.990097 -0.0811051
+ 1.03e+10Hz 0.990009 -0.0818755
+ 1.04e+10Hz 0.989921 -0.0826455
+ 1.05e+10Hz 0.989833 -0.0834151
+ 1.06e+10Hz 0.989744 -0.0841844
+ 1.07e+10Hz 0.989655 -0.0849532
+ 1.08e+10Hz 0.989566 -0.0857216
+ 1.09e+10Hz 0.989477 -0.0864897
+ 1.1e+10Hz 0.989387 -0.0872574
+ 1.11e+10Hz 0.989296 -0.0880247
+ 1.12e+10Hz 0.989206 -0.0887917
+ 1.13e+10Hz 0.989115 -0.0895584
+ 1.14e+10Hz 0.989023 -0.0903247
+ 1.15e+10Hz 0.988932 -0.0910906
+ 1.16e+10Hz 0.98884 -0.0918563
+ 1.17e+10Hz 0.988748 -0.0926217
+ 1.18e+10Hz 0.988655 -0.0933867
+ 1.19e+10Hz 0.988563 -0.0941515
+ 1.2e+10Hz 0.988469 -0.0949159
+ 1.21e+10Hz 0.988376 -0.0956801
+ 1.22e+10Hz 0.988282 -0.096444
+ 1.23e+10Hz 0.988188 -0.0972077
+ 1.24e+10Hz 0.988094 -0.0979711
+ 1.25e+10Hz 0.988 -0.0987343
+ 1.26e+10Hz 0.987905 -0.0994972
+ 1.27e+10Hz 0.98781 -0.10026
+ 1.28e+10Hz 0.987714 -0.101022
+ 1.29e+10Hz 0.987618 -0.101785
+ 1.3e+10Hz 0.987523 -0.102547
+ 1.31e+10Hz 0.987426 -0.103309
+ 1.32e+10Hz 0.98733 -0.10407
+ 1.33e+10Hz 0.987233 -0.104832
+ 1.34e+10Hz 0.987136 -0.105593
+ 1.35e+10Hz 0.987038 -0.106354
+ 1.36e+10Hz 0.986941 -0.107115
+ 1.37e+10Hz 0.986843 -0.107876
+ 1.38e+10Hz 0.986744 -0.108637
+ 1.39e+10Hz 0.986646 -0.109397
+ 1.4e+10Hz 0.986547 -0.110158
+ 1.41e+10Hz 0.986448 -0.110918
+ 1.42e+10Hz 0.986348 -0.111678
+ 1.43e+10Hz 0.986249 -0.112438
+ 1.44e+10Hz 0.986149 -0.113198
+ 1.45e+10Hz 0.986048 -0.113958
+ 1.46e+10Hz 0.985948 -0.114718
+ 1.47e+10Hz 0.985847 -0.115478
+ 1.48e+10Hz 0.985745 -0.116237
+ 1.49e+10Hz 0.985644 -0.116997
+ 1.5e+10Hz 0.985542 -0.117756
+ 1.51e+10Hz 0.98544 -0.118516
+ 1.52e+10Hz 0.985337 -0.119275
+ 1.53e+10Hz 0.985234 -0.120035
+ 1.54e+10Hz 0.985131 -0.120794
+ 1.55e+10Hz 0.985028 -0.121554
+ 1.56e+10Hz 0.984924 -0.122313
+ 1.57e+10Hz 0.98482 -0.123072
+ 1.58e+10Hz 0.984715 -0.123831
+ 1.59e+10Hz 0.98461 -0.124591
+ 1.6e+10Hz 0.984505 -0.12535
+ 1.61e+10Hz 0.984399 -0.126109
+ 1.62e+10Hz 0.984293 -0.126869
+ 1.63e+10Hz 0.984187 -0.127628
+ 1.64e+10Hz 0.98408 -0.128387
+ 1.65e+10Hz 0.983973 -0.129147
+ 1.66e+10Hz 0.983865 -0.129906
+ 1.67e+10Hz 0.983758 -0.130665
+ 1.68e+10Hz 0.983649 -0.131425
+ 1.69e+10Hz 0.983541 -0.132184
+ 1.7e+10Hz 0.983431 -0.132944
+ 1.71e+10Hz 0.983322 -0.133703
+ 1.72e+10Hz 0.983212 -0.134463
+ 1.73e+10Hz 0.983102 -0.135222
+ 1.74e+10Hz 0.982991 -0.135982
+ 1.75e+10Hz 0.98288 -0.136742
+ 1.76e+10Hz 0.982768 -0.137502
+ 1.77e+10Hz 0.982656 -0.138262
+ 1.78e+10Hz 0.982543 -0.139021
+ 1.79e+10Hz 0.98243 -0.139781
+ 1.8e+10Hz 0.982317 -0.140541
+ 1.81e+10Hz 0.982203 -0.141302
+ 1.82e+10Hz 0.982088 -0.142062
+ 1.83e+10Hz 0.981973 -0.142822
+ 1.84e+10Hz 0.981858 -0.143582
+ 1.85e+10Hz 0.981742 -0.144343
+ 1.86e+10Hz 0.981625 -0.145103
+ 1.87e+10Hz 0.981508 -0.145863
+ 1.88e+10Hz 0.981391 -0.146624
+ 1.89e+10Hz 0.981273 -0.147385
+ 1.9e+10Hz 0.981154 -0.148145
+ 1.91e+10Hz 0.981035 -0.148906
+ 1.92e+10Hz 0.980916 -0.149667
+ 1.93e+10Hz 0.980796 -0.150428
+ 1.94e+10Hz 0.980675 -0.151189
+ 1.95e+10Hz 0.980554 -0.15195
+ 1.96e+10Hz 0.980432 -0.152711
+ 1.97e+10Hz 0.980309 -0.153472
+ 1.98e+10Hz 0.980186 -0.154233
+ 1.99e+10Hz 0.980063 -0.154995
+ 2e+10Hz 0.979939 -0.155756
+ 2.01e+10Hz 0.979814 -0.156517
+ 2.02e+10Hz 0.979689 -0.157279
+ 2.03e+10Hz 0.979563 -0.15804
+ 2.04e+10Hz 0.979436 -0.158802
+ 2.05e+10Hz 0.979309 -0.159563
+ 2.06e+10Hz 0.979182 -0.160325
+ 2.07e+10Hz 0.979053 -0.161087
+ 2.08e+10Hz 0.978924 -0.161848
+ 2.09e+10Hz 0.978795 -0.16261
+ 2.1e+10Hz 0.978665 -0.163372
+ 2.11e+10Hz 0.978534 -0.164134
+ 2.12e+10Hz 0.978402 -0.164896
+ 2.13e+10Hz 0.97827 -0.165657
+ 2.14e+10Hz 0.978137 -0.166419
+ 2.15e+10Hz 0.978004 -0.167181
+ 2.16e+10Hz 0.97787 -0.167943
+ 2.17e+10Hz 0.977735 -0.168705
+ 2.18e+10Hz 0.977599 -0.169467
+ 2.19e+10Hz 0.977463 -0.170229
+ 2.2e+10Hz 0.977327 -0.170991
+ 2.21e+10Hz 0.977189 -0.171753
+ 2.22e+10Hz 0.977051 -0.172515
+ 2.23e+10Hz 0.976912 -0.173276
+ 2.24e+10Hz 0.976773 -0.174038
+ 2.25e+10Hz 0.976633 -0.1748
+ 2.26e+10Hz 0.976492 -0.175562
+ 2.27e+10Hz 0.97635 -0.176324
+ 2.28e+10Hz 0.976208 -0.177085
+ 2.29e+10Hz 0.976065 -0.177847
+ 2.3e+10Hz 0.975921 -0.178609
+ 2.31e+10Hz 0.975777 -0.17937
+ 2.32e+10Hz 0.975632 -0.180132
+ 2.33e+10Hz 0.975486 -0.180893
+ 2.34e+10Hz 0.97534 -0.181655
+ 2.35e+10Hz 0.975192 -0.182416
+ 2.36e+10Hz 0.975045 -0.183177
+ 2.37e+10Hz 0.974896 -0.183938
+ 2.38e+10Hz 0.974747 -0.184699
+ 2.39e+10Hz 0.974597 -0.18546
+ 2.4e+10Hz 0.974446 -0.186221
+ 2.41e+10Hz 0.974294 -0.186982
+ 2.42e+10Hz 0.974142 -0.187743
+ 2.43e+10Hz 0.973989 -0.188503
+ 2.44e+10Hz 0.973836 -0.189263
+ 2.45e+10Hz 0.973682 -0.190024
+ 2.46e+10Hz 0.973527 -0.190784
+ 2.47e+10Hz 0.973371 -0.191544
+ 2.48e+10Hz 0.973214 -0.192304
+ 2.49e+10Hz 0.973057 -0.193064
+ 2.5e+10Hz 0.9729 -0.193823
+ 2.51e+10Hz 0.972741 -0.194583
+ 2.52e+10Hz 0.972582 -0.195342
+ 2.53e+10Hz 0.972422 -0.196101
+ 2.54e+10Hz 0.972261 -0.19686
+ 2.55e+10Hz 0.9721 -0.197619
+ 2.56e+10Hz 0.971938 -0.198378
+ 2.57e+10Hz 0.971775 -0.199136
+ 2.58e+10Hz 0.971611 -0.199894
+ 2.59e+10Hz 0.971447 -0.200652
+ 2.6e+10Hz 0.971282 -0.20141
+ 2.61e+10Hz 0.971117 -0.202168
+ 2.62e+10Hz 0.970951 -0.202925
+ 2.63e+10Hz 0.970784 -0.203683
+ 2.64e+10Hz 0.970616 -0.20444
+ 2.65e+10Hz 0.970448 -0.205197
+ 2.66e+10Hz 0.970279 -0.205953
+ 2.67e+10Hz 0.970109 -0.20671
+ 2.68e+10Hz 0.969939 -0.207466
+ 2.69e+10Hz 0.969768 -0.208222
+ 2.7e+10Hz 0.969596 -0.208978
+ 2.71e+10Hz 0.969424 -0.209733
+ 2.72e+10Hz 0.969251 -0.210489
+ 2.73e+10Hz 0.969077 -0.211244
+ 2.74e+10Hz 0.968903 -0.211998
+ 2.75e+10Hz 0.968728 -0.212753
+ 2.76e+10Hz 0.968552 -0.213507
+ 2.77e+10Hz 0.968376 -0.214261
+ 2.78e+10Hz 0.968199 -0.215015
+ 2.79e+10Hz 0.968021 -0.215769
+ 2.8e+10Hz 0.967843 -0.216522
+ 2.81e+10Hz 0.967664 -0.217275
+ 2.82e+10Hz 0.967485 -0.218028
+ 2.83e+10Hz 0.967304 -0.21878
+ 2.84e+10Hz 0.967124 -0.219533
+ 2.85e+10Hz 0.966942 -0.220285
+ 2.86e+10Hz 0.96676 -0.221036
+ 2.87e+10Hz 0.966578 -0.221788
+ 2.88e+10Hz 0.966395 -0.222539
+ 2.89e+10Hz 0.966211 -0.22329
+ 2.9e+10Hz 0.966026 -0.22404
+ 2.91e+10Hz 0.965842 -0.224791
+ 2.92e+10Hz 0.965656 -0.225541
+ 2.93e+10Hz 0.96547 -0.226291
+ 2.94e+10Hz 0.965283 -0.22704
+ 2.95e+10Hz 0.965096 -0.227789
+ 2.96e+10Hz 0.964908 -0.228538
+ 2.97e+10Hz 0.964719 -0.229287
+ 2.98e+10Hz 0.96453 -0.230035
+ 2.99e+10Hz 0.964341 -0.230784
+ 3e+10Hz 0.96415 -0.231531
+ 3.01e+10Hz 0.96396 -0.232279
+ 3.02e+10Hz 0.963768 -0.233026
+ 3.03e+10Hz 0.963577 -0.233773
+ 3.04e+10Hz 0.963384 -0.23452
+ 3.05e+10Hz 0.963191 -0.235266
+ 3.06e+10Hz 0.962998 -0.236013
+ 3.07e+10Hz 0.962804 -0.236758
+ 3.08e+10Hz 0.962609 -0.237504
+ 3.09e+10Hz 0.962414 -0.238249
+ 3.1e+10Hz 0.962219 -0.238994
+ 3.11e+10Hz 0.962023 -0.239739
+ 3.12e+10Hz 0.961826 -0.240484
+ 3.13e+10Hz 0.961629 -0.241228
+ 3.14e+10Hz 0.961431 -0.241972
+ 3.15e+10Hz 0.961233 -0.242716
+ 3.16e+10Hz 0.961034 -0.243459
+ 3.17e+10Hz 0.960835 -0.244202
+ 3.18e+10Hz 0.960636 -0.244945
+ 3.19e+10Hz 0.960435 -0.245688
+ 3.2e+10Hz 0.960235 -0.24643
+ 3.21e+10Hz 0.960034 -0.247172
+ 3.22e+10Hz 0.959832 -0.247914
+ 3.23e+10Hz 0.95963 -0.248656
+ 3.24e+10Hz 0.959427 -0.249397
+ 3.25e+10Hz 0.959224 -0.250138
+ 3.26e+10Hz 0.959021 -0.250879
+ 3.27e+10Hz 0.958817 -0.25162
+ 3.28e+10Hz 0.958612 -0.25236
+ 3.29e+10Hz 0.958407 -0.2531
+ 3.3e+10Hz 0.958202 -0.25384
+ 3.31e+10Hz 0.957996 -0.25458
+ 3.32e+10Hz 0.957789 -0.255319
+ 3.33e+10Hz 0.957583 -0.256058
+ 3.34e+10Hz 0.957375 -0.256797
+ 3.35e+10Hz 0.957168 -0.257536
+ 3.36e+10Hz 0.956959 -0.258275
+ 3.37e+10Hz 0.956751 -0.259013
+ 3.38e+10Hz 0.956542 -0.259751
+ 3.39e+10Hz 0.956332 -0.260489
+ 3.4e+10Hz 0.956122 -0.261227
+ 3.41e+10Hz 0.955911 -0.261964
+ 3.42e+10Hz 0.955701 -0.262701
+ 3.43e+10Hz 0.955489 -0.263438
+ 3.44e+10Hz 0.955277 -0.264175
+ 3.45e+10Hz 0.955065 -0.264912
+ 3.46e+10Hz 0.954852 -0.265649
+ 3.47e+10Hz 0.954639 -0.266385
+ 3.48e+10Hz 0.954426 -0.267121
+ 3.49e+10Hz 0.954212 -0.267857
+ 3.5e+10Hz 0.953997 -0.268593
+ 3.51e+10Hz 0.953782 -0.269328
+ 3.52e+10Hz 0.953567 -0.270064
+ 3.53e+10Hz 0.953351 -0.270799
+ 3.54e+10Hz 0.953134 -0.271534
+ 3.55e+10Hz 0.952918 -0.272269
+ 3.56e+10Hz 0.952701 -0.273003
+ 3.57e+10Hz 0.952483 -0.273738
+ 3.58e+10Hz 0.952265 -0.274472
+ 3.59e+10Hz 0.952046 -0.275207
+ 3.6e+10Hz 0.951827 -0.275941
+ 3.61e+10Hz 0.951608 -0.276675
+ 3.62e+10Hz 0.951388 -0.277409
+ 3.63e+10Hz 0.951168 -0.278142
+ 3.64e+10Hz 0.950947 -0.278876
+ 3.65e+10Hz 0.950725 -0.279609
+ 3.66e+10Hz 0.950504 -0.280342
+ 3.67e+10Hz 0.950282 -0.281075
+ 3.68e+10Hz 0.950059 -0.281808
+ 3.69e+10Hz 0.949836 -0.282541
+ 3.7e+10Hz 0.949612 -0.283274
+ 3.71e+10Hz 0.949388 -0.284007
+ 3.72e+10Hz 0.949164 -0.284739
+ 3.73e+10Hz 0.948939 -0.285471
+ 3.74e+10Hz 0.948713 -0.286204
+ 3.75e+10Hz 0.948487 -0.286936
+ 3.76e+10Hz 0.948261 -0.287668
+ 3.77e+10Hz 0.948034 -0.2884
+ 3.78e+10Hz 0.947807 -0.289132
+ 3.79e+10Hz 0.947579 -0.289863
+ 3.8e+10Hz 0.947351 -0.290595
+ 3.81e+10Hz 0.947122 -0.291326
+ 3.82e+10Hz 0.946893 -0.292058
+ 3.83e+10Hz 0.946663 -0.292789
+ 3.84e+10Hz 0.946433 -0.29352
+ 3.85e+10Hz 0.946202 -0.294251
+ 3.86e+10Hz 0.945971 -0.294982
+ 3.87e+10Hz 0.945739 -0.295713
+ 3.88e+10Hz 0.945507 -0.296444
+ 3.89e+10Hz 0.945274 -0.297175
+ 3.9e+10Hz 0.945041 -0.297905
+ 3.91e+10Hz 0.944807 -0.298636
+ 3.92e+10Hz 0.944573 -0.299366
+ 3.93e+10Hz 0.944338 -0.300097
+ 3.94e+10Hz 0.944103 -0.300827
+ 3.95e+10Hz 0.943867 -0.301557
+ 3.96e+10Hz 0.94363 -0.302287
+ 3.97e+10Hz 0.943394 -0.303017
+ 3.98e+10Hz 0.943156 -0.303747
+ 3.99e+10Hz 0.942918 -0.304477
+ 4e+10Hz 0.94268 -0.305206
+ 4.01e+10Hz 0.942441 -0.305936
+ 4.02e+10Hz 0.942201 -0.306666
+ 4.03e+10Hz 0.941961 -0.307395
+ 4.04e+10Hz 0.94172 -0.308124
+ 4.05e+10Hz 0.941479 -0.308854
+ 4.06e+10Hz 0.941237 -0.309583
+ 4.07e+10Hz 0.940995 -0.310312
+ 4.08e+10Hz 0.940752 -0.311041
+ 4.09e+10Hz 0.940509 -0.31177
+ 4.1e+10Hz 0.940265 -0.312499
+ 4.11e+10Hz 0.94002 -0.313227
+ 4.12e+10Hz 0.939775 -0.313956
+ 4.13e+10Hz 0.939529 -0.314685
+ 4.14e+10Hz 0.939283 -0.315413
+ 4.15e+10Hz 0.939036 -0.316141
+ 4.16e+10Hz 0.938789 -0.31687
+ 4.17e+10Hz 0.938541 -0.317598
+ 4.18e+10Hz 0.938292 -0.318326
+ 4.19e+10Hz 0.938043 -0.319054
+ 4.2e+10Hz 0.937793 -0.319782
+ 4.21e+10Hz 0.937543 -0.320509
+ 4.22e+10Hz 0.937292 -0.321237
+ 4.23e+10Hz 0.93704 -0.321965
+ 4.24e+10Hz 0.936788 -0.322692
+ 4.25e+10Hz 0.936535 -0.323419
+ 4.26e+10Hz 0.936282 -0.324146
+ 4.27e+10Hz 0.936028 -0.324874
+ 4.28e+10Hz 0.935773 -0.3256
+ 4.29e+10Hz 0.935518 -0.326327
+ 4.3e+10Hz 0.935262 -0.327054
+ 4.31e+10Hz 0.935006 -0.327781
+ 4.32e+10Hz 0.934749 -0.328507
+ 4.33e+10Hz 0.934491 -0.329233
+ 4.34e+10Hz 0.934233 -0.32996
+ 4.35e+10Hz 0.933974 -0.330686
+ 4.36e+10Hz 0.933714 -0.331412
+ 4.37e+10Hz 0.933454 -0.332137
+ 4.38e+10Hz 0.933193 -0.332863
+ 4.39e+10Hz 0.932932 -0.333589
+ 4.4e+10Hz 0.932669 -0.334314
+ 4.41e+10Hz 0.932407 -0.335039
+ 4.42e+10Hz 0.932143 -0.335764
+ 4.43e+10Hz 0.931879 -0.336489
+ 4.44e+10Hz 0.931615 -0.337214
+ 4.45e+10Hz 0.93135 -0.337938
+ 4.46e+10Hz 0.931084 -0.338663
+ 4.47e+10Hz 0.930817 -0.339387
+ 4.48e+10Hz 0.93055 -0.340111
+ 4.49e+10Hz 0.930282 -0.340835
+ 4.5e+10Hz 0.930014 -0.341559
+ 4.51e+10Hz 0.929744 -0.342282
+ 4.52e+10Hz 0.929475 -0.343006
+ 4.53e+10Hz 0.929204 -0.343729
+ 4.54e+10Hz 0.928933 -0.344452
+ 4.55e+10Hz 0.928662 -0.345175
+ 4.56e+10Hz 0.928389 -0.345897
+ 4.57e+10Hz 0.928116 -0.34662
+ 4.58e+10Hz 0.927843 -0.347342
+ 4.59e+10Hz 0.927568 -0.348064
+ 4.6e+10Hz 0.927293 -0.348786
+ 4.61e+10Hz 0.927018 -0.349507
+ 4.62e+10Hz 0.926742 -0.350229
+ 4.63e+10Hz 0.926465 -0.35095
+ 4.64e+10Hz 0.926187 -0.351671
+ 4.65e+10Hz 0.925909 -0.352391
+ 4.66e+10Hz 0.92563 -0.353112
+ 4.67e+10Hz 0.925351 -0.353832
+ 4.68e+10Hz 0.925071 -0.354552
+ 4.69e+10Hz 0.92479 -0.355272
+ 4.7e+10Hz 0.924509 -0.355992
+ 4.71e+10Hz 0.924227 -0.356711
+ 4.72e+10Hz 0.923944 -0.35743
+ 4.73e+10Hz 0.923661 -0.358149
+ 4.74e+10Hz 0.923377 -0.358867
+ 4.75e+10Hz 0.923092 -0.359586
+ 4.76e+10Hz 0.922807 -0.360304
+ 4.77e+10Hz 0.922521 -0.361022
+ 4.78e+10Hz 0.922235 -0.361739
+ 4.79e+10Hz 0.921948 -0.362457
+ 4.8e+10Hz 0.92166 -0.363174
+ 4.81e+10Hz 0.921371 -0.36389
+ 4.82e+10Hz 0.921082 -0.364607
+ 4.83e+10Hz 0.920793 -0.365323
+ 4.84e+10Hz 0.920503 -0.366039
+ 4.85e+10Hz 0.920212 -0.366755
+ 4.86e+10Hz 0.91992 -0.36747
+ 4.87e+10Hz 0.919628 -0.368185
+ 4.88e+10Hz 0.919335 -0.3689
+ 4.89e+10Hz 0.919042 -0.369615
+ 4.9e+10Hz 0.918748 -0.370329
+ 4.91e+10Hz 0.918454 -0.371043
+ 4.92e+10Hz 0.918158 -0.371756
+ 4.93e+10Hz 0.917863 -0.37247
+ 4.94e+10Hz 0.917566 -0.373183
+ 4.95e+10Hz 0.917269 -0.373896
+ 4.96e+10Hz 0.916972 -0.374608
+ 4.97e+10Hz 0.916673 -0.37532
+ 4.98e+10Hz 0.916375 -0.376032
+ 4.99e+10Hz 0.916075 -0.376744
+ 5e+10Hz 0.915775 -0.377455
+ 5.01e+10Hz 0.915475 -0.378166
+ 5.02e+10Hz 0.915174 -0.378877
+ 5.03e+10Hz 0.914872 -0.379587
+ 5.04e+10Hz 0.914569 -0.380297
+ 5.05e+10Hz 0.914267 -0.381007
+ 5.06e+10Hz 0.913963 -0.381716
+ 5.07e+10Hz 0.913659 -0.382425
+ 5.08e+10Hz 0.913354 -0.383134
+ 5.09e+10Hz 0.913049 -0.383842
+ 5.1e+10Hz 0.912743 -0.38455
+ 5.11e+10Hz 0.912437 -0.385258
+ 5.12e+10Hz 0.91213 -0.385966
+ 5.13e+10Hz 0.911823 -0.386673
+ 5.14e+10Hz 0.911515 -0.38738
+ 5.15e+10Hz 0.911206 -0.388086
+ 5.16e+10Hz 0.910897 -0.388792
+ 5.17e+10Hz 0.910587 -0.389498
+ 5.18e+10Hz 0.910277 -0.390204
+ 5.19e+10Hz 0.909967 -0.390909
+ 5.2e+10Hz 0.909655 -0.391614
+ 5.21e+10Hz 0.909343 -0.392318
+ 5.22e+10Hz 0.909031 -0.393023
+ 5.23e+10Hz 0.908718 -0.393726
+ 5.24e+10Hz 0.908405 -0.39443
+ 5.25e+10Hz 0.908091 -0.395133
+ 5.26e+10Hz 0.907776 -0.395836
+ 5.27e+10Hz 0.907461 -0.396539
+ 5.28e+10Hz 0.907146 -0.397241
+ 5.29e+10Hz 0.90683 -0.397943
+ 5.3e+10Hz 0.906513 -0.398645
+ 5.31e+10Hz 0.906196 -0.399346
+ 5.32e+10Hz 0.905878 -0.400047
+ 5.33e+10Hz 0.90556 -0.400748
+ 5.34e+10Hz 0.905242 -0.401448
+ 5.35e+10Hz 0.904922 -0.402148
+ 5.36e+10Hz 0.904603 -0.402848
+ 5.37e+10Hz 0.904283 -0.403547
+ 5.38e+10Hz 0.903962 -0.404246
+ 5.39e+10Hz 0.903641 -0.404945
+ 5.4e+10Hz 0.903319 -0.405643
+ 5.41e+10Hz 0.902997 -0.406341
+ 5.42e+10Hz 0.902675 -0.407039
+ 5.43e+10Hz 0.902351 -0.407737
+ 5.44e+10Hz 0.902028 -0.408434
+ 5.45e+10Hz 0.901704 -0.409131
+ 5.46e+10Hz 0.901379 -0.409827
+ 5.47e+10Hz 0.901054 -0.410523
+ 5.48e+10Hz 0.900729 -0.411219
+ 5.49e+10Hz 0.900403 -0.411915
+ 5.5e+10Hz 0.900076 -0.41261
+ 5.51e+10Hz 0.899749 -0.413305
+ 5.52e+10Hz 0.899422 -0.414
+ 5.53e+10Hz 0.899094 -0.414694
+ 5.54e+10Hz 0.898765 -0.415388
+ 5.55e+10Hz 0.898437 -0.416082
+ 5.56e+10Hz 0.898107 -0.416776
+ 5.57e+10Hz 0.897778 -0.417469
+ 5.58e+10Hz 0.897447 -0.418162
+ 5.59e+10Hz 0.897117 -0.418854
+ 5.6e+10Hz 0.896785 -0.419547
+ 5.61e+10Hz 0.896454 -0.420239
+ 5.62e+10Hz 0.896122 -0.420931
+ 5.63e+10Hz 0.895789 -0.421622
+ 5.64e+10Hz 0.895456 -0.422313
+ 5.65e+10Hz 0.895122 -0.423004
+ 5.66e+10Hz 0.894788 -0.423695
+ 5.67e+10Hz 0.894454 -0.424385
+ 5.68e+10Hz 0.894119 -0.425075
+ 5.69e+10Hz 0.893784 -0.425765
+ 5.7e+10Hz 0.893448 -0.426455
+ 5.71e+10Hz 0.893112 -0.427144
+ 5.72e+10Hz 0.892775 -0.427833
+ 5.73e+10Hz 0.892438 -0.428522
+ 5.74e+10Hz 0.8921 -0.42921
+ 5.75e+10Hz 0.891762 -0.429898
+ 5.76e+10Hz 0.891424 -0.430586
+ 5.77e+10Hz 0.891085 -0.431274
+ 5.78e+10Hz 0.890745 -0.431961
+ 5.79e+10Hz 0.890405 -0.432648
+ 5.8e+10Hz 0.890065 -0.433335
+ 5.81e+10Hz 0.889724 -0.434022
+ 5.82e+10Hz 0.889383 -0.434708
+ 5.83e+10Hz 0.889041 -0.435394
+ 5.84e+10Hz 0.888699 -0.43608
+ 5.85e+10Hz 0.888356 -0.436766
+ 5.86e+10Hz 0.888013 -0.437451
+ 5.87e+10Hz 0.887669 -0.438137
+ 5.88e+10Hz 0.887325 -0.438821
+ 5.89e+10Hz 0.886981 -0.439506
+ 5.9e+10Hz 0.886636 -0.440191
+ 5.91e+10Hz 0.88629 -0.440875
+ 5.92e+10Hz 0.885944 -0.441559
+ 5.93e+10Hz 0.885598 -0.442242
+ 5.94e+10Hz 0.885251 -0.442926
+ 5.95e+10Hz 0.884904 -0.443609
+ 5.96e+10Hz 0.884556 -0.444292
+ 5.97e+10Hz 0.884208 -0.444975
+ 5.98e+10Hz 0.883859 -0.445658
+ 5.99e+10Hz 0.88351 -0.44634
+ 6e+10Hz 0.88316 -0.447022
+ 6.01e+10Hz 0.88281 -0.447704
+ 6.02e+10Hz 0.88246 -0.448385
+ 6.03e+10Hz 0.882108 -0.449067
+ 6.04e+10Hz 0.881757 -0.449748
+ 6.05e+10Hz 0.881405 -0.450429
+ 6.06e+10Hz 0.881052 -0.45111
+ 6.07e+10Hz 0.880699 -0.45179
+ 6.08e+10Hz 0.880346 -0.452471
+ 6.09e+10Hz 0.879992 -0.453151
+ 6.1e+10Hz 0.879637 -0.453831
+ 6.11e+10Hz 0.879282 -0.45451
+ 6.12e+10Hz 0.878927 -0.45519
+ 6.13e+10Hz 0.878571 -0.455869
+ 6.14e+10Hz 0.878215 -0.456548
+ 6.15e+10Hz 0.877858 -0.457227
+ 6.16e+10Hz 0.8775 -0.457905
+ 6.17e+10Hz 0.877142 -0.458584
+ 6.18e+10Hz 0.876784 -0.459262
+ 6.19e+10Hz 0.876425 -0.45994
+ 6.2e+10Hz 0.876066 -0.460618
+ 6.21e+10Hz 0.875706 -0.461295
+ 6.22e+10Hz 0.875345 -0.461972
+ 6.23e+10Hz 0.874984 -0.462649
+ 6.24e+10Hz 0.874623 -0.463326
+ 6.25e+10Hz 0.874261 -0.464003
+ 6.26e+10Hz 0.873899 -0.464679
+ 6.27e+10Hz 0.873536 -0.465356
+ 6.28e+10Hz 0.873172 -0.466032
+ 6.29e+10Hz 0.872808 -0.466707
+ 6.3e+10Hz 0.872444 -0.467383
+ 6.31e+10Hz 0.872079 -0.468058
+ 6.32e+10Hz 0.871713 -0.468734
+ 6.33e+10Hz 0.871347 -0.469408
+ 6.34e+10Hz 0.87098 -0.470083
+ 6.35e+10Hz 0.870613 -0.470758
+ 6.36e+10Hz 0.870245 -0.471432
+ 6.37e+10Hz 0.869877 -0.472106
+ 6.38e+10Hz 0.869508 -0.47278
+ 6.39e+10Hz 0.869139 -0.473453
+ 6.4e+10Hz 0.868769 -0.474127
+ 6.41e+10Hz 0.868399 -0.4748
+ 6.42e+10Hz 0.868028 -0.475473
+ 6.43e+10Hz 0.867657 -0.476145
+ 6.44e+10Hz 0.867285 -0.476818
+ 6.45e+10Hz 0.866912 -0.47749
+ 6.46e+10Hz 0.866539 -0.478162
+ 6.47e+10Hz 0.866165 -0.478834
+ 6.48e+10Hz 0.865791 -0.479506
+ 6.49e+10Hz 0.865416 -0.480177
+ 6.5e+10Hz 0.865041 -0.480848
+ 6.51e+10Hz 0.864665 -0.481519
+ 6.52e+10Hz 0.864289 -0.482189
+ 6.53e+10Hz 0.863912 -0.48286
+ 6.54e+10Hz 0.863534 -0.48353
+ 6.55e+10Hz 0.863156 -0.4842
+ 6.56e+10Hz 0.862778 -0.484869
+ 6.57e+10Hz 0.862399 -0.485539
+ 6.58e+10Hz 0.862019 -0.486208
+ 6.59e+10Hz 0.861639 -0.486877
+ 6.6e+10Hz 0.861258 -0.487546
+ 6.61e+10Hz 0.860876 -0.488214
+ 6.62e+10Hz 0.860494 -0.488882
+ 6.63e+10Hz 0.860112 -0.48955
+ 6.64e+10Hz 0.859729 -0.490218
+ 6.65e+10Hz 0.859345 -0.490885
+ 6.66e+10Hz 0.858961 -0.491552
+ 6.67e+10Hz 0.858576 -0.492219
+ 6.68e+10Hz 0.85819 -0.492886
+ 6.69e+10Hz 0.857804 -0.493552
+ 6.7e+10Hz 0.857418 -0.494218
+ 6.71e+10Hz 0.857031 -0.494884
+ 6.72e+10Hz 0.856643 -0.495549
+ 6.73e+10Hz 0.856255 -0.496214
+ 6.74e+10Hz 0.855866 -0.496879
+ 6.75e+10Hz 0.855476 -0.497544
+ 6.76e+10Hz 0.855086 -0.498208
+ 6.77e+10Hz 0.854696 -0.498872
+ 6.78e+10Hz 0.854305 -0.499536
+ 6.79e+10Hz 0.853913 -0.5002
+ 6.8e+10Hz 0.853521 -0.500863
+ 6.81e+10Hz 0.853128 -0.501526
+ 6.82e+10Hz 0.852734 -0.502189
+ 6.83e+10Hz 0.85234 -0.502851
+ 6.84e+10Hz 0.851946 -0.503513
+ 6.85e+10Hz 0.851551 -0.504175
+ 6.86e+10Hz 0.851155 -0.504836
+ 6.87e+10Hz 0.850759 -0.505497
+ 6.88e+10Hz 0.850362 -0.506158
+ 6.89e+10Hz 0.849964 -0.506819
+ 6.9e+10Hz 0.849566 -0.507479
+ 6.91e+10Hz 0.849168 -0.508139
+ 6.92e+10Hz 0.848768 -0.508798
+ 6.93e+10Hz 0.848369 -0.509457
+ 6.94e+10Hz 0.847968 -0.510116
+ 6.95e+10Hz 0.847567 -0.510775
+ 6.96e+10Hz 0.847166 -0.511433
+ 6.97e+10Hz 0.846764 -0.512091
+ 6.98e+10Hz 0.846361 -0.512749
+ 6.99e+10Hz 0.845958 -0.513406
+ 7e+10Hz 0.845554 -0.514063
+ 7.01e+10Hz 0.84515 -0.51472
+ 7.02e+10Hz 0.844745 -0.515376
+ 7.03e+10Hz 0.84434 -0.516032
+ 7.04e+10Hz 0.843934 -0.516687
+ 7.05e+10Hz 0.843527 -0.517343
+ 7.06e+10Hz 0.84312 -0.517998
+ 7.07e+10Hz 0.842712 -0.518652
+ 7.08e+10Hz 0.842304 -0.519306
+ 7.09e+10Hz 0.841895 -0.51996
+ 7.1e+10Hz 0.841486 -0.520614
+ 7.11e+10Hz 0.841076 -0.521267
+ 7.12e+10Hz 0.840665 -0.52192
+ 7.13e+10Hz 0.840254 -0.522572
+ 7.14e+10Hz 0.839843 -0.523224
+ 7.15e+10Hz 0.83943 -0.523876
+ 7.16e+10Hz 0.839018 -0.524527
+ 7.17e+10Hz 0.838605 -0.525178
+ 7.18e+10Hz 0.838191 -0.525829
+ 7.19e+10Hz 0.837776 -0.526479
+ 7.2e+10Hz 0.837362 -0.527129
+ 7.21e+10Hz 0.836946 -0.527779
+ 7.22e+10Hz 0.83653 -0.528428
+ 7.23e+10Hz 0.836114 -0.529077
+ 7.24e+10Hz 0.835697 -0.529725
+ 7.25e+10Hz 0.835279 -0.530373
+ 7.26e+10Hz 0.834861 -0.531021
+ 7.27e+10Hz 0.834442 -0.531668
+ 7.28e+10Hz 0.834023 -0.532315
+ 7.29e+10Hz 0.833604 -0.532961
+ 7.3e+10Hz 0.833183 -0.533608
+ 7.31e+10Hz 0.832763 -0.534253
+ 7.32e+10Hz 0.832341 -0.534899
+ 7.33e+10Hz 0.83192 -0.535544
+ 7.34e+10Hz 0.831497 -0.536188
+ 7.35e+10Hz 0.831075 -0.536833
+ 7.36e+10Hz 0.830651 -0.537476
+ 7.37e+10Hz 0.830227 -0.53812
+ 7.38e+10Hz 0.829803 -0.538763
+ 7.39e+10Hz 0.829378 -0.539406
+ 7.4e+10Hz 0.828953 -0.540048
+ 7.41e+10Hz 0.828527 -0.54069
+ 7.42e+10Hz 0.828101 -0.541331
+ 7.43e+10Hz 0.827674 -0.541972
+ 7.44e+10Hz 0.827246 -0.542613
+ 7.45e+10Hz 0.826818 -0.543254
+ 7.46e+10Hz 0.82639 -0.543894
+ 7.47e+10Hz 0.825961 -0.544533
+ 7.48e+10Hz 0.825532 -0.545172
+ 7.49e+10Hz 0.825102 -0.545811
+ 7.5e+10Hz 0.824672 -0.546449
+ 7.51e+10Hz 0.824241 -0.547087
+ 7.52e+10Hz 0.82381 -0.547725
+ 7.53e+10Hz 0.823378 -0.548362
+ 7.54e+10Hz 0.822946 -0.548999
+ 7.55e+10Hz 0.822513 -0.549636
+ 7.56e+10Hz 0.82208 -0.550272
+ 7.57e+10Hz 0.821646 -0.550907
+ 7.58e+10Hz 0.821212 -0.551542
+ 7.59e+10Hz 0.820777 -0.552177
+ 7.6e+10Hz 0.820342 -0.552812
+ 7.61e+10Hz 0.819906 -0.553446
+ 7.62e+10Hz 0.81947 -0.55408
+ 7.63e+10Hz 0.819034 -0.554713
+ 7.64e+10Hz 0.818597 -0.555346
+ 7.65e+10Hz 0.818159 -0.555978
+ 7.66e+10Hz 0.817721 -0.556611
+ 7.67e+10Hz 0.817283 -0.557242
+ 7.68e+10Hz 0.816844 -0.557874
+ 7.69e+10Hz 0.816405 -0.558505
+ 7.7e+10Hz 0.815965 -0.559135
+ 7.71e+10Hz 0.815525 -0.559765
+ 7.72e+10Hz 0.815084 -0.560395
+ 7.73e+10Hz 0.814643 -0.561025
+ 7.74e+10Hz 0.814202 -0.561654
+ 7.75e+10Hz 0.81376 -0.562282
+ 7.76e+10Hz 0.813317 -0.562911
+ 7.77e+10Hz 0.812874 -0.563539
+ 7.78e+10Hz 0.812431 -0.564166
+ 7.79e+10Hz 0.811987 -0.564793
+ 7.8e+10Hz 0.811543 -0.56542
+ 7.81e+10Hz 0.811098 -0.566047
+ 7.82e+10Hz 0.810653 -0.566673
+ 7.83e+10Hz 0.810208 -0.567298
+ 7.84e+10Hz 0.809762 -0.567924
+ 7.85e+10Hz 0.809315 -0.568549
+ 7.86e+10Hz 0.808868 -0.569173
+ 7.87e+10Hz 0.808421 -0.569797
+ 7.88e+10Hz 0.807973 -0.570421
+ 7.89e+10Hz 0.807525 -0.571044
+ 7.9e+10Hz 0.807076 -0.571668
+ 7.91e+10Hz 0.806627 -0.57229
+ 7.92e+10Hz 0.806178 -0.572913
+ 7.93e+10Hz 0.805728 -0.573535
+ 7.94e+10Hz 0.805278 -0.574156
+ 7.95e+10Hz 0.804827 -0.574777
+ 7.96e+10Hz 0.804376 -0.575398
+ 7.97e+10Hz 0.803924 -0.576019
+ 7.98e+10Hz 0.803472 -0.576639
+ 7.99e+10Hz 0.80302 -0.577259
+ 8e+10Hz 0.802567 -0.577878
+ 8.01e+10Hz 0.802113 -0.578497
+ 8.02e+10Hz 0.80166 -0.579116
+ 8.03e+10Hz 0.801205 -0.579734
+ 8.04e+10Hz 0.800751 -0.580352
+ 8.05e+10Hz 0.800296 -0.58097
+ 8.06e+10Hz 0.79984 -0.581587
+ 8.07e+10Hz 0.799384 -0.582204
+ 8.08e+10Hz 0.798928 -0.582821
+ 8.09e+10Hz 0.798471 -0.583437
+ 8.1e+10Hz 0.798014 -0.584053
+ 8.11e+10Hz 0.797556 -0.584669
+ 8.12e+10Hz 0.797098 -0.585284
+ 8.13e+10Hz 0.79664 -0.585899
+ 8.14e+10Hz 0.796181 -0.586514
+ 8.15e+10Hz 0.795721 -0.587128
+ 8.16e+10Hz 0.795262 -0.587742
+ 8.17e+10Hz 0.794801 -0.588355
+ 8.18e+10Hz 0.794341 -0.588969
+ 8.19e+10Hz 0.79388 -0.589581
+ 8.2e+10Hz 0.793418 -0.590194
+ 8.21e+10Hz 0.792956 -0.590806
+ 8.22e+10Hz 0.792494 -0.591418
+ 8.23e+10Hz 0.792031 -0.59203
+ 8.24e+10Hz 0.791568 -0.592641
+ 8.25e+10Hz 0.791104 -0.593252
+ 8.26e+10Hz 0.79064 -0.593862
+ 8.27e+10Hz 0.790176 -0.594472
+ 8.28e+10Hz 0.789711 -0.595082
+ 8.29e+10Hz 0.789245 -0.595692
+ 8.3e+10Hz 0.788779 -0.596301
+ 8.31e+10Hz 0.788313 -0.59691
+ 8.32e+10Hz 0.787846 -0.597518
+ 8.33e+10Hz 0.787379 -0.598127
+ 8.34e+10Hz 0.786912 -0.598735
+ 8.35e+10Hz 0.786444 -0.599342
+ 8.36e+10Hz 0.785975 -0.599949
+ 8.37e+10Hz 0.785506 -0.600556
+ 8.38e+10Hz 0.785037 -0.601163
+ 8.39e+10Hz 0.784567 -0.601769
+ 8.4e+10Hz 0.784097 -0.602375
+ 8.41e+10Hz 0.783626 -0.602981
+ 8.42e+10Hz 0.783155 -0.603586
+ 8.43e+10Hz 0.782683 -0.604191
+ 8.44e+10Hz 0.782211 -0.604796
+ 8.45e+10Hz 0.781739 -0.6054
+ 8.46e+10Hz 0.781266 -0.606004
+ 8.47e+10Hz 0.780792 -0.606608
+ 8.48e+10Hz 0.780319 -0.607211
+ 8.49e+10Hz 0.779844 -0.607814
+ 8.5e+10Hz 0.779369 -0.608417
+ 8.51e+10Hz 0.778894 -0.609019
+ 8.52e+10Hz 0.778419 -0.609621
+ 8.53e+10Hz 0.777942 -0.610223
+ 8.54e+10Hz 0.777466 -0.610825
+ 8.55e+10Hz 0.776989 -0.611426
+ 8.56e+10Hz 0.776511 -0.612026
+ 8.57e+10Hz 0.776033 -0.612627
+ 8.58e+10Hz 0.775555 -0.613227
+ 8.59e+10Hz 0.775076 -0.613827
+ 8.6e+10Hz 0.774596 -0.614426
+ 8.61e+10Hz 0.774117 -0.615025
+ 8.62e+10Hz 0.773636 -0.615624
+ 8.63e+10Hz 0.773155 -0.616223
+ 8.64e+10Hz 0.772674 -0.616821
+ 8.65e+10Hz 0.772192 -0.617419
+ 8.66e+10Hz 0.77171 -0.618016
+ 8.67e+10Hz 0.771228 -0.618614
+ 8.68e+10Hz 0.770744 -0.61921
+ 8.69e+10Hz 0.770261 -0.619807
+ 8.7e+10Hz 0.769777 -0.620403
+ 8.71e+10Hz 0.769292 -0.620999
+ 8.72e+10Hz 0.768807 -0.621594
+ 8.73e+10Hz 0.768321 -0.62219
+ 8.74e+10Hz 0.767835 -0.622784
+ 8.75e+10Hz 0.767349 -0.623379
+ 8.76e+10Hz 0.766862 -0.623973
+ 8.77e+10Hz 0.766374 -0.624567
+ 8.78e+10Hz 0.765886 -0.625161
+ 8.79e+10Hz 0.765398 -0.625754
+ 8.8e+10Hz 0.764909 -0.626346
+ 8.81e+10Hz 0.76442 -0.626939
+ 8.82e+10Hz 0.76393 -0.627531
+ 8.83e+10Hz 0.763439 -0.628123
+ 8.84e+10Hz 0.762948 -0.628714
+ 8.85e+10Hz 0.762457 -0.629305
+ 8.86e+10Hz 0.761965 -0.629896
+ 8.87e+10Hz 0.761473 -0.630487
+ 8.88e+10Hz 0.76098 -0.631077
+ 8.89e+10Hz 0.760487 -0.631666
+ 8.9e+10Hz 0.759993 -0.632256
+ 8.91e+10Hz 0.759499 -0.632845
+ 8.92e+10Hz 0.759004 -0.633433
+ 8.93e+10Hz 0.758508 -0.634021
+ 8.94e+10Hz 0.758013 -0.634609
+ 8.95e+10Hz 0.757516 -0.635197
+ 8.96e+10Hz 0.757019 -0.635784
+ 8.97e+10Hz 0.756522 -0.636371
+ 8.98e+10Hz 0.756024 -0.636957
+ 8.99e+10Hz 0.755526 -0.637543
+ 9e+10Hz 0.755027 -0.638129
+ 9.01e+10Hz 0.754528 -0.638715
+ 9.02e+10Hz 0.754028 -0.639299
+ 9.03e+10Hz 0.753528 -0.639884
+ 9.04e+10Hz 0.753027 -0.640468
+ 9.05e+10Hz 0.752526 -0.641052
+ 9.06e+10Hz 0.752024 -0.641636
+ 9.07e+10Hz 0.751522 -0.642219
+ 9.08e+10Hz 0.751019 -0.642801
+ 9.09e+10Hz 0.750516 -0.643384
+ 9.1e+10Hz 0.750012 -0.643966
+ 9.11e+10Hz 0.749508 -0.644547
+ 9.12e+10Hz 0.749003 -0.645128
+ 9.13e+10Hz 0.748498 -0.645709
+ 9.14e+10Hz 0.747992 -0.64629
+ 9.15e+10Hz 0.747486 -0.64687
+ 9.16e+10Hz 0.74698 -0.647449
+ 9.17e+10Hz 0.746472 -0.648028
+ 9.18e+10Hz 0.745965 -0.648607
+ 9.19e+10Hz 0.745456 -0.649186
+ 9.2e+10Hz 0.744948 -0.649764
+ 9.21e+10Hz 0.744439 -0.650341
+ 9.22e+10Hz 0.743929 -0.650919
+ 9.23e+10Hz 0.743419 -0.651495
+ 9.24e+10Hz 0.742908 -0.652072
+ 9.25e+10Hz 0.742397 -0.652648
+ 9.26e+10Hz 0.741885 -0.653223
+ 9.27e+10Hz 0.741373 -0.653799
+ 9.28e+10Hz 0.740861 -0.654373
+ 9.29e+10Hz 0.740347 -0.654948
+ 9.3e+10Hz 0.739834 -0.655522
+ 9.31e+10Hz 0.73932 -0.656095
+ 9.32e+10Hz 0.738805 -0.656668
+ 9.33e+10Hz 0.73829 -0.657241
+ 9.34e+10Hz 0.737775 -0.657813
+ 9.35e+10Hz 0.737259 -0.658385
+ 9.36e+10Hz 0.736742 -0.658956
+ 9.37e+10Hz 0.736225 -0.659527
+ 9.38e+10Hz 0.735708 -0.660098
+ 9.39e+10Hz 0.73519 -0.660668
+ 9.4e+10Hz 0.734671 -0.661238
+ 9.41e+10Hz 0.734153 -0.661807
+ 9.42e+10Hz 0.733633 -0.662376
+ 9.43e+10Hz 0.733113 -0.662944
+ 9.44e+10Hz 0.732593 -0.663512
+ 9.45e+10Hz 0.732072 -0.66408
+ 9.46e+10Hz 0.731551 -0.664647
+ 9.47e+10Hz 0.731029 -0.665214
+ 9.48e+10Hz 0.730507 -0.66578
+ 9.49e+10Hz 0.729984 -0.666346
+ 9.5e+10Hz 0.729461 -0.666911
+ 9.51e+10Hz 0.728938 -0.667476
+ 9.52e+10Hz 0.728414 -0.66804
+ 9.53e+10Hz 0.727889 -0.668605
+ 9.54e+10Hz 0.727364 -0.669168
+ 9.55e+10Hz 0.726839 -0.669731
+ 9.56e+10Hz 0.726313 -0.670294
+ 9.57e+10Hz 0.725787 -0.670856
+ 9.58e+10Hz 0.72526 -0.671418
+ 9.59e+10Hz 0.724733 -0.671979
+ 9.6e+10Hz 0.724205 -0.67254
+ 9.61e+10Hz 0.723677 -0.673101
+ 9.62e+10Hz 0.723148 -0.673661
+ 9.63e+10Hz 0.722619 -0.67422
+ 9.64e+10Hz 0.72209 -0.674779
+ 9.65e+10Hz 0.72156 -0.675338
+ 9.66e+10Hz 0.721029 -0.675896
+ 9.67e+10Hz 0.720498 -0.676454
+ 9.68e+10Hz 0.719967 -0.677011
+ 9.69e+10Hz 0.719436 -0.677568
+ 9.7e+10Hz 0.718903 -0.678125
+ 9.71e+10Hz 0.718371 -0.678681
+ 9.72e+10Hz 0.717838 -0.679236
+ 9.73e+10Hz 0.717304 -0.679791
+ 9.74e+10Hz 0.71677 -0.680346
+ 9.75e+10Hz 0.716236 -0.6809
+ 9.76e+10Hz 0.715701 -0.681453
+ 9.77e+10Hz 0.715166 -0.682007
+ 9.78e+10Hz 0.714631 -0.682559
+ 9.79e+10Hz 0.714095 -0.683112
+ 9.8e+10Hz 0.713558 -0.683664
+ 9.81e+10Hz 0.713021 -0.684215
+ 9.82e+10Hz 0.712484 -0.684766
+ 9.83e+10Hz 0.711946 -0.685316
+ 9.84e+10Hz 0.711408 -0.685866
+ 9.85e+10Hz 0.71087 -0.686416
+ 9.86e+10Hz 0.710331 -0.686965
+ 9.87e+10Hz 0.709791 -0.687514
+ 9.88e+10Hz 0.709252 -0.688062
+ 9.89e+10Hz 0.708712 -0.68861
+ 9.9e+10Hz 0.708171 -0.689157
+ 9.91e+10Hz 0.70763 -0.689704
+ 9.92e+10Hz 0.707089 -0.69025
+ 9.93e+10Hz 0.706547 -0.690796
+ 9.94e+10Hz 0.706004 -0.691342
+ 9.95e+10Hz 0.705462 -0.691887
+ 9.96e+10Hz 0.704919 -0.692431
+ 9.97e+10Hz 0.704375 -0.692975
+ 9.98e+10Hz 0.703832 -0.693519
+ 9.99e+10Hz 0.703287 -0.694062
+ 1e+11Hz 0.702743 -0.694605
+ 1.001e+11Hz 0.702198 -0.695147
+ 1.002e+11Hz 0.701652 -0.695689
+ 1.003e+11Hz 0.701106 -0.696231
+ 1.004e+11Hz 0.70056 -0.696772
+ 1.005e+11Hz 0.700014 -0.697312
+ 1.006e+11Hz 0.699467 -0.697852
+ 1.007e+11Hz 0.698919 -0.698392
+ 1.008e+11Hz 0.698372 -0.698931
+ 1.009e+11Hz 0.697823 -0.69947
+ 1.01e+11Hz 0.697275 -0.700008
+ 1.011e+11Hz 0.696726 -0.700546
+ 1.012e+11Hz 0.696177 -0.701083
+ 1.013e+11Hz 0.695627 -0.70162
+ 1.014e+11Hz 0.695077 -0.702157
+ 1.015e+11Hz 0.694526 -0.702693
+ 1.016e+11Hz 0.693975 -0.703229
+ 1.017e+11Hz 0.693424 -0.703764
+ 1.018e+11Hz 0.692873 -0.704299
+ 1.019e+11Hz 0.692321 -0.704833
+ 1.02e+11Hz 0.691768 -0.705367
+ 1.021e+11Hz 0.691215 -0.7059
+ 1.022e+11Hz 0.690662 -0.706433
+ 1.023e+11Hz 0.690109 -0.706966
+ 1.024e+11Hz 0.689555 -0.707498
+ 1.025e+11Hz 0.689 -0.70803
+ 1.026e+11Hz 0.688446 -0.708561
+ 1.027e+11Hz 0.687891 -0.709092
+ 1.028e+11Hz 0.687335 -0.709622
+ 1.029e+11Hz 0.686779 -0.710152
+ 1.03e+11Hz 0.686223 -0.710682
+ 1.031e+11Hz 0.685667 -0.711211
+ 1.032e+11Hz 0.68511 -0.71174
+ 1.033e+11Hz 0.684552 -0.712268
+ 1.034e+11Hz 0.683995 -0.712796
+ 1.035e+11Hz 0.683437 -0.713323
+ 1.036e+11Hz 0.682878 -0.71385
+ 1.037e+11Hz 0.682319 -0.714377
+ 1.038e+11Hz 0.68176 -0.714903
+ 1.039e+11Hz 0.681201 -0.715428
+ 1.04e+11Hz 0.680641 -0.715954
+ 1.041e+11Hz 0.68008 -0.716479
+ 1.042e+11Hz 0.67952 -0.717003
+ 1.043e+11Hz 0.678958 -0.717527
+ 1.044e+11Hz 0.678397 -0.718051
+ 1.045e+11Hz 0.677835 -0.718574
+ 1.046e+11Hz 0.677273 -0.719097
+ 1.047e+11Hz 0.67671 -0.719619
+ 1.048e+11Hz 0.676147 -0.720141
+ 1.049e+11Hz 0.675584 -0.720662
+ 1.05e+11Hz 0.67502 -0.721183
+ 1.051e+11Hz 0.674456 -0.721704
+ 1.052e+11Hz 0.673891 -0.722224
+ 1.053e+11Hz 0.673327 -0.722744
+ 1.054e+11Hz 0.672761 -0.723264
+ 1.055e+11Hz 0.672196 -0.723783
+ 1.056e+11Hz 0.67163 -0.724301
+ 1.057e+11Hz 0.671063 -0.72482
+ 1.058e+11Hz 0.670496 -0.725337
+ 1.059e+11Hz 0.669929 -0.725855
+ 1.06e+11Hz 0.669362 -0.726372
+ 1.061e+11Hz 0.668794 -0.726888
+ 1.062e+11Hz 0.668225 -0.727404
+ 1.063e+11Hz 0.667657 -0.72792
+ 1.064e+11Hz 0.667087 -0.728435
+ 1.065e+11Hz 0.666518 -0.72895
+ 1.066e+11Hz 0.665948 -0.729465
+ 1.067e+11Hz 0.665378 -0.729979
+ 1.068e+11Hz 0.664807 -0.730493
+ 1.069e+11Hz 0.664236 -0.731006
+ 1.07e+11Hz 0.663665 -0.731519
+ 1.071e+11Hz 0.663093 -0.732031
+ 1.072e+11Hz 0.662521 -0.732543
+ 1.073e+11Hz 0.661948 -0.733055
+ 1.074e+11Hz 0.661375 -0.733566
+ 1.075e+11Hz 0.660801 -0.734077
+ 1.076e+11Hz 0.660228 -0.734587
+ 1.077e+11Hz 0.659653 -0.735097
+ 1.078e+11Hz 0.659079 -0.735607
+ 1.079e+11Hz 0.658504 -0.736116
+ 1.08e+11Hz 0.657928 -0.736625
+ 1.081e+11Hz 0.657353 -0.737133
+ 1.082e+11Hz 0.656776 -0.737641
+ 1.083e+11Hz 0.6562 -0.738148
+ 1.084e+11Hz 0.655623 -0.738655
+ 1.085e+11Hz 0.655045 -0.739162
+ 1.086e+11Hz 0.654468 -0.739668
+ 1.087e+11Hz 0.653889 -0.740174
+ 1.088e+11Hz 0.653311 -0.74068
+ 1.089e+11Hz 0.652732 -0.741185
+ 1.09e+11Hz 0.652152 -0.741689
+ 1.091e+11Hz 0.651573 -0.742194
+ 1.092e+11Hz 0.650992 -0.742697
+ 1.093e+11Hz 0.650412 -0.743201
+ 1.094e+11Hz 0.649831 -0.743704
+ 1.095e+11Hz 0.649249 -0.744206
+ 1.096e+11Hz 0.648667 -0.744708
+ 1.097e+11Hz 0.648085 -0.74521
+ 1.098e+11Hz 0.647502 -0.745711
+ 1.099e+11Hz 0.646919 -0.746212
+ 1.1e+11Hz 0.646336 -0.746713
+ 1.101e+11Hz 0.645752 -0.747213
+ 1.102e+11Hz 0.645167 -0.747712
+ 1.103e+11Hz 0.644583 -0.748212
+ 1.104e+11Hz 0.643998 -0.74871
+ 1.105e+11Hz 0.643412 -0.749209
+ 1.106e+11Hz 0.642826 -0.749706
+ 1.107e+11Hz 0.64224 -0.750204
+ 1.108e+11Hz 0.641653 -0.750701
+ 1.109e+11Hz 0.641065 -0.751198
+ 1.11e+11Hz 0.640478 -0.751694
+ 1.111e+11Hz 0.63989 -0.75219
+ 1.112e+11Hz 0.639301 -0.752685
+ 1.113e+11Hz 0.638712 -0.75318
+ 1.114e+11Hz 0.638123 -0.753674
+ 1.115e+11Hz 0.637533 -0.754168
+ 1.116e+11Hz 0.636943 -0.754662
+ 1.117e+11Hz 0.636352 -0.755155
+ 1.118e+11Hz 0.635761 -0.755648
+ 1.119e+11Hz 0.63517 -0.75614
+ 1.12e+11Hz 0.634578 -0.756632
+ 1.121e+11Hz 0.633986 -0.757123
+ 1.122e+11Hz 0.633393 -0.757614
+ 1.123e+11Hz 0.6328 -0.758105
+ 1.124e+11Hz 0.632206 -0.758595
+ 1.125e+11Hz 0.631612 -0.759084
+ 1.126e+11Hz 0.631018 -0.759573
+ 1.127e+11Hz 0.630423 -0.760062
+ 1.128e+11Hz 0.629828 -0.76055
+ 1.129e+11Hz 0.629232 -0.761038
+ 1.13e+11Hz 0.628636 -0.761526
+ 1.131e+11Hz 0.628039 -0.762012
+ 1.132e+11Hz 0.627442 -0.762499
+ 1.133e+11Hz 0.626845 -0.762985
+ 1.134e+11Hz 0.626247 -0.76347
+ 1.135e+11Hz 0.625649 -0.763955
+ 1.136e+11Hz 0.62505 -0.76444
+ 1.137e+11Hz 0.624451 -0.764924
+ 1.138e+11Hz 0.623852 -0.765408
+ 1.139e+11Hz 0.623252 -0.765891
+ 1.14e+11Hz 0.622651 -0.766374
+ 1.141e+11Hz 0.622051 -0.766856
+ 1.142e+11Hz 0.621449 -0.767338
+ 1.143e+11Hz 0.620848 -0.767819
+ 1.144e+11Hz 0.620246 -0.7683
+ 1.145e+11Hz 0.619643 -0.76878
+ 1.146e+11Hz 0.61904 -0.76926
+ 1.147e+11Hz 0.618437 -0.76974
+ 1.148e+11Hz 0.617833 -0.770218
+ 1.149e+11Hz 0.617229 -0.770697
+ 1.15e+11Hz 0.616625 -0.771175
+ 1.151e+11Hz 0.61602 -0.771652
+ 1.152e+11Hz 0.615414 -0.772129
+ 1.153e+11Hz 0.614808 -0.772606
+ 1.154e+11Hz 0.614202 -0.773082
+ 1.155e+11Hz 0.613596 -0.773557
+ 1.156e+11Hz 0.612989 -0.774032
+ 1.157e+11Hz 0.612381 -0.774507
+ 1.158e+11Hz 0.611773 -0.774981
+ 1.159e+11Hz 0.611165 -0.775455
+ 1.16e+11Hz 0.610556 -0.775928
+ 1.161e+11Hz 0.609947 -0.7764
+ 1.162e+11Hz 0.609338 -0.776872
+ 1.163e+11Hz 0.608728 -0.777344
+ 1.164e+11Hz 0.608117 -0.777815
+ 1.165e+11Hz 0.607507 -0.778286
+ 1.166e+11Hz 0.606895 -0.778756
+ 1.167e+11Hz 0.606284 -0.779225
+ 1.168e+11Hz 0.605672 -0.779694
+ 1.169e+11Hz 0.60506 -0.780163
+ 1.17e+11Hz 0.604447 -0.780631
+ 1.171e+11Hz 0.603834 -0.781099
+ 1.172e+11Hz 0.60322 -0.781566
+ 1.173e+11Hz 0.602606 -0.782032
+ 1.174e+11Hz 0.601992 -0.782498
+ 1.175e+11Hz 0.601377 -0.782964
+ 1.176e+11Hz 0.600762 -0.783429
+ 1.177e+11Hz 0.600146 -0.783893
+ 1.178e+11Hz 0.59953 -0.784357
+ 1.179e+11Hz 0.598914 -0.784821
+ 1.18e+11Hz 0.598297 -0.785284
+ 1.181e+11Hz 0.59768 -0.785746
+ 1.182e+11Hz 0.597063 -0.786208
+ 1.183e+11Hz 0.596445 -0.786669
+ 1.184e+11Hz 0.595827 -0.78713
+ 1.185e+11Hz 0.595208 -0.78759
+ 1.186e+11Hz 0.594589 -0.78805
+ 1.187e+11Hz 0.593969 -0.78851
+ 1.188e+11Hz 0.59335 -0.788968
+ 1.189e+11Hz 0.592729 -0.789427
+ 1.19e+11Hz 0.592109 -0.789884
+ 1.191e+11Hz 0.591488 -0.790342
+ 1.192e+11Hz 0.590867 -0.790798
+ 1.193e+11Hz 0.590245 -0.791254
+ 1.194e+11Hz 0.589623 -0.79171
+ 1.195e+11Hz 0.589001 -0.792165
+ 1.196e+11Hz 0.588378 -0.79262
+ 1.197e+11Hz 0.587755 -0.793074
+ 1.198e+11Hz 0.587131 -0.793527
+ 1.199e+11Hz 0.586507 -0.79398
+ 1.2e+11Hz 0.585883 -0.794433
+ 1.201e+11Hz 0.585258 -0.794885
+ 1.202e+11Hz 0.584633 -0.795336
+ 1.203e+11Hz 0.584008 -0.795787
+ 1.204e+11Hz 0.583382 -0.796237
+ 1.205e+11Hz 0.582756 -0.796687
+ 1.206e+11Hz 0.58213 -0.797137
+ 1.207e+11Hz 0.581503 -0.797585
+ 1.208e+11Hz 0.580876 -0.798033
+ 1.209e+11Hz 0.580248 -0.798481
+ 1.21e+11Hz 0.579621 -0.798928
+ 1.211e+11Hz 0.578993 -0.799375
+ 1.212e+11Hz 0.578364 -0.799821
+ 1.213e+11Hz 0.577735 -0.800267
+ 1.214e+11Hz 0.577106 -0.800712
+ 1.215e+11Hz 0.576476 -0.801156
+ 1.216e+11Hz 0.575846 -0.8016
+ 1.217e+11Hz 0.575216 -0.802044
+ 1.218e+11Hz 0.574586 -0.802487
+ 1.219e+11Hz 0.573955 -0.802929
+ 1.22e+11Hz 0.573324 -0.803371
+ 1.221e+11Hz 0.572692 -0.803812
+ 1.222e+11Hz 0.57206 -0.804253
+ 1.223e+11Hz 0.571428 -0.804693
+ 1.224e+11Hz 0.570795 -0.805133
+ 1.225e+11Hz 0.570162 -0.805572
+ 1.226e+11Hz 0.569529 -0.806011
+ 1.227e+11Hz 0.568895 -0.806449
+ 1.228e+11Hz 0.568261 -0.806887
+ 1.229e+11Hz 0.567627 -0.807324
+ 1.23e+11Hz 0.566993 -0.807761
+ 1.231e+11Hz 0.566358 -0.808197
+ 1.232e+11Hz 0.565723 -0.808632
+ 1.233e+11Hz 0.565087 -0.809067
+ 1.234e+11Hz 0.564451 -0.809502
+ 1.235e+11Hz 0.563815 -0.809936
+ 1.236e+11Hz 0.563178 -0.810369
+ 1.237e+11Hz 0.562542 -0.810802
+ 1.238e+11Hz 0.561904 -0.811234
+ 1.239e+11Hz 0.561267 -0.811666
+ 1.24e+11Hz 0.560629 -0.812098
+ 1.241e+11Hz 0.559991 -0.812528
+ 1.242e+11Hz 0.559353 -0.812959
+ 1.243e+11Hz 0.558714 -0.813389
+ 1.244e+11Hz 0.558075 -0.813818
+ 1.245e+11Hz 0.557436 -0.814247
+ 1.246e+11Hz 0.556796 -0.814675
+ 1.247e+11Hz 0.556156 -0.815103
+ 1.248e+11Hz 0.555516 -0.81553
+ 1.249e+11Hz 0.554875 -0.815956
+ 1.25e+11Hz 0.554234 -0.816383
+ 1.251e+11Hz 0.553593 -0.816808
+ 1.252e+11Hz 0.552951 -0.817233
+ 1.253e+11Hz 0.552309 -0.817658
+ 1.254e+11Hz 0.551667 -0.818082
+ 1.255e+11Hz 0.551025 -0.818506
+ 1.256e+11Hz 0.550382 -0.818929
+ 1.257e+11Hz 0.549739 -0.819351
+ 1.258e+11Hz 0.549096 -0.819773
+ 1.259e+11Hz 0.548452 -0.820195
+ 1.26e+11Hz 0.547808 -0.820616
+ 1.261e+11Hz 0.547164 -0.821037
+ 1.262e+11Hz 0.546519 -0.821457
+ 1.263e+11Hz 0.545874 -0.821876
+ 1.264e+11Hz 0.545229 -0.822295
+ 1.265e+11Hz 0.544583 -0.822714
+ 1.266e+11Hz 0.543937 -0.823132
+ 1.267e+11Hz 0.543291 -0.823549
+ 1.268e+11Hz 0.542645 -0.823966
+ 1.269e+11Hz 0.541998 -0.824383
+ 1.27e+11Hz 0.541351 -0.824799
+ 1.271e+11Hz 0.540704 -0.825214
+ 1.272e+11Hz 0.540056 -0.825629
+ 1.273e+11Hz 0.539408 -0.826044
+ 1.274e+11Hz 0.53876 -0.826457
+ 1.275e+11Hz 0.538111 -0.826871
+ 1.276e+11Hz 0.537462 -0.827284
+ 1.277e+11Hz 0.536813 -0.827696
+ 1.278e+11Hz 0.536164 -0.828108
+ 1.279e+11Hz 0.535514 -0.82852
+ 1.28e+11Hz 0.534864 -0.828931
+ 1.281e+11Hz 0.534213 -0.829341
+ 1.282e+11Hz 0.533562 -0.829751
+ 1.283e+11Hz 0.532911 -0.830161
+ 1.284e+11Hz 0.53226 -0.83057
+ 1.285e+11Hz 0.531608 -0.830978
+ 1.286e+11Hz 0.530956 -0.831386
+ 1.287e+11Hz 0.530304 -0.831794
+ 1.288e+11Hz 0.529652 -0.832201
+ 1.289e+11Hz 0.528999 -0.832607
+ 1.29e+11Hz 0.528346 -0.833013
+ 1.291e+11Hz 0.527692 -0.833419
+ 1.292e+11Hz 0.527038 -0.833824
+ 1.293e+11Hz 0.526384 -0.834228
+ 1.294e+11Hz 0.52573 -0.834632
+ 1.295e+11Hz 0.525075 -0.835036
+ 1.296e+11Hz 0.52442 -0.835439
+ 1.297e+11Hz 0.523764 -0.835841
+ 1.298e+11Hz 0.523109 -0.836244
+ 1.299e+11Hz 0.522453 -0.836645
+ 1.3e+11Hz 0.521796 -0.837046
+ 1.301e+11Hz 0.52114 -0.837447
+ 1.302e+11Hz 0.520483 -0.837847
+ 1.303e+11Hz 0.519826 -0.838246
+ 1.304e+11Hz 0.519168 -0.838645
+ 1.305e+11Hz 0.51851 -0.839044
+ 1.306e+11Hz 0.517852 -0.839442
+ 1.307e+11Hz 0.517193 -0.83984
+ 1.308e+11Hz 0.516535 -0.840237
+ 1.309e+11Hz 0.515875 -0.840634
+ 1.31e+11Hz 0.515216 -0.84103
+ 1.311e+11Hz 0.514556 -0.841425
+ 1.312e+11Hz 0.513896 -0.84182
+ 1.313e+11Hz 0.513236 -0.842215
+ 1.314e+11Hz 0.512575 -0.842609
+ 1.315e+11Hz 0.511914 -0.843003
+ 1.316e+11Hz 0.511252 -0.843396
+ 1.317e+11Hz 0.510591 -0.843789
+ 1.318e+11Hz 0.509928 -0.844181
+ 1.319e+11Hz 0.509266 -0.844572
+ 1.32e+11Hz 0.508603 -0.844964
+ 1.321e+11Hz 0.50794 -0.845354
+ 1.322e+11Hz 0.507277 -0.845744
+ 1.323e+11Hz 0.506613 -0.846134
+ 1.324e+11Hz 0.505949 -0.846523
+ 1.325e+11Hz 0.505285 -0.846912
+ 1.326e+11Hz 0.50462 -0.8473
+ 1.327e+11Hz 0.503955 -0.847688
+ 1.328e+11Hz 0.50329 -0.848075
+ 1.329e+11Hz 0.502624 -0.848461
+ 1.33e+11Hz 0.501958 -0.848847
+ 1.331e+11Hz 0.501292 -0.849233
+ 1.332e+11Hz 0.500625 -0.849618
+ 1.333e+11Hz 0.499958 -0.850003
+ 1.334e+11Hz 0.499291 -0.850387
+ 1.335e+11Hz 0.498623 -0.85077
+ 1.336e+11Hz 0.497955 -0.851154
+ 1.337e+11Hz 0.497287 -0.851536
+ 1.338e+11Hz 0.496618 -0.851918
+ 1.339e+11Hz 0.495949 -0.8523
+ 1.34e+11Hz 0.49528 -0.852681
+ 1.341e+11Hz 0.49461 -0.853061
+ 1.342e+11Hz 0.49394 -0.853441
+ 1.343e+11Hz 0.49327 -0.853821
+ 1.344e+11Hz 0.492599 -0.8542
+ 1.345e+11Hz 0.491928 -0.854578
+ 1.346e+11Hz 0.491257 -0.854956
+ 1.347e+11Hz 0.490585 -0.855333
+ 1.348e+11Hz 0.489913 -0.85571
+ 1.349e+11Hz 0.489241 -0.856087
+ 1.35e+11Hz 0.488568 -0.856462
+ 1.351e+11Hz 0.487895 -0.856838
+ 1.352e+11Hz 0.487222 -0.857212
+ 1.353e+11Hz 0.486548 -0.857587
+ 1.354e+11Hz 0.485874 -0.85796
+ 1.355e+11Hz 0.4852 -0.858334
+ 1.356e+11Hz 0.484525 -0.858706
+ 1.357e+11Hz 0.48385 -0.859078
+ 1.358e+11Hz 0.483175 -0.85945
+ 1.359e+11Hz 0.482499 -0.859821
+ 1.36e+11Hz 0.481823 -0.860191
+ 1.361e+11Hz 0.481147 -0.860561
+ 1.362e+11Hz 0.48047 -0.860931
+ 1.363e+11Hz 0.479793 -0.8613
+ 1.364e+11Hz 0.479116 -0.861668
+ 1.365e+11Hz 0.478438 -0.862036
+ 1.366e+11Hz 0.47776 -0.862403
+ 1.367e+11Hz 0.477082 -0.86277
+ 1.368e+11Hz 0.476403 -0.863136
+ 1.369e+11Hz 0.475724 -0.863501
+ 1.37e+11Hz 0.475044 -0.863866
+ 1.371e+11Hz 0.474365 -0.864231
+ 1.372e+11Hz 0.473685 -0.864595
+ 1.373e+11Hz 0.473004 -0.864958
+ 1.374e+11Hz 0.472323 -0.865321
+ 1.375e+11Hz 0.471642 -0.865683
+ 1.376e+11Hz 0.470961 -0.866045
+ 1.377e+11Hz 0.470279 -0.866406
+ 1.378e+11Hz 0.469597 -0.866767
+ 1.379e+11Hz 0.468915 -0.867127
+ 1.38e+11Hz 0.468232 -0.867486
+ 1.381e+11Hz 0.467549 -0.867845
+ 1.382e+11Hz 0.466866 -0.868203
+ 1.383e+11Hz 0.466182 -0.868561
+ 1.384e+11Hz 0.465498 -0.868918
+ 1.385e+11Hz 0.464814 -0.869275
+ 1.386e+11Hz 0.464129 -0.869631
+ 1.387e+11Hz 0.463444 -0.869986
+ 1.388e+11Hz 0.462759 -0.870341
+ 1.389e+11Hz 0.462073 -0.870696
+ 1.39e+11Hz 0.461387 -0.871049
+ 1.391e+11Hz 0.460701 -0.871403
+ 1.392e+11Hz 0.460014 -0.871755
+ 1.393e+11Hz 0.459328 -0.872107
+ 1.394e+11Hz 0.45864 -0.872459
+ 1.395e+11Hz 0.457953 -0.872809
+ 1.396e+11Hz 0.457265 -0.87316
+ 1.397e+11Hz 0.456577 -0.873509
+ 1.398e+11Hz 0.455888 -0.873858
+ 1.399e+11Hz 0.4552 -0.874207
+ 1.4e+11Hz 0.45451 -0.874555
+ 1.401e+11Hz 0.453821 -0.874902
+ 1.402e+11Hz 0.453131 -0.875249
+ 1.403e+11Hz 0.452441 -0.875595
+ 1.404e+11Hz 0.451751 -0.87594
+ 1.405e+11Hz 0.45106 -0.876285
+ 1.406e+11Hz 0.450369 -0.87663
+ 1.407e+11Hz 0.449678 -0.876974
+ 1.408e+11Hz 0.448987 -0.877317
+ 1.409e+11Hz 0.448295 -0.877659
+ 1.41e+11Hz 0.447603 -0.878001
+ 1.411e+11Hz 0.44691 -0.878343
+ 1.412e+11Hz 0.446218 -0.878683
+ 1.413e+11Hz 0.445524 -0.879023
+ 1.414e+11Hz 0.444831 -0.879363
+ 1.415e+11Hz 0.444138 -0.879702
+ 1.416e+11Hz 0.443444 -0.88004
+ 1.417e+11Hz 0.44275 -0.880378
+ 1.418e+11Hz 0.442055 -0.880715
+ 1.419e+11Hz 0.44136 -0.881052
+ 1.42e+11Hz 0.440665 -0.881388
+ 1.421e+11Hz 0.43997 -0.881723
+ 1.422e+11Hz 0.439274 -0.882058
+ 1.423e+11Hz 0.438578 -0.882392
+ 1.424e+11Hz 0.437882 -0.882725
+ 1.425e+11Hz 0.437186 -0.883058
+ 1.426e+11Hz 0.436489 -0.883391
+ 1.427e+11Hz 0.435792 -0.883722
+ 1.428e+11Hz 0.435095 -0.884053
+ 1.429e+11Hz 0.434397 -0.884384
+ 1.43e+11Hz 0.433699 -0.884714
+ 1.431e+11Hz 0.433001 -0.885043
+ 1.432e+11Hz 0.432303 -0.885371
+ 1.433e+11Hz 0.431604 -0.885699
+ 1.434e+11Hz 0.430906 -0.886027
+ 1.435e+11Hz 0.430206 -0.886354
+ 1.436e+11Hz 0.429507 -0.88668
+ 1.437e+11Hz 0.428807 -0.887005
+ 1.438e+11Hz 0.428107 -0.88733
+ 1.439e+11Hz 0.427407 -0.887655
+ 1.44e+11Hz 0.426707 -0.887978
+ 1.441e+11Hz 0.426006 -0.888301
+ 1.442e+11Hz 0.425305 -0.888624
+ 1.443e+11Hz 0.424604 -0.888946
+ 1.444e+11Hz 0.423903 -0.889267
+ 1.445e+11Hz 0.423201 -0.889588
+ 1.446e+11Hz 0.422499 -0.889908
+ 1.447e+11Hz 0.421797 -0.890227
+ 1.448e+11Hz 0.421094 -0.890546
+ 1.449e+11Hz 0.420392 -0.890864
+ 1.45e+11Hz 0.419689 -0.891182
+ 1.451e+11Hz 0.418986 -0.891499
+ 1.452e+11Hz 0.418282 -0.891815
+ 1.453e+11Hz 0.417579 -0.892131
+ 1.454e+11Hz 0.416875 -0.892446
+ 1.455e+11Hz 0.416171 -0.89276
+ 1.456e+11Hz 0.415466 -0.893074
+ 1.457e+11Hz 0.414762 -0.893387
+ 1.458e+11Hz 0.414057 -0.8937
+ 1.459e+11Hz 0.413352 -0.894012
+ 1.46e+11Hz 0.412647 -0.894323
+ 1.461e+11Hz 0.411941 -0.894634
+ 1.462e+11Hz 0.411235 -0.894944
+ 1.463e+11Hz 0.410529 -0.895254
+ 1.464e+11Hz 0.409823 -0.895563
+ 1.465e+11Hz 0.409117 -0.895871
+ 1.466e+11Hz 0.40841 -0.896179
+ 1.467e+11Hz 0.407703 -0.896486
+ 1.468e+11Hz 0.406996 -0.896793
+ 1.469e+11Hz 0.406289 -0.897099
+ 1.47e+11Hz 0.405581 -0.897404
+ 1.471e+11Hz 0.404874 -0.897709
+ 1.472e+11Hz 0.404166 -0.898013
+ 1.473e+11Hz 0.403458 -0.898316
+ 1.474e+11Hz 0.402749 -0.898619
+ 1.475e+11Hz 0.402041 -0.898922
+ 1.476e+11Hz 0.401332 -0.899223
+ 1.477e+11Hz 0.400623 -0.899524
+ 1.478e+11Hz 0.399914 -0.899825
+ 1.479e+11Hz 0.399204 -0.900125
+ 1.48e+11Hz 0.398494 -0.900424
+ 1.481e+11Hz 0.397785 -0.900723
+ 1.482e+11Hz 0.397074 -0.901021
+ 1.483e+11Hz 0.396364 -0.901318
+ 1.484e+11Hz 0.395654 -0.901615
+ 1.485e+11Hz 0.394943 -0.901911
+ 1.486e+11Hz 0.394232 -0.902207
+ 1.487e+11Hz 0.393521 -0.902502
+ 1.488e+11Hz 0.39281 -0.902796
+ 1.489e+11Hz 0.392098 -0.90309
+ 1.49e+11Hz 0.391386 -0.903383
+ 1.491e+11Hz 0.390675 -0.903676
+ 1.492e+11Hz 0.389962 -0.903968
+ 1.493e+11Hz 0.38925 -0.904259
+ 1.494e+11Hz 0.388538 -0.90455
+ 1.495e+11Hz 0.387825 -0.90484
+ 1.496e+11Hz 0.387112 -0.90513
+ 1.497e+11Hz 0.386399 -0.905419
+ 1.498e+11Hz 0.385685 -0.905707
+ 1.499e+11Hz 0.384972 -0.905995
+ 1.5e+11Hz 0.384258 -0.906282
+ 1.501e+11Hz 0.383544 -0.906569
+ 1.502e+11Hz 0.38283 -0.906855
+ 1.503e+11Hz 0.382116 -0.907141
+ 1.504e+11Hz 0.381401 -0.907425
+ 1.505e+11Hz 0.380686 -0.90771
+ 1.506e+11Hz 0.379972 -0.907993
+ 1.507e+11Hz 0.379256 -0.908276
+ 1.508e+11Hz 0.378541 -0.908559
+ 1.509e+11Hz 0.377826 -0.908841
+ 1.51e+11Hz 0.37711 -0.909122
+ 1.511e+11Hz 0.376394 -0.909403
+ 1.512e+11Hz 0.375678 -0.909683
+ 1.513e+11Hz 0.374962 -0.909962
+ 1.514e+11Hz 0.374245 -0.910241
+ 1.515e+11Hz 0.373528 -0.91052
+ 1.516e+11Hz 0.372811 -0.910797
+ 1.517e+11Hz 0.372094 -0.911074
+ 1.518e+11Hz 0.371377 -0.911351
+ 1.519e+11Hz 0.37066 -0.911627
+ 1.52e+11Hz 0.369942 -0.911902
+ 1.521e+11Hz 0.369224 -0.912177
+ 1.522e+11Hz 0.368506 -0.912451
+ 1.523e+11Hz 0.367788 -0.912725
+ 1.524e+11Hz 0.367069 -0.912998
+ 1.525e+11Hz 0.366351 -0.91327
+ 1.526e+11Hz 0.365632 -0.913542
+ 1.527e+11Hz 0.364913 -0.913813
+ 1.528e+11Hz 0.364193 -0.914084
+ 1.529e+11Hz 0.363474 -0.914354
+ 1.53e+11Hz 0.362754 -0.914623
+ 1.531e+11Hz 0.362034 -0.914892
+ 1.532e+11Hz 0.361314 -0.915161
+ 1.533e+11Hz 0.360594 -0.915428
+ 1.534e+11Hz 0.359874 -0.915695
+ 1.535e+11Hz 0.359153 -0.915962
+ 1.536e+11Hz 0.358432 -0.916228
+ 1.537e+11Hz 0.357711 -0.916493
+ 1.538e+11Hz 0.35699 -0.916758
+ 1.539e+11Hz 0.356269 -0.917022
+ 1.54e+11Hz 0.355547 -0.917285
+ 1.541e+11Hz 0.354825 -0.917548
+ 1.542e+11Hz 0.354103 -0.91781
+ 1.543e+11Hz 0.353381 -0.918072
+ 1.544e+11Hz 0.352659 -0.918333
+ 1.545e+11Hz 0.351936 -0.918594
+ 1.546e+11Hz 0.351213 -0.918854
+ 1.547e+11Hz 0.35049 -0.919113
+ 1.548e+11Hz 0.349767 -0.919372
+ 1.549e+11Hz 0.349044 -0.91963
+ 1.55e+11Hz 0.34832 -0.919888
+ 1.551e+11Hz 0.347596 -0.920144
+ 1.552e+11Hz 0.346872 -0.920401
+ 1.553e+11Hz 0.346148 -0.920657
+ 1.554e+11Hz 0.345424 -0.920912
+ 1.555e+11Hz 0.344699 -0.921166
+ 1.556e+11Hz 0.343974 -0.92142
+ 1.557e+11Hz 0.343249 -0.921673
+ 1.558e+11Hz 0.342524 -0.921926
+ 1.559e+11Hz 0.341799 -0.922178
+ 1.56e+11Hz 0.341073 -0.92243
+ 1.561e+11Hz 0.340348 -0.922681
+ 1.562e+11Hz 0.339622 -0.922931
+ 1.563e+11Hz 0.338895 -0.923181
+ 1.564e+11Hz 0.338169 -0.92343
+ 1.565e+11Hz 0.337443 -0.923678
+ 1.566e+11Hz 0.336716 -0.923926
+ 1.567e+11Hz 0.335989 -0.924173
+ 1.568e+11Hz 0.335262 -0.92442
+ 1.569e+11Hz 0.334535 -0.924666
+ 1.57e+11Hz 0.333807 -0.924911
+ 1.571e+11Hz 0.333079 -0.925156
+ 1.572e+11Hz 0.332351 -0.9254
+ 1.573e+11Hz 0.331623 -0.925643
+ 1.574e+11Hz 0.330895 -0.925886
+ 1.575e+11Hz 0.330167 -0.926129
+ 1.576e+11Hz 0.329438 -0.92637
+ 1.577e+11Hz 0.328709 -0.926611
+ 1.578e+11Hz 0.32798 -0.926852
+ 1.579e+11Hz 0.327251 -0.927091
+ 1.58e+11Hz 0.326521 -0.927331
+ 1.581e+11Hz 0.325792 -0.927569
+ 1.582e+11Hz 0.325062 -0.927807
+ 1.583e+11Hz 0.324332 -0.928044
+ 1.584e+11Hz 0.323602 -0.928281
+ 1.585e+11Hz 0.322872 -0.928517
+ 1.586e+11Hz 0.322141 -0.928752
+ 1.587e+11Hz 0.32141 -0.928987
+ 1.588e+11Hz 0.320679 -0.929221
+ 1.589e+11Hz 0.319948 -0.929454
+ 1.59e+11Hz 0.319217 -0.929687
+ 1.591e+11Hz 0.318486 -0.929919
+ 1.592e+11Hz 0.317754 -0.930151
+ 1.593e+11Hz 0.317022 -0.930382
+ 1.594e+11Hz 0.31629 -0.930612
+ 1.595e+11Hz 0.315558 -0.930842
+ 1.596e+11Hz 0.314826 -0.931071
+ 1.597e+11Hz 0.314093 -0.931299
+ 1.598e+11Hz 0.313361 -0.931526
+ 1.599e+11Hz 0.312628 -0.931753
+ 1.6e+11Hz 0.311895 -0.93198
+ 1.601e+11Hz 0.311162 -0.932206
+ 1.602e+11Hz 0.310428 -0.932431
+ 1.603e+11Hz 0.309695 -0.932655
+ 1.604e+11Hz 0.308961 -0.932879
+ 1.605e+11Hz 0.308227 -0.933102
+ 1.606e+11Hz 0.307493 -0.933324
+ 1.607e+11Hz 0.306759 -0.933546
+ 1.608e+11Hz 0.306025 -0.933767
+ 1.609e+11Hz 0.305291 -0.933988
+ 1.61e+11Hz 0.304556 -0.934207
+ 1.611e+11Hz 0.303821 -0.934426
+ 1.612e+11Hz 0.303086 -0.934645
+ 1.613e+11Hz 0.302351 -0.934863
+ 1.614e+11Hz 0.301616 -0.93508
+ 1.615e+11Hz 0.300881 -0.935296
+ 1.616e+11Hz 0.300145 -0.935512
+ 1.617e+11Hz 0.299409 -0.935727
+ 1.618e+11Hz 0.298674 -0.935942
+ 1.619e+11Hz 0.297938 -0.936155
+ 1.62e+11Hz 0.297202 -0.936369
+ 1.621e+11Hz 0.296465 -0.936581
+ 1.622e+11Hz 0.295729 -0.936793
+ 1.623e+11Hz 0.294993 -0.937004
+ 1.624e+11Hz 0.294256 -0.937214
+ 1.625e+11Hz 0.293519 -0.937424
+ 1.626e+11Hz 0.292782 -0.937633
+ 1.627e+11Hz 0.292046 -0.937842
+ 1.628e+11Hz 0.291308 -0.938049
+ 1.629e+11Hz 0.290571 -0.938256
+ 1.63e+11Hz 0.289834 -0.938463
+ 1.631e+11Hz 0.289096 -0.938668
+ 1.632e+11Hz 0.288359 -0.938873
+ 1.633e+11Hz 0.287621 -0.939078
+ 1.634e+11Hz 0.286883 -0.939281
+ 1.635e+11Hz 0.286145 -0.939484
+ 1.636e+11Hz 0.285407 -0.939687
+ 1.637e+11Hz 0.284669 -0.939888
+ 1.638e+11Hz 0.283931 -0.940089
+ 1.639e+11Hz 0.283193 -0.940289
+ 1.64e+11Hz 0.282455 -0.940489
+ 1.641e+11Hz 0.281716 -0.940688
+ 1.642e+11Hz 0.280977 -0.940886
+ 1.643e+11Hz 0.280239 -0.941084
+ 1.644e+11Hz 0.2795 -0.941281
+ 1.645e+11Hz 0.278761 -0.941477
+ 1.646e+11Hz 0.278022 -0.941672
+ 1.647e+11Hz 0.277283 -0.941867
+ 1.648e+11Hz 0.276544 -0.942061
+ 1.649e+11Hz 0.275805 -0.942255
+ 1.65e+11Hz 0.275066 -0.942447
+ 1.651e+11Hz 0.274327 -0.94264
+ 1.652e+11Hz 0.273587 -0.942831
+ 1.653e+11Hz 0.272848 -0.943022
+ 1.654e+11Hz 0.272108 -0.943212
+ 1.655e+11Hz 0.271369 -0.943401
+ 1.656e+11Hz 0.270629 -0.94359
+ 1.657e+11Hz 0.269889 -0.943778
+ 1.658e+11Hz 0.26915 -0.943965
+ 1.659e+11Hz 0.26841 -0.944152
+ 1.66e+11Hz 0.26767 -0.944338
+ 1.661e+11Hz 0.26693 -0.944523
+ 1.662e+11Hz 0.26619 -0.944708
+ 1.663e+11Hz 0.26545 -0.944892
+ 1.664e+11Hz 0.26471 -0.945075
+ 1.665e+11Hz 0.26397 -0.945258
+ 1.666e+11Hz 0.26323 -0.94544
+ 1.667e+11Hz 0.26249 -0.945621
+ 1.668e+11Hz 0.26175 -0.945802
+ 1.669e+11Hz 0.26101 -0.945982
+ 1.67e+11Hz 0.26027 -0.946161
+ 1.671e+11Hz 0.259529 -0.946339
+ 1.672e+11Hz 0.258789 -0.946517
+ 1.673e+11Hz 0.258049 -0.946695
+ 1.674e+11Hz 0.257309 -0.946871
+ 1.675e+11Hz 0.256568 -0.947047
+ 1.676e+11Hz 0.255828 -0.947223
+ 1.677e+11Hz 0.255088 -0.947397
+ 1.678e+11Hz 0.254348 -0.947571
+ 1.679e+11Hz 0.253607 -0.947744
+ 1.68e+11Hz 0.252867 -0.947917
+ 1.681e+11Hz 0.252127 -0.948089
+ 1.682e+11Hz 0.251386 -0.94826
+ 1.683e+11Hz 0.250646 -0.948431
+ 1.684e+11Hz 0.249906 -0.948601
+ 1.685e+11Hz 0.249165 -0.948771
+ 1.686e+11Hz 0.248425 -0.948939
+ 1.687e+11Hz 0.247685 -0.949108
+ 1.688e+11Hz 0.246944 -0.949275
+ 1.689e+11Hz 0.246204 -0.949442
+ 1.69e+11Hz 0.245464 -0.949608
+ 1.691e+11Hz 0.244724 -0.949774
+ 1.692e+11Hz 0.243983 -0.949939
+ 1.693e+11Hz 0.243243 -0.950103
+ 1.694e+11Hz 0.242503 -0.950266
+ 1.695e+11Hz 0.241763 -0.950429
+ 1.696e+11Hz 0.241023 -0.950592
+ 1.697e+11Hz 0.240283 -0.950754
+ 1.698e+11Hz 0.239543 -0.950915
+ 1.699e+11Hz 0.238803 -0.951075
+ 1.7e+11Hz 0.238063 -0.951235
+ 1.701e+11Hz 0.237323 -0.951394
+ 1.702e+11Hz 0.236583 -0.951553
+ 1.703e+11Hz 0.235843 -0.951711
+ 1.704e+11Hz 0.235103 -0.951869
+ 1.705e+11Hz 0.234363 -0.952025
+ 1.706e+11Hz 0.233623 -0.952182
+ 1.707e+11Hz 0.232884 -0.952337
+ 1.708e+11Hz 0.232144 -0.952492
+ 1.709e+11Hz 0.231404 -0.952647
+ 1.71e+11Hz 0.230665 -0.952801
+ 1.711e+11Hz 0.229925 -0.952954
+ 1.712e+11Hz 0.229185 -0.953106
+ 1.713e+11Hz 0.228446 -0.953258
+ 1.714e+11Hz 0.227706 -0.95341
+ 1.715e+11Hz 0.226967 -0.953561
+ 1.716e+11Hz 0.226228 -0.953711
+ 1.717e+11Hz 0.225488 -0.953861
+ 1.718e+11Hz 0.224749 -0.95401
+ 1.719e+11Hz 0.22401 -0.954158
+ 1.72e+11Hz 0.223271 -0.954306
+ 1.721e+11Hz 0.222532 -0.954453
+ 1.722e+11Hz 0.221793 -0.9546
+ 1.723e+11Hz 0.221054 -0.954747
+ 1.724e+11Hz 0.220315 -0.954892
+ 1.725e+11Hz 0.219576 -0.955037
+ 1.726e+11Hz 0.218837 -0.955182
+ 1.727e+11Hz 0.218098 -0.955326
+ 1.728e+11Hz 0.21736 -0.955469
+ 1.729e+11Hz 0.216621 -0.955612
+ 1.73e+11Hz 0.215882 -0.955754
+ 1.731e+11Hz 0.215144 -0.955896
+ 1.732e+11Hz 0.214405 -0.956037
+ 1.733e+11Hz 0.213667 -0.956178
+ 1.734e+11Hz 0.212929 -0.956318
+ 1.735e+11Hz 0.21219 -0.956458
+ 1.736e+11Hz 0.211452 -0.956597
+ 1.737e+11Hz 0.210714 -0.956735
+ 1.738e+11Hz 0.209976 -0.956873
+ 1.739e+11Hz 0.209237 -0.95701
+ 1.74e+11Hz 0.208499 -0.957147
+ 1.741e+11Hz 0.207761 -0.957284
+ 1.742e+11Hz 0.207023 -0.957419
+ 1.743e+11Hz 0.206286 -0.957555
+ 1.744e+11Hz 0.205548 -0.957689
+ 1.745e+11Hz 0.20481 -0.957824
+ 1.746e+11Hz 0.204072 -0.957957
+ 1.747e+11Hz 0.203335 -0.958091
+ 1.748e+11Hz 0.202597 -0.958223
+ 1.749e+11Hz 0.201859 -0.958356
+ 1.75e+11Hz 0.201122 -0.958487
+ 1.751e+11Hz 0.200384 -0.958618
+ 1.752e+11Hz 0.199647 -0.958749
+ 1.753e+11Hz 0.19891 -0.958879
+ 1.754e+11Hz 0.198172 -0.959009
+ 1.755e+11Hz 0.197435 -0.959138
+ 1.756e+11Hz 0.196698 -0.959267
+ 1.757e+11Hz 0.195961 -0.959395
+ 1.758e+11Hz 0.195223 -0.959523
+ 1.759e+11Hz 0.194486 -0.95965
+ 1.76e+11Hz 0.193749 -0.959776
+ 1.761e+11Hz 0.193012 -0.959903
+ 1.762e+11Hz 0.192275 -0.960028
+ 1.763e+11Hz 0.191538 -0.960154
+ 1.764e+11Hz 0.190801 -0.960278
+ 1.765e+11Hz 0.190064 -0.960402
+ 1.766e+11Hz 0.189328 -0.960526
+ 1.767e+11Hz 0.188591 -0.96065
+ 1.768e+11Hz 0.187854 -0.960772
+ 1.769e+11Hz 0.187117 -0.960895
+ 1.77e+11Hz 0.186381 -0.961017
+ 1.771e+11Hz 0.185644 -0.961138
+ 1.772e+11Hz 0.184907 -0.961259
+ 1.773e+11Hz 0.184171 -0.961379
+ 1.774e+11Hz 0.183434 -0.961499
+ 1.775e+11Hz 0.182697 -0.961619
+ 1.776e+11Hz 0.181961 -0.961738
+ 1.777e+11Hz 0.181224 -0.961856
+ 1.778e+11Hz 0.180488 -0.961974
+ 1.779e+11Hz 0.179751 -0.962092
+ 1.78e+11Hz 0.179015 -0.962209
+ 1.781e+11Hz 0.178278 -0.962326
+ 1.782e+11Hz 0.177542 -0.962442
+ 1.783e+11Hz 0.176805 -0.962558
+ 1.784e+11Hz 0.176069 -0.962673
+ 1.785e+11Hz 0.175333 -0.962788
+ 1.786e+11Hz 0.174596 -0.962902
+ 1.787e+11Hz 0.17386 -0.963016
+ 1.788e+11Hz 0.173123 -0.96313
+ 1.789e+11Hz 0.172387 -0.963243
+ 1.79e+11Hz 0.171651 -0.963355
+ 1.791e+11Hz 0.170914 -0.963468
+ 1.792e+11Hz 0.170178 -0.963579
+ 1.793e+11Hz 0.169441 -0.96369
+ 1.794e+11Hz 0.168705 -0.963801
+ 1.795e+11Hz 0.167968 -0.963911
+ 1.796e+11Hz 0.167232 -0.964021
+ 1.797e+11Hz 0.166496 -0.964131
+ 1.798e+11Hz 0.165759 -0.96424
+ 1.799e+11Hz 0.165023 -0.964348
+ 1.8e+11Hz 0.164286 -0.964456
+ 1.801e+11Hz 0.16355 -0.964564
+ 1.802e+11Hz 0.162813 -0.964671
+ 1.803e+11Hz 0.162077 -0.964778
+ 1.804e+11Hz 0.16134 -0.964884
+ 1.805e+11Hz 0.160604 -0.96499
+ 1.806e+11Hz 0.159867 -0.965095
+ 1.807e+11Hz 0.15913 -0.9652
+ 1.808e+11Hz 0.158394 -0.965304
+ 1.809e+11Hz 0.157657 -0.965408
+ 1.81e+11Hz 0.15692 -0.965512
+ 1.811e+11Hz 0.156184 -0.965615
+ 1.812e+11Hz 0.155447 -0.965718
+ 1.813e+11Hz 0.15471 -0.96582
+ 1.814e+11Hz 0.153973 -0.965921
+ 1.815e+11Hz 0.153236 -0.966023
+ 1.816e+11Hz 0.152499 -0.966124
+ 1.817e+11Hz 0.151762 -0.966224
+ 1.818e+11Hz 0.151025 -0.966324
+ 1.819e+11Hz 0.150288 -0.966423
+ 1.82e+11Hz 0.149551 -0.966522
+ 1.821e+11Hz 0.148814 -0.966621
+ 1.822e+11Hz 0.148077 -0.966719
+ 1.823e+11Hz 0.14734 -0.966817
+ 1.824e+11Hz 0.146602 -0.966914
+ 1.825e+11Hz 0.145865 -0.967011
+ 1.826e+11Hz 0.145128 -0.967107
+ 1.827e+11Hz 0.14439 -0.967203
+ 1.828e+11Hz 0.143653 -0.967298
+ 1.829e+11Hz 0.142915 -0.967393
+ 1.83e+11Hz 0.142178 -0.967488
+ 1.831e+11Hz 0.14144 -0.967582
+ 1.832e+11Hz 0.140702 -0.967675
+ 1.833e+11Hz 0.139965 -0.967768
+ 1.834e+11Hz 0.139227 -0.967861
+ 1.835e+11Hz 0.138489 -0.967953
+ 1.836e+11Hz 0.137751 -0.968045
+ 1.837e+11Hz 0.137013 -0.968136
+ 1.838e+11Hz 0.136275 -0.968227
+ 1.839e+11Hz 0.135537 -0.968317
+ 1.84e+11Hz 0.134799 -0.968407
+ 1.841e+11Hz 0.13406 -0.968496
+ 1.842e+11Hz 0.133322 -0.968585
+ 1.843e+11Hz 0.132584 -0.968673
+ 1.844e+11Hz 0.131845 -0.968761
+ 1.845e+11Hz 0.131107 -0.968849
+ 1.846e+11Hz 0.130368 -0.968936
+ 1.847e+11Hz 0.129629 -0.969022
+ 1.848e+11Hz 0.128891 -0.969109
+ 1.849e+11Hz 0.128152 -0.969194
+ 1.85e+11Hz 0.127413 -0.969279
+ 1.851e+11Hz 0.126674 -0.969364
+ 1.852e+11Hz 0.125935 -0.969448
+ 1.853e+11Hz 0.125196 -0.969532
+ 1.854e+11Hz 0.124457 -0.969615
+ 1.855e+11Hz 0.123717 -0.969698
+ 1.856e+11Hz 0.122978 -0.96978
+ 1.857e+11Hz 0.122239 -0.969862
+ 1.858e+11Hz 0.121499 -0.969943
+ 1.859e+11Hz 0.120759 -0.970024
+ 1.86e+11Hz 0.12002 -0.970104
+ 1.861e+11Hz 0.11928 -0.970184
+ 1.862e+11Hz 0.11854 -0.970263
+ 1.863e+11Hz 0.1178 -0.970342
+ 1.864e+11Hz 0.11706 -0.97042
+ 1.865e+11Hz 0.11632 -0.970498
+ 1.866e+11Hz 0.11558 -0.970576
+ 1.867e+11Hz 0.11484 -0.970652
+ 1.868e+11Hz 0.1141 -0.970729
+ 1.869e+11Hz 0.113359 -0.970805
+ 1.87e+11Hz 0.112619 -0.97088
+ 1.871e+11Hz 0.111878 -0.970955
+ 1.872e+11Hz 0.111138 -0.971029
+ 1.873e+11Hz 0.110397 -0.971103
+ 1.874e+11Hz 0.109656 -0.971177
+ 1.875e+11Hz 0.108915 -0.971249
+ 1.876e+11Hz 0.108175 -0.971322
+ 1.877e+11Hz 0.107434 -0.971394
+ 1.878e+11Hz 0.106692 -0.971465
+ 1.879e+11Hz 0.105951 -0.971536
+ 1.88e+11Hz 0.10521 -0.971606
+ 1.881e+11Hz 0.104469 -0.971676
+ 1.882e+11Hz 0.103727 -0.971745
+ 1.883e+11Hz 0.102986 -0.971814
+ 1.884e+11Hz 0.102244 -0.971883
+ 1.885e+11Hz 0.101503 -0.97195
+ 1.886e+11Hz 0.100761 -0.972018
+ 1.887e+11Hz 0.100019 -0.972084
+ 1.888e+11Hz 0.0992772 -0.972151
+ 1.889e+11Hz 0.0985352 -0.972216
+ 1.89e+11Hz 0.0977932 -0.972282
+ 1.891e+11Hz 0.0970511 -0.972346
+ 1.892e+11Hz 0.0963089 -0.972411
+ 1.893e+11Hz 0.0955666 -0.972474
+ 1.894e+11Hz 0.0948242 -0.972537
+ 1.895e+11Hz 0.0940818 -0.9726
+ 1.896e+11Hz 0.0933393 -0.972662
+ 1.897e+11Hz 0.0925967 -0.972724
+ 1.898e+11Hz 0.0918541 -0.972785
+ 1.899e+11Hz 0.0911114 -0.972845
+ 1.9e+11Hz 0.0903686 -0.972905
+ 1.901e+11Hz 0.0896257 -0.972965
+ 1.902e+11Hz 0.0888827 -0.973024
+ 1.903e+11Hz 0.0881397 -0.973082
+ 1.904e+11Hz 0.0873966 -0.97314
+ 1.905e+11Hz 0.0866534 -0.973198
+ 1.906e+11Hz 0.0859102 -0.973254
+ 1.907e+11Hz 0.0851669 -0.973311
+ 1.908e+11Hz 0.0844235 -0.973367
+ 1.909e+11Hz 0.08368 -0.973422
+ 1.91e+11Hz 0.0829365 -0.973477
+ 1.911e+11Hz 0.0821929 -0.973531
+ 1.912e+11Hz 0.0814492 -0.973584
+ 1.913e+11Hz 0.0807055 -0.973638
+ 1.914e+11Hz 0.0799617 -0.97369
+ 1.915e+11Hz 0.0792178 -0.973742
+ 1.916e+11Hz 0.0784739 -0.973794
+ 1.917e+11Hz 0.0777299 -0.973845
+ 1.918e+11Hz 0.0769858 -0.973895
+ 1.919e+11Hz 0.0762416 -0.973945
+ 1.92e+11Hz 0.0754974 -0.973995
+ 1.921e+11Hz 0.0747532 -0.974043
+ 1.922e+11Hz 0.0740088 -0.974092
+ 1.923e+11Hz 0.0732644 -0.97414
+ 1.924e+11Hz 0.0725199 -0.974187
+ 1.925e+11Hz 0.0717754 -0.974233
+ 1.926e+11Hz 0.0710308 -0.97428
+ 1.927e+11Hz 0.0702861 -0.974325
+ 1.928e+11Hz 0.0695414 -0.97437
+ 1.929e+11Hz 0.0687966 -0.974415
+ 1.93e+11Hz 0.0680518 -0.974459
+ 1.931e+11Hz 0.0673068 -0.974502
+ 1.932e+11Hz 0.0665619 -0.974545
+ 1.933e+11Hz 0.0658168 -0.974588
+ 1.934e+11Hz 0.0650717 -0.974629
+ 1.935e+11Hz 0.0643266 -0.974671
+ 1.936e+11Hz 0.0635814 -0.974711
+ 1.937e+11Hz 0.0628361 -0.974752
+ 1.938e+11Hz 0.0620907 -0.974791
+ 1.939e+11Hz 0.0613453 -0.97483
+ 1.94e+11Hz 0.0605999 -0.974869
+ 1.941e+11Hz 0.0598544 -0.974907
+ 1.942e+11Hz 0.0591088 -0.974944
+ 1.943e+11Hz 0.0583632 -0.974981
+ 1.944e+11Hz 0.0576175 -0.975018
+ 1.945e+11Hz 0.0568717 -0.975054
+ 1.946e+11Hz 0.0561259 -0.975089
+ 1.947e+11Hz 0.0553801 -0.975123
+ 1.948e+11Hz 0.0546342 -0.975158
+ 1.949e+11Hz 0.0538882 -0.975191
+ 1.95e+11Hz 0.0531422 -0.975224
+ 1.951e+11Hz 0.0523961 -0.975257
+ 1.952e+11Hz 0.05165 -0.975289
+ 1.953e+11Hz 0.0509038 -0.97532
+ 1.954e+11Hz 0.0501575 -0.975351
+ 1.955e+11Hz 0.0494112 -0.975381
+ 1.956e+11Hz 0.0486649 -0.975411
+ 1.957e+11Hz 0.0479185 -0.97544
+ 1.958e+11Hz 0.047172 -0.975469
+ 1.959e+11Hz 0.0464255 -0.975497
+ 1.96e+11Hz 0.045679 -0.975525
+ 1.961e+11Hz 0.0449323 -0.975552
+ 1.962e+11Hz 0.0441857 -0.975578
+ 1.963e+11Hz 0.043439 -0.975604
+ 1.964e+11Hz 0.0426922 -0.975629
+ 1.965e+11Hz 0.0419454 -0.975654
+ 1.966e+11Hz 0.0411985 -0.975678
+ 1.967e+11Hz 0.0404515 -0.975702
+ 1.968e+11Hz 0.0397046 -0.975725
+ 1.969e+11Hz 0.0389575 -0.975748
+ 1.97e+11Hz 0.0382104 -0.97577
+ 1.971e+11Hz 0.0374633 -0.975791
+ 1.972e+11Hz 0.0367161 -0.975812
+ 1.973e+11Hz 0.0359689 -0.975832
+ 1.974e+11Hz 0.0352216 -0.975852
+ 1.975e+11Hz 0.0344743 -0.975871
+ 1.976e+11Hz 0.0337269 -0.97589
+ 1.977e+11Hz 0.0329794 -0.975908
+ 1.978e+11Hz 0.032232 -0.975925
+ 1.979e+11Hz 0.0314844 -0.975942
+ 1.98e+11Hz 0.0307368 -0.975958
+ 1.981e+11Hz 0.0299892 -0.975974
+ 1.982e+11Hz 0.0292415 -0.975989
+ 1.983e+11Hz 0.0284938 -0.976004
+ 1.984e+11Hz 0.027746 -0.976018
+ 1.985e+11Hz 0.0269982 -0.976031
+ 1.986e+11Hz 0.0262503 -0.976044
+ 1.987e+11Hz 0.0255024 -0.976057
+ 1.988e+11Hz 0.0247544 -0.976068
+ 1.989e+11Hz 0.0240064 -0.97608
+ 1.99e+11Hz 0.0232584 -0.97609
+ 1.991e+11Hz 0.0225103 -0.9761
+ 1.992e+11Hz 0.0217621 -0.97611
+ 1.993e+11Hz 0.0210139 -0.976119
+ 1.994e+11Hz 0.0202657 -0.976127
+ 1.995e+11Hz 0.0195174 -0.976135
+ 1.996e+11Hz 0.018769 -0.976142
+ 1.997e+11Hz 0.0180206 -0.976148
+ 1.998e+11Hz 0.0172722 -0.976154
+ 1.999e+11Hz 0.0165238 -0.97616
+ 2e+11Hz 0.0157752 -0.976165
+ 2.001e+11Hz 0.0150267 -0.976169
+ 2.002e+11Hz 0.0142781 -0.976173
+ 2.003e+11Hz 0.0135295 -0.976176
+ 2.004e+11Hz 0.0127808 -0.976178
+ 2.005e+11Hz 0.0120321 -0.97618
+ 2.006e+11Hz 0.0112833 -0.976181
+ 2.007e+11Hz 0.0105345 -0.976182
+ 2.008e+11Hz 0.00978566 -0.976182
+ 2.009e+11Hz 0.00903679 -0.976182
+ 2.01e+11Hz 0.00828787 -0.976181
+ 2.011e+11Hz 0.00753892 -0.976179
+ 2.012e+11Hz 0.00678993 -0.976177
+ 2.013e+11Hz 0.00604091 -0.976174
+ 2.014e+11Hz 0.00529185 -0.97617
+ 2.015e+11Hz 0.00454275 -0.976166
+ 2.016e+11Hz 0.00379363 -0.976162
+ 2.017e+11Hz 0.00304447 -0.976156
+ 2.018e+11Hz 0.00229528 -0.97615
+ 2.019e+11Hz 0.00154605 -0.976144
+ 2.02e+11Hz 0.000796802 -0.976137
+ 2.021e+11Hz 4.7521e-05 -0.976129
+ 2.022e+11Hz -0.000701788 -0.976121
+ 2.023e+11Hz -0.00145112 -0.976112
+ 2.024e+11Hz -0.00220049 -0.976102
+ 2.025e+11Hz -0.00294987 -0.976092
+ 2.026e+11Hz -0.00369929 -0.976081
+ 2.027e+11Hz -0.00444872 -0.97607
+ 2.028e+11Hz -0.00519818 -0.976058
+ 2.029e+11Hz -0.00594765 -0.976045
+ 2.03e+11Hz -0.00669715 -0.976032
+ 2.031e+11Hz -0.00744666 -0.976018
+ 2.032e+11Hz -0.00819619 -0.976004
+ 2.033e+11Hz -0.00894573 -0.975988
+ 2.034e+11Hz -0.00969529 -0.975973
+ 2.035e+11Hz -0.0104449 -0.975956
+ 2.036e+11Hz -0.0111944 -0.975939
+ 2.037e+11Hz -0.011944 -0.975922
+ 2.038e+11Hz -0.0126936 -0.975903
+ 2.039e+11Hz -0.0134432 -0.975884
+ 2.04e+11Hz -0.0141928 -0.975865
+ 2.041e+11Hz -0.0149425 -0.975845
+ 2.042e+11Hz -0.0156921 -0.975824
+ 2.043e+11Hz -0.0164417 -0.975802
+ 2.044e+11Hz -0.0171913 -0.97578
+ 2.045e+11Hz -0.0179409 -0.975758
+ 2.046e+11Hz -0.0186905 -0.975734
+ 2.047e+11Hz -0.0194401 -0.97571
+ 2.048e+11Hz -0.0201897 -0.975686
+ 2.049e+11Hz -0.0209393 -0.97566
+ 2.05e+11Hz -0.0216888 -0.975634
+ 2.051e+11Hz -0.0224384 -0.975608
+ 2.052e+11Hz -0.0231879 -0.975581
+ 2.053e+11Hz -0.0239374 -0.975553
+ 2.054e+11Hz -0.0246869 -0.975524
+ 2.055e+11Hz -0.0254363 -0.975495
+ 2.056e+11Hz -0.0261858 -0.975465
+ 2.057e+11Hz -0.0269352 -0.975435
+ 2.058e+11Hz -0.0276845 -0.975403
+ 2.059e+11Hz -0.0284339 -0.975372
+ 2.06e+11Hz -0.0291832 -0.975339
+ 2.061e+11Hz -0.0299325 -0.975306
+ 2.062e+11Hz -0.0306817 -0.975272
+ 2.063e+11Hz -0.0314309 -0.975238
+ 2.064e+11Hz -0.03218 -0.975203
+ 2.065e+11Hz -0.0329291 -0.975167
+ 2.066e+11Hz -0.0336781 -0.975131
+ 2.067e+11Hz -0.0344271 -0.975094
+ 2.068e+11Hz -0.035176 -0.975056
+ 2.069e+11Hz -0.0359249 -0.975017
+ 2.07e+11Hz -0.0366737 -0.974978
+ 2.071e+11Hz -0.0374225 -0.974939
+ 2.072e+11Hz -0.0381711 -0.974898
+ 2.073e+11Hz -0.0389197 -0.974857
+ 2.074e+11Hz -0.0396683 -0.974816
+ 2.075e+11Hz -0.0404167 -0.974773
+ 2.076e+11Hz -0.0411651 -0.97473
+ 2.077e+11Hz -0.0419134 -0.974686
+ 2.078e+11Hz -0.0426616 -0.974642
+ 2.079e+11Hz -0.0434098 -0.974597
+ 2.08e+11Hz -0.0441578 -0.974551
+ 2.081e+11Hz -0.0449058 -0.974505
+ 2.082e+11Hz -0.0456536 -0.974458
+ 2.083e+11Hz -0.0464014 -0.97441
+ 2.084e+11Hz -0.047149 -0.974362
+ 2.085e+11Hz -0.0478966 -0.974313
+ 2.086e+11Hz -0.048644 -0.974263
+ 2.087e+11Hz -0.0493913 -0.974213
+ 2.088e+11Hz -0.0501385 -0.974162
+ 2.089e+11Hz -0.0508856 -0.974111
+ 2.09e+11Hz -0.0516326 -0.974058
+ 2.091e+11Hz -0.0523794 -0.974005
+ 2.092e+11Hz -0.0531262 -0.973952
+ 2.093e+11Hz -0.0538728 -0.973897
+ 2.094e+11Hz -0.0546192 -0.973843
+ 2.095e+11Hz -0.0553656 -0.973787
+ 2.096e+11Hz -0.0561117 -0.973731
+ 2.097e+11Hz -0.0568578 -0.973674
+ 2.098e+11Hz -0.0576037 -0.973616
+ 2.099e+11Hz -0.0583494 -0.973558
+ 2.1e+11Hz -0.059095 -0.973499
+ 2.101e+11Hz -0.0598405 -0.97344
+ 2.102e+11Hz -0.0605858 -0.97338
+ 2.103e+11Hz -0.0613309 -0.973319
+ 2.104e+11Hz -0.0620758 -0.973257
+ 2.105e+11Hz -0.0628206 -0.973195
+ 2.106e+11Hz -0.0635652 -0.973133
+ 2.107e+11Hz -0.0643097 -0.973069
+ 2.108e+11Hz -0.065054 -0.973005
+ 2.109e+11Hz -0.0657981 -0.972941
+ 2.11e+11Hz -0.066542 -0.972875
+ 2.111e+11Hz -0.0672857 -0.97281
+ 2.112e+11Hz -0.0680292 -0.972743
+ 2.113e+11Hz -0.0687726 -0.972676
+ 2.114e+11Hz -0.0695157 -0.972608
+ 2.115e+11Hz -0.0702587 -0.97254
+ 2.116e+11Hz -0.0710014 -0.972471
+ 2.117e+11Hz -0.071744 -0.972401
+ 2.118e+11Hz -0.0724863 -0.972331
+ 2.119e+11Hz -0.0732284 -0.97226
+ 2.12e+11Hz -0.0739704 -0.972189
+ 2.121e+11Hz -0.0747121 -0.972116
+ 2.122e+11Hz -0.0754535 -0.972044
+ 2.123e+11Hz -0.0761948 -0.97197
+ 2.124e+11Hz -0.0769359 -0.971897
+ 2.125e+11Hz -0.0776767 -0.971822
+ 2.126e+11Hz -0.0784173 -0.971747
+ 2.127e+11Hz -0.0791577 -0.971671
+ 2.128e+11Hz -0.0798978 -0.971595
+ 2.129e+11Hz -0.0806377 -0.971518
+ 2.13e+11Hz -0.0813774 -0.971441
+ 2.131e+11Hz -0.0821168 -0.971363
+ 2.132e+11Hz -0.082856 -0.971284
+ 2.133e+11Hz -0.0835949 -0.971205
+ 2.134e+11Hz -0.0843336 -0.971125
+ 2.135e+11Hz -0.0850721 -0.971045
+ 2.136e+11Hz -0.0858103 -0.970964
+ 2.137e+11Hz -0.0865482 -0.970883
+ 2.138e+11Hz -0.0872859 -0.970801
+ 2.139e+11Hz -0.0880233 -0.970718
+ 2.14e+11Hz -0.0887605 -0.970635
+ 2.141e+11Hz -0.0894975 -0.970552
+ 2.142e+11Hz -0.0902341 -0.970468
+ 2.143e+11Hz -0.0909705 -0.970383
+ 2.144e+11Hz -0.0917067 -0.970298
+ 2.145e+11Hz -0.0924426 -0.970212
+ 2.146e+11Hz -0.0931782 -0.970126
+ 2.147e+11Hz -0.0939135 -0.970039
+ 2.148e+11Hz -0.0946486 -0.969952
+ 2.149e+11Hz -0.0953834 -0.969864
+ 2.15e+11Hz -0.096118 -0.969776
+ 2.151e+11Hz -0.0968523 -0.969687
+ 2.152e+11Hz -0.0975863 -0.969597
+ 2.153e+11Hz -0.09832 -0.969508
+ 2.154e+11Hz -0.0990535 -0.969417
+ 2.155e+11Hz -0.0997867 -0.969327
+ 2.156e+11Hz -0.10052 -0.969235
+ 2.157e+11Hz -0.101252 -0.969144
+ 2.158e+11Hz -0.101985 -0.969051
+ 2.159e+11Hz -0.102717 -0.968959
+ 2.16e+11Hz -0.103449 -0.968866
+ 2.161e+11Hz -0.10418 -0.968772
+ 2.162e+11Hz -0.104911 -0.968678
+ 2.163e+11Hz -0.105642 -0.968583
+ 2.164e+11Hz -0.106373 -0.968488
+ 2.165e+11Hz -0.107104 -0.968393
+ 2.166e+11Hz -0.107834 -0.968297
+ 2.167e+11Hz -0.108564 -0.968201
+ 2.168e+11Hz -0.109293 -0.968104
+ 2.169e+11Hz -0.110023 -0.968007
+ 2.17e+11Hz -0.110752 -0.96791
+ 2.171e+11Hz -0.111481 -0.967812
+ 2.172e+11Hz -0.112209 -0.967713
+ 2.173e+11Hz -0.112937 -0.967615
+ 2.174e+11Hz -0.113666 -0.967515
+ 2.175e+11Hz -0.114393 -0.967416
+ 2.176e+11Hz -0.115121 -0.967316
+ 2.177e+11Hz -0.115848 -0.967216
+ 2.178e+11Hz -0.116575 -0.967115
+ 2.179e+11Hz -0.117302 -0.967014
+ 2.18e+11Hz -0.118028 -0.966912
+ 2.181e+11Hz -0.118754 -0.96681
+ 2.182e+11Hz -0.11948 -0.966708
+ 2.183e+11Hz -0.120206 -0.966606
+ 2.184e+11Hz -0.120932 -0.966503
+ 2.185e+11Hz -0.121657 -0.966399
+ 2.186e+11Hz -0.122382 -0.966296
+ 2.187e+11Hz -0.123106 -0.966192
+ 2.188e+11Hz -0.123831 -0.966087
+ 2.189e+11Hz -0.124555 -0.965983
+ 2.19e+11Hz -0.125279 -0.965878
+ 2.191e+11Hz -0.126003 -0.965772
+ 2.192e+11Hz -0.126727 -0.965667
+ 2.193e+11Hz -0.12745 -0.965561
+ 2.194e+11Hz -0.128173 -0.965454
+ 2.195e+11Hz -0.128896 -0.965348
+ 2.196e+11Hz -0.129619 -0.965241
+ 2.197e+11Hz -0.130341 -0.965134
+ 2.198e+11Hz -0.131063 -0.965026
+ 2.199e+11Hz -0.131786 -0.964918
+ 2.2e+11Hz -0.132507 -0.96481
+ 2.201e+11Hz -0.133229 -0.964702
+ 2.202e+11Hz -0.133951 -0.964593
+ 2.203e+11Hz -0.134672 -0.964484
+ 2.204e+11Hz -0.135393 -0.964375
+ 2.205e+11Hz -0.136114 -0.964265
+ 2.206e+11Hz -0.136835 -0.964155
+ 2.207e+11Hz -0.137555 -0.964045
+ 2.208e+11Hz -0.138275 -0.963935
+ 2.209e+11Hz -0.138996 -0.963824
+ 2.21e+11Hz -0.139716 -0.963713
+ 2.211e+11Hz -0.140436 -0.963602
+ 2.212e+11Hz -0.141155 -0.963491
+ 2.213e+11Hz -0.141875 -0.963379
+ 2.214e+11Hz -0.142594 -0.963267
+ 2.215e+11Hz -0.143314 -0.963155
+ 2.216e+11Hz -0.144033 -0.963042
+ 2.217e+11Hz -0.144752 -0.96293
+ 2.218e+11Hz -0.145471 -0.962817
+ 2.219e+11Hz -0.14619 -0.962703
+ 2.22e+11Hz -0.146908 -0.96259
+ 2.221e+11Hz -0.147627 -0.962476
+ 2.222e+11Hz -0.148346 -0.962362
+ 2.223e+11Hz -0.149064 -0.962248
+ 2.224e+11Hz -0.149782 -0.962134
+ 2.225e+11Hz -0.1505 -0.962019
+ 2.226e+11Hz -0.151219 -0.961904
+ 2.227e+11Hz -0.151937 -0.961789
+ 2.228e+11Hz -0.152655 -0.961673
+ 2.229e+11Hz -0.153372 -0.961558
+ 2.23e+11Hz -0.15409 -0.961442
+ 2.231e+11Hz -0.154808 -0.961326
+ 2.232e+11Hz -0.155526 -0.96121
+ 2.233e+11Hz -0.156243 -0.961093
+ 2.234e+11Hz -0.156961 -0.960976
+ 2.235e+11Hz -0.157679 -0.960859
+ 2.236e+11Hz -0.158396 -0.960742
+ 2.237e+11Hz -0.159114 -0.960625
+ 2.238e+11Hz -0.159831 -0.960507
+ 2.239e+11Hz -0.160549 -0.960389
+ 2.24e+11Hz -0.161266 -0.960271
+ 2.241e+11Hz -0.161984 -0.960152
+ 2.242e+11Hz -0.162701 -0.960034
+ 2.243e+11Hz -0.163419 -0.959915
+ 2.244e+11Hz -0.164136 -0.959796
+ 2.245e+11Hz -0.164854 -0.959677
+ 2.246e+11Hz -0.165571 -0.959557
+ 2.247e+11Hz -0.166289 -0.959437
+ 2.248e+11Hz -0.167006 -0.959317
+ 2.249e+11Hz -0.167724 -0.959197
+ 2.25e+11Hz -0.168442 -0.959076
+ 2.251e+11Hz -0.169159 -0.958955
+ 2.252e+11Hz -0.169877 -0.958834
+ 2.253e+11Hz -0.170595 -0.958713
+ 2.254e+11Hz -0.171313 -0.958592
+ 2.255e+11Hz -0.172031 -0.95847
+ 2.256e+11Hz -0.172749 -0.958348
+ 2.257e+11Hz -0.173467 -0.958225
+ 2.258e+11Hz -0.174185 -0.958103
+ 2.259e+11Hz -0.174904 -0.95798
+ 2.26e+11Hz -0.175622 -0.957857
+ 2.261e+11Hz -0.176341 -0.957734
+ 2.262e+11Hz -0.177059 -0.95761
+ 2.263e+11Hz -0.177778 -0.957486
+ 2.264e+11Hz -0.178497 -0.957362
+ 2.265e+11Hz -0.179216 -0.957238
+ 2.266e+11Hz -0.179935 -0.957113
+ 2.267e+11Hz -0.180654 -0.956988
+ 2.268e+11Hz -0.181374 -0.956862
+ 2.269e+11Hz -0.182093 -0.956737
+ 2.27e+11Hz -0.182813 -0.956611
+ 2.271e+11Hz -0.183533 -0.956485
+ 2.272e+11Hz -0.184252 -0.956358
+ 2.273e+11Hz -0.184973 -0.956231
+ 2.274e+11Hz -0.185693 -0.956104
+ 2.275e+11Hz -0.186413 -0.955977
+ 2.276e+11Hz -0.187134 -0.955849
+ 2.277e+11Hz -0.187855 -0.955721
+ 2.278e+11Hz -0.188576 -0.955592
+ 2.279e+11Hz -0.189297 -0.955464
+ 2.28e+11Hz -0.190018 -0.955335
+ 2.281e+11Hz -0.19074 -0.955205
+ 2.282e+11Hz -0.191461 -0.955075
+ 2.283e+11Hz -0.192183 -0.954945
+ 2.284e+11Hz -0.192905 -0.954815
+ 2.285e+11Hz -0.193627 -0.954684
+ 2.286e+11Hz -0.19435 -0.954552
+ 2.287e+11Hz -0.195073 -0.954421
+ 2.288e+11Hz -0.195796 -0.954289
+ 2.289e+11Hz -0.196519 -0.954156
+ 2.29e+11Hz -0.197242 -0.954023
+ 2.291e+11Hz -0.197965 -0.95389
+ 2.292e+11Hz -0.198689 -0.953757
+ 2.293e+11Hz -0.199413 -0.953623
+ 2.294e+11Hz -0.200137 -0.953488
+ 2.295e+11Hz -0.200862 -0.953353
+ 2.296e+11Hz -0.201587 -0.953218
+ 2.297e+11Hz -0.202311 -0.953082
+ 2.298e+11Hz -0.203037 -0.952946
+ 2.299e+11Hz -0.203762 -0.95281
+ 2.3e+11Hz -0.204487 -0.952673
+ 2.301e+11Hz -0.205213 -0.952535
+ 2.302e+11Hz -0.205939 -0.952397
+ 2.303e+11Hz -0.206666 -0.952259
+ 2.304e+11Hz -0.207392 -0.95212
+ 2.305e+11Hz -0.208119 -0.95198
+ 2.306e+11Hz -0.208846 -0.951841
+ 2.307e+11Hz -0.209573 -0.9517
+ 2.308e+11Hz -0.210301 -0.951559
+ 2.309e+11Hz -0.211029 -0.951418
+ 2.31e+11Hz -0.211757 -0.951276
+ 2.311e+11Hz -0.212485 -0.951134
+ 2.312e+11Hz -0.213213 -0.950991
+ 2.313e+11Hz -0.213942 -0.950848
+ 2.314e+11Hz -0.214671 -0.950704
+ 2.315e+11Hz -0.2154 -0.950559
+ 2.316e+11Hz -0.21613 -0.950414
+ 2.317e+11Hz -0.21686 -0.950268
+ 2.318e+11Hz -0.21759 -0.950122
+ 2.319e+11Hz -0.21832 -0.949976
+ 2.32e+11Hz -0.21905 -0.949828
+ 2.321e+11Hz -0.219781 -0.94968
+ 2.322e+11Hz -0.220512 -0.949532
+ 2.323e+11Hz -0.221243 -0.949383
+ 2.324e+11Hz -0.221974 -0.949233
+ 2.325e+11Hz -0.222706 -0.949083
+ 2.326e+11Hz -0.223438 -0.948932
+ 2.327e+11Hz -0.22417 -0.948781
+ 2.328e+11Hz -0.224902 -0.948629
+ 2.329e+11Hz -0.225635 -0.948476
+ 2.33e+11Hz -0.226368 -0.948323
+ 2.331e+11Hz -0.227101 -0.948169
+ 2.332e+11Hz -0.227834 -0.948014
+ 2.333e+11Hz -0.228568 -0.947859
+ 2.334e+11Hz -0.229301 -0.947703
+ 2.335e+11Hz -0.230035 -0.947546
+ 2.336e+11Hz -0.230769 -0.947389
+ 2.337e+11Hz -0.231504 -0.947231
+ 2.338e+11Hz -0.232238 -0.947073
+ 2.339e+11Hz -0.232973 -0.946913
+ 2.34e+11Hz -0.233708 -0.946753
+ 2.341e+11Hz -0.234443 -0.946593
+ 2.342e+11Hz -0.235178 -0.946431
+ 2.343e+11Hz -0.235914 -0.946269
+ 2.344e+11Hz -0.23665 -0.946107
+ 2.345e+11Hz -0.237385 -0.945943
+ 2.346e+11Hz -0.238122 -0.945779
+ 2.347e+11Hz -0.238858 -0.945614
+ 2.348e+11Hz -0.239594 -0.945448
+ 2.349e+11Hz -0.240331 -0.945282
+ 2.35e+11Hz -0.241068 -0.945115
+ 2.351e+11Hz -0.241805 -0.944947
+ 2.352e+11Hz -0.242542 -0.944778
+ 2.353e+11Hz -0.243279 -0.944609
+ 2.354e+11Hz -0.244016 -0.944439
+ 2.355e+11Hz -0.244754 -0.944268
+ 2.356e+11Hz -0.245491 -0.944096
+ 2.357e+11Hz -0.246229 -0.943924
+ 2.358e+11Hz -0.246967 -0.943751
+ 2.359e+11Hz -0.247705 -0.943577
+ 2.36e+11Hz -0.248443 -0.943402
+ 2.361e+11Hz -0.249182 -0.943227
+ 2.362e+11Hz -0.24992 -0.94305
+ 2.363e+11Hz -0.250659 -0.942873
+ 2.364e+11Hz -0.251397 -0.942695
+ 2.365e+11Hz -0.252136 -0.942517
+ 2.366e+11Hz -0.252875 -0.942337
+ 2.367e+11Hz -0.253614 -0.942157
+ 2.368e+11Hz -0.254353 -0.941976
+ 2.369e+11Hz -0.255092 -0.941794
+ 2.37e+11Hz -0.255831 -0.941611
+ 2.371e+11Hz -0.25657 -0.941427
+ 2.372e+11Hz -0.257309 -0.941243
+ 2.373e+11Hz -0.258049 -0.941058
+ 2.374e+11Hz -0.258788 -0.940872
+ 2.375e+11Hz -0.259527 -0.940685
+ 2.376e+11Hz -0.260267 -0.940497
+ 2.377e+11Hz -0.261006 -0.940309
+ 2.378e+11Hz -0.261746 -0.94012
+ 2.379e+11Hz -0.262485 -0.93993
+ 2.38e+11Hz -0.263225 -0.939739
+ 2.381e+11Hz -0.263964 -0.939547
+ 2.382e+11Hz -0.264704 -0.939354
+ 2.383e+11Hz -0.265443 -0.939161
+ 2.384e+11Hz -0.266183 -0.938966
+ 2.385e+11Hz -0.266923 -0.938771
+ 2.386e+11Hz -0.267662 -0.938575
+ 2.387e+11Hz -0.268402 -0.938378
+ 2.388e+11Hz -0.269141 -0.938181
+ 2.389e+11Hz -0.26988 -0.937982
+ 2.39e+11Hz -0.27062 -0.937783
+ 2.391e+11Hz -0.271359 -0.937582
+ 2.392e+11Hz -0.272098 -0.937381
+ 2.393e+11Hz -0.272838 -0.937179
+ 2.394e+11Hz -0.273577 -0.936976
+ 2.395e+11Hz -0.274316 -0.936773
+ 2.396e+11Hz -0.275055 -0.936568
+ 2.397e+11Hz -0.275794 -0.936363
+ 2.398e+11Hz -0.276533 -0.936157
+ 2.399e+11Hz -0.277272 -0.93595
+ 2.4e+11Hz -0.27801 -0.935742
+ 2.401e+11Hz -0.278749 -0.935533
+ 2.402e+11Hz -0.279487 -0.935324
+ 2.403e+11Hz -0.280226 -0.935113
+ 2.404e+11Hz -0.280964 -0.934902
+ 2.405e+11Hz -0.281702 -0.93469
+ 2.406e+11Hz -0.28244 -0.934477
+ 2.407e+11Hz -0.283178 -0.934263
+ 2.408e+11Hz -0.283916 -0.934048
+ 2.409e+11Hz -0.284653 -0.933833
+ 2.41e+11Hz -0.285391 -0.933617
+ 2.411e+11Hz -0.286128 -0.933399
+ 2.412e+11Hz -0.286865 -0.933181
+ 2.413e+11Hz -0.287602 -0.932963
+ 2.414e+11Hz -0.288339 -0.932743
+ 2.415e+11Hz -0.289076 -0.932522
+ 2.416e+11Hz -0.289812 -0.932301
+ 2.417e+11Hz -0.290549 -0.932079
+ 2.418e+11Hz -0.291285 -0.931856
+ 2.419e+11Hz -0.292021 -0.931632
+ 2.42e+11Hz -0.292756 -0.931407
+ 2.421e+11Hz -0.293492 -0.931182
+ 2.422e+11Hz -0.294227 -0.930956
+ 2.423e+11Hz -0.294962 -0.930728
+ 2.424e+11Hz -0.295697 -0.930501
+ 2.425e+11Hz -0.296432 -0.930272
+ 2.426e+11Hz -0.297166 -0.930042
+ 2.427e+11Hz -0.297901 -0.929812
+ 2.428e+11Hz -0.298635 -0.929581
+ 2.429e+11Hz -0.299368 -0.929349
+ 2.43e+11Hz -0.300102 -0.929116
+ 2.431e+11Hz -0.300835 -0.928882
+ 2.432e+11Hz -0.301568 -0.928648
+ 2.433e+11Hz -0.302301 -0.928413
+ 2.434e+11Hz -0.303034 -0.928177
+ 2.435e+11Hz -0.303766 -0.92794
+ 2.436e+11Hz -0.304498 -0.927703
+ 2.437e+11Hz -0.30523 -0.927464
+ 2.438e+11Hz -0.305962 -0.927225
+ 2.439e+11Hz -0.306693 -0.926985
+ 2.44e+11Hz -0.307424 -0.926745
+ 2.441e+11Hz -0.308155 -0.926503
+ 2.442e+11Hz -0.308885 -0.926261
+ 2.443e+11Hz -0.309616 -0.926018
+ 2.444e+11Hz -0.310345 -0.925774
+ 2.445e+11Hz -0.311075 -0.92553
+ 2.446e+11Hz -0.311805 -0.925285
+ 2.447e+11Hz -0.312534 -0.925039
+ 2.448e+11Hz -0.313262 -0.924792
+ 2.449e+11Hz -0.313991 -0.924545
+ 2.45e+11Hz -0.314719 -0.924296
+ 2.451e+11Hz -0.315447 -0.924047
+ 2.452e+11Hz -0.316175 -0.923798
+ 2.453e+11Hz -0.316902 -0.923547
+ 2.454e+11Hz -0.317629 -0.923296
+ 2.455e+11Hz -0.318356 -0.923044
+ 2.456e+11Hz -0.319082 -0.922791
+ 2.457e+11Hz -0.319808 -0.922538
+ 2.458e+11Hz -0.320534 -0.922284
+ 2.459e+11Hz -0.321259 -0.922029
+ 2.46e+11Hz -0.321985 -0.921774
+ 2.461e+11Hz -0.32271 -0.921517
+ 2.462e+11Hz -0.323434 -0.92126
+ 2.463e+11Hz -0.324158 -0.921003
+ 2.464e+11Hz -0.324882 -0.920744
+ 2.465e+11Hz -0.325606 -0.920485
+ 2.466e+11Hz -0.326329 -0.920225
+ 2.467e+11Hz -0.327052 -0.919965
+ 2.468e+11Hz -0.327775 -0.919704
+ 2.469e+11Hz -0.328497 -0.919442
+ 2.47e+11Hz -0.329219 -0.919179
+ 2.471e+11Hz -0.329941 -0.918916
+ 2.472e+11Hz -0.330662 -0.918652
+ 2.473e+11Hz -0.331383 -0.918388
+ 2.474e+11Hz -0.332103 -0.918122
+ 2.475e+11Hz -0.332824 -0.917856
+ 2.476e+11Hz -0.333544 -0.91759
+ 2.477e+11Hz -0.334264 -0.917322
+ 2.478e+11Hz -0.334983 -0.917054
+ 2.479e+11Hz -0.335702 -0.916786
+ 2.48e+11Hz -0.336421 -0.916516
+ 2.481e+11Hz -0.337139 -0.916247
+ 2.482e+11Hz -0.337857 -0.915976
+ 2.483e+11Hz -0.338575 -0.915705
+ 2.484e+11Hz -0.339292 -0.915433
+ 2.485e+11Hz -0.340009 -0.91516
+ 2.486e+11Hz -0.340726 -0.914887
+ 2.487e+11Hz -0.341442 -0.914613
+ 2.488e+11Hz -0.342158 -0.914338
+ 2.489e+11Hz -0.342874 -0.914063
+ 2.49e+11Hz -0.343589 -0.913787
+ 2.491e+11Hz -0.344304 -0.913511
+ 2.492e+11Hz -0.345019 -0.913234
+ 2.493e+11Hz -0.345733 -0.912956
+ 2.494e+11Hz -0.346447 -0.912678
+ 2.495e+11Hz -0.347161 -0.912399
+ 2.496e+11Hz -0.347874 -0.912119
+ 2.497e+11Hz -0.348587 -0.911839
+ 2.498e+11Hz -0.3493 -0.911558
+ 2.499e+11Hz -0.350012 -0.911276
+ 2.5e+11Hz -0.350724 -0.910994
+ 2.501e+11Hz -0.351436 -0.910712
+ 2.502e+11Hz -0.352147 -0.910428
+ 2.503e+11Hz -0.352858 -0.910144
+ 2.504e+11Hz -0.353569 -0.909859
+ 2.505e+11Hz -0.354279 -0.909574
+ 2.506e+11Hz -0.354989 -0.909288
+ 2.507e+11Hz -0.355699 -0.909002
+ 2.508e+11Hz -0.356408 -0.908715
+ 2.509e+11Hz -0.357117 -0.908427
+ 2.51e+11Hz -0.357826 -0.908139
+ 2.511e+11Hz -0.358534 -0.90785
+ 2.512e+11Hz -0.359242 -0.90756
+ 2.513e+11Hz -0.35995 -0.90727
+ 2.514e+11Hz -0.360657 -0.906979
+ 2.515e+11Hz -0.361364 -0.906688
+ 2.516e+11Hz -0.36207 -0.906396
+ 2.517e+11Hz -0.362777 -0.906103
+ 2.518e+11Hz -0.363483 -0.90581
+ 2.519e+11Hz -0.364188 -0.905516
+ 2.52e+11Hz -0.364894 -0.905221
+ 2.521e+11Hz -0.365598 -0.904926
+ 2.522e+11Hz -0.366303 -0.904631
+ 2.523e+11Hz -0.367007 -0.904334
+ 2.524e+11Hz -0.367711 -0.904038
+ 2.525e+11Hz -0.368415 -0.90374
+ 2.526e+11Hz -0.369118 -0.903442
+ 2.527e+11Hz -0.369821 -0.903143
+ 2.528e+11Hz -0.370523 -0.902844
+ 2.529e+11Hz -0.371226 -0.902544
+ 2.53e+11Hz -0.371928 -0.902244
+ 2.531e+11Hz -0.372629 -0.901943
+ 2.532e+11Hz -0.37333 -0.901641
+ 2.533e+11Hz -0.374031 -0.901339
+ 2.534e+11Hz -0.374732 -0.901036
+ 2.535e+11Hz -0.375432 -0.900732
+ 2.536e+11Hz -0.376131 -0.900428
+ 2.537e+11Hz -0.376831 -0.900123
+ 2.538e+11Hz -0.37753 -0.899818
+ 2.539e+11Hz -0.378229 -0.899512
+ 2.54e+11Hz -0.378927 -0.899206
+ 2.541e+11Hz -0.379625 -0.898899
+ 2.542e+11Hz -0.380323 -0.898591
+ 2.543e+11Hz -0.38102 -0.898283
+ 2.544e+11Hz -0.381717 -0.897974
+ 2.545e+11Hz -0.382414 -0.897664
+ 2.546e+11Hz -0.38311 -0.897354
+ 2.547e+11Hz -0.383806 -0.897044
+ 2.548e+11Hz -0.384502 -0.896732
+ 2.549e+11Hz -0.385197 -0.896421
+ 2.55e+11Hz -0.385892 -0.896108
+ 2.551e+11Hz -0.386586 -0.895795
+ 2.552e+11Hz -0.38728 -0.895481
+ 2.553e+11Hz -0.387974 -0.895167
+ 2.554e+11Hz -0.388667 -0.894852
+ 2.555e+11Hz -0.38936 -0.894537
+ 2.556e+11Hz -0.390053 -0.894221
+ 2.557e+11Hz -0.390745 -0.893904
+ 2.558e+11Hz -0.391437 -0.893587
+ 2.559e+11Hz -0.392128 -0.893269
+ 2.56e+11Hz -0.392819 -0.892951
+ 2.561e+11Hz -0.39351 -0.892632
+ 2.562e+11Hz -0.3942 -0.892312
+ 2.563e+11Hz -0.39489 -0.891992
+ 2.564e+11Hz -0.39558 -0.891672
+ 2.565e+11Hz -0.396269 -0.89135
+ 2.566e+11Hz -0.396958 -0.891028
+ 2.567e+11Hz -0.397646 -0.890706
+ 2.568e+11Hz -0.398334 -0.890383
+ 2.569e+11Hz -0.399022 -0.890059
+ 2.57e+11Hz -0.399709 -0.889735
+ 2.571e+11Hz -0.400396 -0.88941
+ 2.572e+11Hz -0.401082 -0.889085
+ 2.573e+11Hz -0.401768 -0.888759
+ 2.574e+11Hz -0.402454 -0.888432
+ 2.575e+11Hz -0.403139 -0.888105
+ 2.576e+11Hz -0.403824 -0.887778
+ 2.577e+11Hz -0.404508 -0.887449
+ 2.578e+11Hz -0.405192 -0.887121
+ 2.579e+11Hz -0.405875 -0.886791
+ 2.58e+11Hz -0.406558 -0.886461
+ 2.581e+11Hz -0.407241 -0.886131
+ 2.582e+11Hz -0.407923 -0.8858
+ 2.583e+11Hz -0.408605 -0.885468
+ 2.584e+11Hz -0.409286 -0.885136
+ 2.585e+11Hz -0.409967 -0.884803
+ 2.586e+11Hz -0.410648 -0.88447
+ 2.587e+11Hz -0.411328 -0.884136
+ 2.588e+11Hz -0.412007 -0.883802
+ 2.589e+11Hz -0.412686 -0.883467
+ 2.59e+11Hz -0.413365 -0.883131
+ 2.591e+11Hz -0.414043 -0.882795
+ 2.592e+11Hz -0.414721 -0.882458
+ 2.593e+11Hz -0.415398 -0.882121
+ 2.594e+11Hz -0.416075 -0.881784
+ 2.595e+11Hz -0.416752 -0.881446
+ 2.596e+11Hz -0.417428 -0.881107
+ 2.597e+11Hz -0.418103 -0.880768
+ 2.598e+11Hz -0.418778 -0.880428
+ 2.599e+11Hz -0.419453 -0.880088
+ 2.6e+11Hz -0.420127 -0.879747
+ 2.601e+11Hz -0.420801 -0.879405
+ 2.602e+11Hz -0.421474 -0.879064
+ 2.603e+11Hz -0.422146 -0.878721
+ 2.604e+11Hz -0.422819 -0.878379
+ 2.605e+11Hz -0.42349 -0.878035
+ 2.606e+11Hz -0.424162 -0.877691
+ 2.607e+11Hz -0.424832 -0.877347
+ 2.608e+11Hz -0.425503 -0.877002
+ 2.609e+11Hz -0.426173 -0.876657
+ 2.61e+11Hz -0.426842 -0.876311
+ 2.611e+11Hz -0.427511 -0.875965
+ 2.612e+11Hz -0.428179 -0.875618
+ 2.613e+11Hz -0.428847 -0.875271
+ 2.614e+11Hz -0.429514 -0.874923
+ 2.615e+11Hz -0.430181 -0.874575
+ 2.616e+11Hz -0.430847 -0.874227
+ 2.617e+11Hz -0.431513 -0.873878
+ 2.618e+11Hz -0.432179 -0.873528
+ 2.619e+11Hz -0.432843 -0.873178
+ 2.62e+11Hz -0.433508 -0.872828
+ 2.621e+11Hz -0.434172 -0.872477
+ 2.622e+11Hz -0.434835 -0.872126
+ 2.623e+11Hz -0.435498 -0.871774
+ 2.624e+11Hz -0.43616 -0.871422
+ 2.625e+11Hz -0.436822 -0.87107
+ 2.626e+11Hz -0.437484 -0.870717
+ 2.627e+11Hz -0.438144 -0.870364
+ 2.628e+11Hz -0.438805 -0.87001
+ 2.629e+11Hz -0.439465 -0.869656
+ 2.63e+11Hz -0.440124 -0.869301
+ 2.631e+11Hz -0.440783 -0.868947
+ 2.632e+11Hz -0.441441 -0.868591
+ 2.633e+11Hz -0.442099 -0.868236
+ 2.634e+11Hz -0.442756 -0.86788
+ 2.635e+11Hz -0.443413 -0.867523
+ 2.636e+11Hz -0.444069 -0.867167
+ 2.637e+11Hz -0.444725 -0.86681
+ 2.638e+11Hz -0.44538 -0.866452
+ 2.639e+11Hz -0.446035 -0.866094
+ 2.64e+11Hz -0.44669 -0.865736
+ 2.641e+11Hz -0.447343 -0.865378
+ 2.642e+11Hz -0.447997 -0.865019
+ 2.643e+11Hz -0.448649 -0.86466
+ 2.644e+11Hz -0.449302 -0.8643
+ 2.645e+11Hz -0.449954 -0.863941
+ 2.646e+11Hz -0.450605 -0.863581
+ 2.647e+11Hz -0.451256 -0.86322
+ 2.648e+11Hz -0.451906 -0.86286
+ 2.649e+11Hz -0.452556 -0.862499
+ 2.65e+11Hz -0.453205 -0.862137
+ 2.651e+11Hz -0.453854 -0.861776
+ 2.652e+11Hz -0.454503 -0.861414
+ 2.653e+11Hz -0.455151 -0.861052
+ 2.654e+11Hz -0.455798 -0.86069
+ 2.655e+11Hz -0.456445 -0.860327
+ 2.656e+11Hz -0.457092 -0.859964
+ 2.657e+11Hz -0.457738 -0.859601
+ 2.658e+11Hz -0.458384 -0.859238
+ 2.659e+11Hz -0.459029 -0.858874
+ 2.66e+11Hz -0.459673 -0.85851
+ 2.661e+11Hz -0.460318 -0.858146
+ 2.662e+11Hz -0.460962 -0.857782
+ 2.663e+11Hz -0.461605 -0.857418
+ 2.664e+11Hz -0.462248 -0.857053
+ 2.665e+11Hz -0.46289 -0.856688
+ 2.666e+11Hz -0.463532 -0.856323
+ 2.667e+11Hz -0.464174 -0.855957
+ 2.668e+11Hz -0.464815 -0.855592
+ 2.669e+11Hz -0.465456 -0.855226
+ 2.67e+11Hz -0.466097 -0.85486
+ 2.671e+11Hz -0.466737 -0.854494
+ 2.672e+11Hz -0.467376 -0.854128
+ 2.673e+11Hz -0.468015 -0.853761
+ 2.674e+11Hz -0.468654 -0.853395
+ 2.675e+11Hz -0.469293 -0.853028
+ 2.676e+11Hz -0.469931 -0.852661
+ 2.677e+11Hz -0.470568 -0.852293
+ 2.678e+11Hz -0.471205 -0.851926
+ 2.679e+11Hz -0.471842 -0.851559
+ 2.68e+11Hz -0.472479 -0.851191
+ 2.681e+11Hz -0.473115 -0.850823
+ 2.682e+11Hz -0.473751 -0.850455
+ 2.683e+11Hz -0.474386 -0.850087
+ 2.684e+11Hz -0.475022 -0.849719
+ 2.685e+11Hz -0.475656 -0.849351
+ 2.686e+11Hz -0.476291 -0.848982
+ 2.687e+11Hz -0.476925 -0.848613
+ 2.688e+11Hz -0.477559 -0.848245
+ 2.689e+11Hz -0.478193 -0.847876
+ 2.69e+11Hz -0.478826 -0.847507
+ 2.691e+11Hz -0.479459 -0.847138
+ 2.692e+11Hz -0.480091 -0.846768
+ 2.693e+11Hz -0.480724 -0.846399
+ 2.694e+11Hz -0.481356 -0.846029
+ 2.695e+11Hz -0.481988 -0.84566
+ 2.696e+11Hz -0.482619 -0.84529
+ 2.697e+11Hz -0.483251 -0.84492
+ 2.698e+11Hz -0.483882 -0.84455
+ 2.699e+11Hz -0.484513 -0.84418
+ 2.7e+11Hz -0.485143 -0.84381
+ 2.701e+11Hz -0.485774 -0.84344
+ 2.702e+11Hz -0.486404 -0.843069
+ 2.703e+11Hz -0.487034 -0.842699
+ 2.704e+11Hz -0.487664 -0.842328
+ 2.705e+11Hz -0.488293 -0.841957
+ 2.706e+11Hz -0.488923 -0.841586
+ 2.707e+11Hz -0.489552 -0.841215
+ 2.708e+11Hz -0.490181 -0.840844
+ 2.709e+11Hz -0.49081 -0.840473
+ 2.71e+11Hz -0.491439 -0.840102
+ 2.711e+11Hz -0.492067 -0.83973
+ 2.712e+11Hz -0.492696 -0.839359
+ 2.713e+11Hz -0.493324 -0.838987
+ 2.714e+11Hz -0.493952 -0.838615
+ 2.715e+11Hz -0.49458 -0.838243
+ 2.716e+11Hz -0.495208 -0.837871
+ 2.717e+11Hz -0.495836 -0.837499
+ 2.718e+11Hz -0.496464 -0.837127
+ 2.719e+11Hz -0.497092 -0.836754
+ 2.72e+11Hz -0.497719 -0.836382
+ 2.721e+11Hz -0.498347 -0.836009
+ 2.722e+11Hz -0.498974 -0.835636
+ 2.723e+11Hz -0.499601 -0.835263
+ 2.724e+11Hz -0.500229 -0.83489
+ 2.725e+11Hz -0.500856 -0.834517
+ 2.726e+11Hz -0.501483 -0.834144
+ 2.727e+11Hz -0.50211 -0.83377
+ 2.728e+11Hz -0.502738 -0.833396
+ 2.729e+11Hz -0.503365 -0.833022
+ 2.73e+11Hz -0.503992 -0.832648
+ 2.731e+11Hz -0.504619 -0.832274
+ 2.732e+11Hz -0.505246 -0.8319
+ 2.733e+11Hz -0.505873 -0.831525
+ 2.734e+11Hz -0.5065 -0.83115
+ 2.735e+11Hz -0.507127 -0.830775
+ 2.736e+11Hz -0.507755 -0.8304
+ 2.737e+11Hz -0.508382 -0.830025
+ 2.738e+11Hz -0.509009 -0.829649
+ 2.739e+11Hz -0.509636 -0.829273
+ 2.74e+11Hz -0.510264 -0.828897
+ 2.741e+11Hz -0.510891 -0.828521
+ 2.742e+11Hz -0.511519 -0.828145
+ 2.743e+11Hz -0.512146 -0.827768
+ 2.744e+11Hz -0.512774 -0.827391
+ 2.745e+11Hz -0.513401 -0.827014
+ 2.746e+11Hz -0.514029 -0.826636
+ 2.747e+11Hz -0.514657 -0.826259
+ 2.748e+11Hz -0.515285 -0.825881
+ 2.749e+11Hz -0.515913 -0.825502
+ 2.75e+11Hz -0.516541 -0.825124
+ 2.751e+11Hz -0.517169 -0.824745
+ 2.752e+11Hz -0.517798 -0.824366
+ 2.753e+11Hz -0.518426 -0.823987
+ 2.754e+11Hz -0.519055 -0.823607
+ 2.755e+11Hz -0.519683 -0.823227
+ 2.756e+11Hz -0.520312 -0.822846
+ 2.757e+11Hz -0.520941 -0.822466
+ 2.758e+11Hz -0.52157 -0.822084
+ 2.759e+11Hz -0.522199 -0.821703
+ 2.76e+11Hz -0.522829 -0.821321
+ 2.761e+11Hz -0.523458 -0.820939
+ 2.762e+11Hz -0.524088 -0.820556
+ 2.763e+11Hz -0.524718 -0.820174
+ 2.764e+11Hz -0.525348 -0.81979
+ 2.765e+11Hz -0.525978 -0.819406
+ 2.766e+11Hz -0.526608 -0.819022
+ 2.767e+11Hz -0.527238 -0.818638
+ 2.768e+11Hz -0.527869 -0.818253
+ 2.769e+11Hz -0.5285 -0.817867
+ 2.77e+11Hz -0.529131 -0.817481
+ 2.771e+11Hz -0.529762 -0.817095
+ 2.772e+11Hz -0.530393 -0.816708
+ 2.773e+11Hz -0.531024 -0.816321
+ 2.774e+11Hz -0.531656 -0.815933
+ 2.775e+11Hz -0.532287 -0.815545
+ 2.776e+11Hz -0.532919 -0.815156
+ 2.777e+11Hz -0.533551 -0.814767
+ 2.778e+11Hz -0.534184 -0.814377
+ 2.779e+11Hz -0.534816 -0.813987
+ 2.78e+11Hz -0.535448 -0.813596
+ 2.781e+11Hz -0.536081 -0.813205
+ 2.782e+11Hz -0.536714 -0.812813
+ 2.783e+11Hz -0.537347 -0.81242
+ 2.784e+11Hz -0.53798 -0.812027
+ 2.785e+11Hz -0.538613 -0.811633
+ 2.786e+11Hz -0.539247 -0.811239
+ 2.787e+11Hz -0.53988 -0.810844
+ 2.788e+11Hz -0.540514 -0.810449
+ 2.789e+11Hz -0.541148 -0.810053
+ 2.79e+11Hz -0.541782 -0.809656
+ 2.791e+11Hz -0.542416 -0.809258
+ 2.792e+11Hz -0.54305 -0.80886
+ 2.793e+11Hz -0.543685 -0.808462
+ 2.794e+11Hz -0.544319 -0.808062
+ 2.795e+11Hz -0.544954 -0.807662
+ 2.796e+11Hz -0.545589 -0.807262
+ 2.797e+11Hz -0.546224 -0.80686
+ 2.798e+11Hz -0.546859 -0.806458
+ 2.799e+11Hz -0.547494 -0.806055
+ 2.8e+11Hz -0.548129 -0.805652
+ 2.801e+11Hz -0.548765 -0.805248
+ 2.802e+11Hz -0.5494 -0.804843
+ 2.803e+11Hz -0.550036 -0.804437
+ 2.804e+11Hz -0.550671 -0.804031
+ 2.805e+11Hz -0.551307 -0.803623
+ 2.806e+11Hz -0.551943 -0.803215
+ 2.807e+11Hz -0.552579 -0.802807
+ 2.808e+11Hz -0.553215 -0.802397
+ 2.809e+11Hz -0.553851 -0.801987
+ 2.81e+11Hz -0.554487 -0.801576
+ 2.811e+11Hz -0.555123 -0.801164
+ 2.812e+11Hz -0.555759 -0.800751
+ 2.813e+11Hz -0.556395 -0.800338
+ 2.814e+11Hz -0.557031 -0.799923
+ 2.815e+11Hz -0.557667 -0.799508
+ 2.816e+11Hz -0.558303 -0.799092
+ 2.817e+11Hz -0.55894 -0.798675
+ 2.818e+11Hz -0.559576 -0.798258
+ 2.819e+11Hz -0.560212 -0.797839
+ 2.82e+11Hz -0.560848 -0.79742
+ 2.821e+11Hz -0.561484 -0.797
+ 2.822e+11Hz -0.56212 -0.796579
+ 2.823e+11Hz -0.562756 -0.796157
+ 2.824e+11Hz -0.563392 -0.795734
+ 2.825e+11Hz -0.564028 -0.79531
+ 2.826e+11Hz -0.564664 -0.794885
+ 2.827e+11Hz -0.5653 -0.79446
+ 2.828e+11Hz -0.565935 -0.794033
+ 2.829e+11Hz -0.566571 -0.793606
+ 2.83e+11Hz -0.567207 -0.793178
+ 2.831e+11Hz -0.567842 -0.792749
+ 2.832e+11Hz -0.568477 -0.792319
+ 2.833e+11Hz -0.569112 -0.791888
+ 2.834e+11Hz -0.569747 -0.791456
+ 2.835e+11Hz -0.570382 -0.791023
+ 2.836e+11Hz -0.571017 -0.790589
+ 2.837e+11Hz -0.571651 -0.790155
+ 2.838e+11Hz -0.572285 -0.789719
+ 2.839e+11Hz -0.572919 -0.789283
+ 2.84e+11Hz -0.573553 -0.788845
+ 2.841e+11Hz -0.574187 -0.788407
+ 2.842e+11Hz -0.57482 -0.787968
+ 2.843e+11Hz -0.575454 -0.787527
+ 2.844e+11Hz -0.576087 -0.787086
+ 2.845e+11Hz -0.57672 -0.786644
+ 2.846e+11Hz -0.577352 -0.786201
+ 2.847e+11Hz -0.577984 -0.785757
+ 2.848e+11Hz -0.578616 -0.785312
+ 2.849e+11Hz -0.579248 -0.784866
+ 2.85e+11Hz -0.579879 -0.784419
+ 2.851e+11Hz -0.58051 -0.783972
+ 2.852e+11Hz -0.581141 -0.783523
+ 2.853e+11Hz -0.581772 -0.783073
+ 2.854e+11Hz -0.582402 -0.782623
+ 2.855e+11Hz -0.583032 -0.782171
+ 2.856e+11Hz -0.583661 -0.781719
+ 2.857e+11Hz -0.58429 -0.781265
+ 2.858e+11Hz -0.584919 -0.780811
+ 2.859e+11Hz -0.585547 -0.780356
+ 2.86e+11Hz -0.586175 -0.779899
+ 2.861e+11Hz -0.586802 -0.779442
+ 2.862e+11Hz -0.58743 -0.778984
+ 2.863e+11Hz -0.588056 -0.778525
+ 2.864e+11Hz -0.588683 -0.778065
+ 2.865e+11Hz -0.589308 -0.777605
+ 2.866e+11Hz -0.589934 -0.777143
+ 2.867e+11Hz -0.590559 -0.77668
+ 2.868e+11Hz -0.591183 -0.776217
+ 2.869e+11Hz -0.591807 -0.775752
+ 2.87e+11Hz -0.592431 -0.775287
+ 2.871e+11Hz -0.593054 -0.77482
+ 2.872e+11Hz -0.593677 -0.774353
+ 2.873e+11Hz -0.594299 -0.773885
+ 2.874e+11Hz -0.59492 -0.773416
+ 2.875e+11Hz -0.595541 -0.772947
+ 2.876e+11Hz -0.596162 -0.772476
+ 2.877e+11Hz -0.596782 -0.772004
+ 2.878e+11Hz -0.597401 -0.771532
+ 2.879e+11Hz -0.59802 -0.771059
+ 2.88e+11Hz -0.598638 -0.770585
+ 2.881e+11Hz -0.599256 -0.77011
+ 2.882e+11Hz -0.599873 -0.769634
+ 2.883e+11Hz -0.60049 -0.769157
+ 2.884e+11Hz -0.601106 -0.76868
+ 2.885e+11Hz -0.601722 -0.768201
+ 2.886e+11Hz -0.602336 -0.767722
+ 2.887e+11Hz -0.602951 -0.767242
+ 2.888e+11Hz -0.603564 -0.766762
+ 2.889e+11Hz -0.604177 -0.76628
+ 2.89e+11Hz -0.60479 -0.765798
+ 2.891e+11Hz -0.605402 -0.765315
+ 2.892e+11Hz -0.606013 -0.764831
+ 2.893e+11Hz -0.606623 -0.764346
+ 2.894e+11Hz -0.607233 -0.763861
+ 2.895e+11Hz -0.607843 -0.763374
+ 2.896e+11Hz -0.608451 -0.762888
+ 2.897e+11Hz -0.609059 -0.7624
+ 2.898e+11Hz -0.609666 -0.761911
+ 2.899e+11Hz -0.610273 -0.761422
+ 2.9e+11Hz -0.610879 -0.760932
+ 2.901e+11Hz -0.611484 -0.760442
+ 2.902e+11Hz -0.612089 -0.759951
+ 2.903e+11Hz -0.612693 -0.759459
+ 2.904e+11Hz -0.613296 -0.758966
+ 2.905e+11Hz -0.613899 -0.758473
+ 2.906e+11Hz -0.614501 -0.757978
+ 2.907e+11Hz -0.615102 -0.757484
+ 2.908e+11Hz -0.615703 -0.756988
+ 2.909e+11Hz -0.616302 -0.756492
+ 2.91e+11Hz -0.616902 -0.755996
+ 2.911e+11Hz -0.6175 -0.755498
+ 2.912e+11Hz -0.618098 -0.755
+ 2.913e+11Hz -0.618695 -0.754502
+ 2.914e+11Hz -0.619291 -0.754003
+ 2.915e+11Hz -0.619887 -0.753503
+ 2.916e+11Hz -0.620482 -0.753003
+ 2.917e+11Hz -0.621076 -0.752502
+ 2.918e+11Hz -0.62167 -0.752
+ 2.919e+11Hz -0.622262 -0.751498
+ 2.92e+11Hz -0.622855 -0.750995
+ 2.921e+11Hz -0.623446 -0.750492
+ 2.922e+11Hz -0.624037 -0.749988
+ 2.923e+11Hz -0.624627 -0.749484
+ 2.924e+11Hz -0.625216 -0.748979
+ 2.925e+11Hz -0.625805 -0.748473
+ 2.926e+11Hz -0.626392 -0.747967
+ 2.927e+11Hz -0.62698 -0.747461
+ 2.928e+11Hz -0.627566 -0.746954
+ 2.929e+11Hz -0.628152 -0.746446
+ 2.93e+11Hz -0.628737 -0.745938
+ 2.931e+11Hz -0.629322 -0.74543
+ 2.932e+11Hz -0.629905 -0.744921
+ 2.933e+11Hz -0.630488 -0.744411
+ 2.934e+11Hz -0.631071 -0.743901
+ 2.935e+11Hz -0.631652 -0.743391
+ 2.936e+11Hz -0.632233 -0.74288
+ 2.937e+11Hz -0.632813 -0.742369
+ 2.938e+11Hz -0.633393 -0.741857
+ 2.939e+11Hz -0.633972 -0.741345
+ 2.94e+11Hz -0.63455 -0.740832
+ 2.941e+11Hz -0.635128 -0.740319
+ 2.942e+11Hz -0.635705 -0.739805
+ 2.943e+11Hz -0.636281 -0.739291
+ 2.944e+11Hz -0.636856 -0.738777
+ 2.945e+11Hz -0.637431 -0.738262
+ 2.946e+11Hz -0.638005 -0.737747
+ 2.947e+11Hz -0.638579 -0.737231
+ 2.948e+11Hz -0.639152 -0.736716
+ 2.949e+11Hz -0.639724 -0.736199
+ 2.95e+11Hz -0.640296 -0.735682
+ 2.951e+11Hz -0.640867 -0.735165
+ 2.952e+11Hz -0.641437 -0.734648
+ 2.953e+11Hz -0.642007 -0.73413
+ 2.954e+11Hz -0.642576 -0.733612
+ 2.955e+11Hz -0.643144 -0.733093
+ 2.956e+11Hz -0.643712 -0.732574
+ 2.957e+11Hz -0.644279 -0.732055
+ 2.958e+11Hz -0.644846 -0.731535
+ 2.959e+11Hz -0.645412 -0.731015
+ 2.96e+11Hz -0.645978 -0.730494
+ 2.961e+11Hz -0.646542 -0.729974
+ 2.962e+11Hz -0.647107 -0.729452
+ 2.963e+11Hz -0.64767 -0.728931
+ 2.964e+11Hz -0.648233 -0.728409
+ 2.965e+11Hz -0.648796 -0.727887
+ 2.966e+11Hz -0.649358 -0.727364
+ 2.967e+11Hz -0.649919 -0.726842
+ 2.968e+11Hz -0.65048 -0.726318
+ 2.969e+11Hz -0.65104 -0.725795
+ 2.97e+11Hz -0.651599 -0.725271
+ 2.971e+11Hz -0.652158 -0.724747
+ 2.972e+11Hz -0.652717 -0.724222
+ 2.973e+11Hz -0.653275 -0.723698
+ 2.974e+11Hz -0.653832 -0.723172
+ 2.975e+11Hz -0.654389 -0.722647
+ 2.976e+11Hz -0.654946 -0.722121
+ 2.977e+11Hz -0.655501 -0.721595
+ 2.978e+11Hz -0.656057 -0.721069
+ 2.979e+11Hz -0.656612 -0.720542
+ 2.98e+11Hz -0.657166 -0.720015
+ 2.981e+11Hz -0.65772 -0.719487
+ 2.982e+11Hz -0.658273 -0.718959
+ 2.983e+11Hz -0.658826 -0.718431
+ 2.984e+11Hz -0.659378 -0.717903
+ 2.985e+11Hz -0.659929 -0.717374
+ 2.986e+11Hz -0.660481 -0.716845
+ 2.987e+11Hz -0.661031 -0.716316
+ 2.988e+11Hz -0.661582 -0.715786
+ 2.989e+11Hz -0.662131 -0.715256
+ 2.99e+11Hz -0.662681 -0.714725
+ 2.991e+11Hz -0.66323 -0.714194
+ 2.992e+11Hz -0.663778 -0.713663
+ 2.993e+11Hz -0.664326 -0.713132
+ 2.994e+11Hz -0.664873 -0.7126
+ 2.995e+11Hz -0.66542 -0.712068
+ 2.996e+11Hz -0.665967 -0.711535
+ 2.997e+11Hz -0.666513 -0.711002
+ 2.998e+11Hz -0.667058 -0.710469
+ 2.999e+11Hz -0.667603 -0.709936
+ 3e+11Hz -0.668148 -0.709402
+ ]

A22 %vd(20 3) %vd(22, 3) xfer4
.model xfer4 xfer R_I=true table=[
+ 0Hz 0.0047718 0
+ 1e+08Hz 0.00477202 3.3416e-06
+ 2e+08Hz 0.00477265 6.6748e-06
+ 3e+08Hz 0.0047737 9.99121e-06
+ 4e+08Hz 0.00477517 1.32825e-05
+ 5e+08Hz 0.00477706 1.65402e-05
+ 6e+08Hz 0.00477937 1.9756e-05
+ 7e+08Hz 0.0047821 2.29215e-05
+ 8e+08Hz 0.00478524 2.60286e-05
+ 9e+08Hz 0.0047888 2.90688e-05
+ 1e+09Hz 0.00479277 3.20341e-05
+ 1.1e+09Hz 0.00479716 3.49161e-05
+ 1.2e+09Hz 0.00480195 3.77067e-05
+ 1.3e+09Hz 0.00480715 4.03978e-05
+ 1.4e+09Hz 0.00481276 4.29814e-05
+ 1.5e+09Hz 0.00481877 4.54495e-05
+ 1.6e+09Hz 0.00482518 4.77941e-05
+ 1.7e+09Hz 0.00483198 5.00074e-05
+ 1.8e+09Hz 0.00483919 5.20816e-05
+ 1.9e+09Hz 0.00484678 5.40089e-05
+ 2e+09Hz 0.00485476 5.57818e-05
+ 2.1e+09Hz 0.00486313 5.73926e-05
+ 2.2e+09Hz 0.00487188 5.88339e-05
+ 2.3e+09Hz 0.00488101 6.00983e-05
+ 2.4e+09Hz 0.00489051 6.11784e-05
+ 2.5e+09Hz 0.00490038 6.20672e-05
+ 2.6e+09Hz 0.00491061 6.27574e-05
+ 2.7e+09Hz 0.00492121 6.32421e-05
+ 2.8e+09Hz 0.00493216 6.35144e-05
+ 2.9e+09Hz 0.00494347 6.35675e-05
+ 3e+09Hz 0.00495512 6.33948e-05
+ 3.1e+09Hz 0.00496711 6.29896e-05
+ 3.2e+09Hz 0.00497945 6.23456e-05
+ 3.3e+09Hz 0.00499211 6.14564e-05
+ 3.4e+09Hz 0.0050051 6.03159e-05
+ 3.5e+09Hz 0.00501841 5.89179e-05
+ 3.6e+09Hz 0.00503204 5.72566e-05
+ 3.7e+09Hz 0.00504598 5.53262e-05
+ 3.8e+09Hz 0.00506022 5.3121e-05
+ 3.9e+09Hz 0.00507476 5.06354e-05
+ 4e+09Hz 0.00508959 4.78642e-05
+ 4.1e+09Hz 0.00510471 4.48019e-05
+ 4.2e+09Hz 0.00512011 4.14436e-05
+ 4.3e+09Hz 0.00513579 3.77843e-05
+ 4.4e+09Hz 0.00515173 3.38191e-05
+ 4.5e+09Hz 0.00516793 2.95435e-05
+ 4.6e+09Hz 0.00518439 2.49528e-05
+ 4.7e+09Hz 0.0052011 2.00428e-05
+ 4.8e+09Hz 0.00521804 1.48093e-05
+ 4.9e+09Hz 0.00523522 9.24808e-06
+ 5e+09Hz 0.00525263 3.3554e-06
+ 5.1e+09Hz 0.00527026 -2.87253e-06
+ 5.2e+09Hz 0.00528811 -9.43928e-06
+ 5.3e+09Hz 0.00530616 -1.63483e-05
+ 5.4e+09Hz 0.00532441 -2.36027e-05
+ 5.5e+09Hz 0.00534285 -3.12058e-05
+ 5.6e+09Hz 0.00536148 -3.91605e-05
+ 5.7e+09Hz 0.00538029 -4.74694e-05
+ 5.8e+09Hz 0.00539927 -5.61353e-05
+ 5.9e+09Hz 0.00541841 -6.51606e-05
+ 6e+09Hz 0.00543771 -7.45476e-05
+ 6.1e+09Hz 0.00545716 -8.42984e-05
+ 6.2e+09Hz 0.00547675 -9.44149e-05
+ 6.3e+09Hz 0.00549648 -0.000104899
+ 6.4e+09Hz 0.00551633 -0.000115753
+ 6.5e+09Hz 0.0055363 -0.000126977
+ 6.6e+09Hz 0.00555639 -0.000138573
+ 6.7e+09Hz 0.00557658 -0.000150542
+ 6.8e+09Hz 0.00559687 -0.000162886
+ 6.9e+09Hz 0.00561724 -0.000175605
+ 7e+09Hz 0.00563771 -0.0001887
+ 7.1e+09Hz 0.00565825 -0.00020217
+ 7.2e+09Hz 0.00567885 -0.000216018
+ 7.3e+09Hz 0.00569952 -0.000230243
+ 7.4e+09Hz 0.00572024 -0.000244844
+ 7.5e+09Hz 0.00574101 -0.000259822
+ 7.6e+09Hz 0.00576182 -0.000275178
+ 7.7e+09Hz 0.00578266 -0.000290909
+ 7.8e+09Hz 0.00580352 -0.000307016
+ 7.9e+09Hz 0.00582441 -0.000323498
+ 8e+09Hz 0.0058453 -0.000340355
+ 8.1e+09Hz 0.0058662 -0.000357584
+ 8.2e+09Hz 0.00588709 -0.000375186
+ 8.3e+09Hz 0.00590798 -0.000393159
+ 8.4e+09Hz 0.00592884 -0.000411502
+ 8.5e+09Hz 0.00594969 -0.000430212
+ 8.6e+09Hz 0.0059705 -0.000449289
+ 8.7e+09Hz 0.00599128 -0.00046873
+ 8.8e+09Hz 0.00601201 -0.000488534
+ 8.9e+09Hz 0.0060327 -0.000508699
+ 9e+09Hz 0.00605332 -0.000529222
+ 9.1e+09Hz 0.00607388 -0.000550101
+ 9.2e+09Hz 0.00609438 -0.000571334
+ 9.3e+09Hz 0.0061148 -0.000592918
+ 9.4e+09Hz 0.00613513 -0.00061485
+ 9.5e+09Hz 0.00615538 -0.000637128
+ 9.6e+09Hz 0.00617553 -0.000659749
+ 9.7e+09Hz 0.00619559 -0.00068271
+ 9.8e+09Hz 0.00621554 -0.000706007
+ 9.9e+09Hz 0.00623537 -0.000729638
+ 1e+10Hz 0.00625509 -0.0007536
+ 1.01e+10Hz 0.00627469 -0.000777888
+ 1.02e+10Hz 0.00629416 -0.000802499
+ 1.03e+10Hz 0.0063135 -0.00082743
+ 1.04e+10Hz 0.0063327 -0.000852677
+ 1.05e+10Hz 0.00635175 -0.000878236
+ 1.06e+10Hz 0.00637065 -0.000904103
+ 1.07e+10Hz 0.00638941 -0.000930275
+ 1.08e+10Hz 0.006408 -0.000956747
+ 1.09e+10Hz 0.00642643 -0.000983515
+ 1.1e+10Hz 0.00644469 -0.00101058
+ 1.11e+10Hz 0.00646278 -0.00103792
+ 1.12e+10Hz 0.00648069 -0.00106555
+ 1.13e+10Hz 0.00649842 -0.00109346
+ 1.14e+10Hz 0.00651597 -0.00112165
+ 1.15e+10Hz 0.00653332 -0.0011501
+ 1.16e+10Hz 0.00655049 -0.00117882
+ 1.17e+10Hz 0.00656745 -0.0012078
+ 1.18e+10Hz 0.00658422 -0.00123704
+ 1.19e+10Hz 0.00660078 -0.00126653
+ 1.2e+10Hz 0.00661713 -0.00129626
+ 1.21e+10Hz 0.00663328 -0.00132624
+ 1.22e+10Hz 0.0066492 -0.00135645
+ 1.23e+10Hz 0.00666491 -0.0013869
+ 1.24e+10Hz 0.0066804 -0.00141757
+ 1.25e+10Hz 0.00669567 -0.00144846
+ 1.26e+10Hz 0.00671071 -0.00147957
+ 1.27e+10Hz 0.00672552 -0.00151089
+ 1.28e+10Hz 0.0067401 -0.00154242
+ 1.29e+10Hz 0.00675444 -0.00157415
+ 1.3e+10Hz 0.00676855 -0.00160607
+ 1.31e+10Hz 0.00678242 -0.00163819
+ 1.32e+10Hz 0.00679605 -0.00167049
+ 1.33e+10Hz 0.00680944 -0.00170297
+ 1.34e+10Hz 0.00682259 -0.00173563
+ 1.35e+10Hz 0.00683548 -0.00176846
+ 1.36e+10Hz 0.00684813 -0.00180146
+ 1.37e+10Hz 0.00686054 -0.00183461
+ 1.38e+10Hz 0.00687269 -0.00186792
+ 1.39e+10Hz 0.00688459 -0.00190138
+ 1.4e+10Hz 0.00689623 -0.00193498
+ 1.41e+10Hz 0.00690763 -0.00196872
+ 1.42e+10Hz 0.00691877 -0.00200259
+ 1.43e+10Hz 0.00692965 -0.0020366
+ 1.44e+10Hz 0.00694028 -0.00207073
+ 1.45e+10Hz 0.00695065 -0.00210497
+ 1.46e+10Hz 0.00696076 -0.00213933
+ 1.47e+10Hz 0.00697062 -0.0021738
+ 1.48e+10Hz 0.00698022 -0.00220837
+ 1.49e+10Hz 0.00698956 -0.00224303
+ 1.5e+10Hz 0.00699865 -0.00227779
+ 1.51e+10Hz 0.00700747 -0.00231264
+ 1.52e+10Hz 0.00701604 -0.00234757
+ 1.53e+10Hz 0.00702435 -0.00238258
+ 1.54e+10Hz 0.00703241 -0.00241767
+ 1.55e+10Hz 0.00704021 -0.00245282
+ 1.56e+10Hz 0.00704775 -0.00248803
+ 1.57e+10Hz 0.00705504 -0.0025233
+ 1.58e+10Hz 0.00706207 -0.00255863
+ 1.59e+10Hz 0.00706885 -0.00259401
+ 1.6e+10Hz 0.00707538 -0.00262943
+ 1.61e+10Hz 0.00708166 -0.00266489
+ 1.62e+10Hz 0.00708769 -0.00270038
+ 1.63e+10Hz 0.00709347 -0.00273591
+ 1.64e+10Hz 0.007099 -0.00277146
+ 1.65e+10Hz 0.00710429 -0.00280704
+ 1.66e+10Hz 0.00710933 -0.00284263
+ 1.67e+10Hz 0.00711413 -0.00287824
+ 1.68e+10Hz 0.00711869 -0.00291386
+ 1.69e+10Hz 0.007123 -0.00294948
+ 1.7e+10Hz 0.00712709 -0.0029851
+ 1.71e+10Hz 0.00713093 -0.00302072
+ 1.72e+10Hz 0.00713454 -0.00305634
+ 1.73e+10Hz 0.00713792 -0.00309194
+ 1.74e+10Hz 0.00714107 -0.00312753
+ 1.75e+10Hz 0.007144 -0.0031631
+ 1.76e+10Hz 0.0071467 -0.00319865
+ 1.77e+10Hz 0.00714917 -0.00323418
+ 1.78e+10Hz 0.00715143 -0.00326967
+ 1.79e+10Hz 0.00715346 -0.00330514
+ 1.8e+10Hz 0.00715529 -0.00334057
+ 1.81e+10Hz 0.0071569 -0.00337596
+ 1.82e+10Hz 0.0071583 -0.00341131
+ 1.83e+10Hz 0.00715949 -0.00344661
+ 1.84e+10Hz 0.00716048 -0.00348187
+ 1.85e+10Hz 0.00716126 -0.00351707
+ 1.86e+10Hz 0.00716185 -0.00355222
+ 1.87e+10Hz 0.00716224 -0.00358732
+ 1.88e+10Hz 0.00716243 -0.00362236
+ 1.89e+10Hz 0.00716244 -0.00365733
+ 1.9e+10Hz 0.00716225 -0.00369224
+ 1.91e+10Hz 0.00716189 -0.00372709
+ 1.92e+10Hz 0.00716134 -0.00376186
+ 1.93e+10Hz 0.00716061 -0.00379657
+ 1.94e+10Hz 0.00715971 -0.0038312
+ 1.95e+10Hz 0.00715863 -0.00386576
+ 1.96e+10Hz 0.00715739 -0.00390024
+ 1.97e+10Hz 0.00715598 -0.00393464
+ 1.98e+10Hz 0.00715441 -0.00396895
+ 1.99e+10Hz 0.00715267 -0.00400319
+ 2e+10Hz 0.00715079 -0.00403734
+ 2.01e+10Hz 0.00714874 -0.00407141
+ 2.02e+10Hz 0.00714655 -0.00410539
+ 2.03e+10Hz 0.00714421 -0.00413928
+ 2.04e+10Hz 0.00714173 -0.00417308
+ 2.05e+10Hz 0.0071391 -0.00420679
+ 2.06e+10Hz 0.00713634 -0.0042404
+ 2.07e+10Hz 0.00713345 -0.00427393
+ 2.08e+10Hz 0.00713043 -0.00430736
+ 2.09e+10Hz 0.00712727 -0.00434069
+ 2.1e+10Hz 0.007124 -0.00437393
+ 2.11e+10Hz 0.0071206 -0.00440707
+ 2.12e+10Hz 0.00711709 -0.00444012
+ 2.13e+10Hz 0.00711346 -0.00447306
+ 2.14e+10Hz 0.00710972 -0.00450591
+ 2.15e+10Hz 0.00710587 -0.00453866
+ 2.16e+10Hz 0.00710192 -0.00457131
+ 2.17e+10Hz 0.00709786 -0.00460386
+ 2.18e+10Hz 0.00709371 -0.00463632
+ 2.19e+10Hz 0.00708946 -0.00466867
+ 2.2e+10Hz 0.00708512 -0.00470093
+ 2.21e+10Hz 0.00708069 -0.00473308
+ 2.22e+10Hz 0.00707617 -0.00476514
+ 2.23e+10Hz 0.00707157 -0.0047971
+ 2.24e+10Hz 0.00706689 -0.00482896
+ 2.25e+10Hz 0.00706213 -0.00486072
+ 2.26e+10Hz 0.0070573 -0.00489238
+ 2.27e+10Hz 0.00705239 -0.00492395
+ 2.28e+10Hz 0.00704742 -0.00495542
+ 2.29e+10Hz 0.00704238 -0.0049868
+ 2.3e+10Hz 0.00703728 -0.00501808
+ 2.31e+10Hz 0.00703211 -0.00504927
+ 2.32e+10Hz 0.00702689 -0.00508036
+ 2.33e+10Hz 0.00702161 -0.00511136
+ 2.34e+10Hz 0.00701628 -0.00514227
+ 2.35e+10Hz 0.0070109 -0.00517309
+ 2.36e+10Hz 0.00700547 -0.00520382
+ 2.37e+10Hz 0.00699999 -0.00523446
+ 2.38e+10Hz 0.00699447 -0.00526501
+ 2.39e+10Hz 0.00698891 -0.00529548
+ 2.4e+10Hz 0.00698331 -0.00532587
+ 2.41e+10Hz 0.00697767 -0.00535617
+ 2.42e+10Hz 0.006972 -0.00538639
+ 2.43e+10Hz 0.0069663 -0.00541653
+ 2.44e+10Hz 0.00696057 -0.00544659
+ 2.45e+10Hz 0.0069548 -0.00547657
+ 2.46e+10Hz 0.00694902 -0.00550648
+ 2.47e+10Hz 0.0069432 -0.00553631
+ 2.48e+10Hz 0.00693737 -0.00556607
+ 2.49e+10Hz 0.00693151 -0.00559576
+ 2.5e+10Hz 0.00692563 -0.00562538
+ 2.51e+10Hz 0.00691974 -0.00565493
+ 2.52e+10Hz 0.00691383 -0.00568442
+ 2.53e+10Hz 0.0069079 -0.00571384
+ 2.54e+10Hz 0.00690196 -0.0057432
+ 2.55e+10Hz 0.00689601 -0.0057725
+ 2.56e+10Hz 0.00689004 -0.00580175
+ 2.57e+10Hz 0.00688407 -0.00583093
+ 2.58e+10Hz 0.00687809 -0.00586006
+ 2.59e+10Hz 0.0068721 -0.00588914
+ 2.6e+10Hz 0.00686611 -0.00591816
+ 2.61e+10Hz 0.00686011 -0.00594714
+ 2.62e+10Hz 0.0068541 -0.00597607
+ 2.63e+10Hz 0.0068481 -0.00600495
+ 2.64e+10Hz 0.00684208 -0.00603379
+ 2.65e+10Hz 0.00683607 -0.00606259
+ 2.66e+10Hz 0.00683006 -0.00609135
+ 2.67e+10Hz 0.00682404 -0.00612007
+ 2.68e+10Hz 0.00681803 -0.00614876
+ 2.69e+10Hz 0.00681201 -0.00617741
+ 2.7e+10Hz 0.006806 -0.00620604
+ 2.71e+10Hz 0.00679998 -0.00623463
+ 2.72e+10Hz 0.00679397 -0.00626319
+ 2.73e+10Hz 0.00678796 -0.00629173
+ 2.74e+10Hz 0.00678195 -0.00632025
+ 2.75e+10Hz 0.00677594 -0.00634874
+ 2.76e+10Hz 0.00676994 -0.00637721
+ 2.77e+10Hz 0.00676394 -0.00640566
+ 2.78e+10Hz 0.00675793 -0.0064341
+ 2.79e+10Hz 0.00675193 -0.00646252
+ 2.8e+10Hz 0.00674593 -0.00649093
+ 2.81e+10Hz 0.00673994 -0.00651933
+ 2.82e+10Hz 0.00673394 -0.00654773
+ 2.83e+10Hz 0.00672795 -0.00657611
+ 2.84e+10Hz 0.00672195 -0.00660449
+ 2.85e+10Hz 0.00671596 -0.00663286
+ 2.86e+10Hz 0.00670996 -0.00666123
+ 2.87e+10Hz 0.00670396 -0.0066896
+ 2.88e+10Hz 0.00669797 -0.00671798
+ 2.89e+10Hz 0.00669197 -0.00674635
+ 2.9e+10Hz 0.00668596 -0.00677473
+ 2.91e+10Hz 0.00667996 -0.00680312
+ 2.92e+10Hz 0.00667394 -0.00683151
+ 2.93e+10Hz 0.00666793 -0.00685991
+ 2.94e+10Hz 0.00666191 -0.00688833
+ 2.95e+10Hz 0.00665588 -0.00691675
+ 2.96e+10Hz 0.00664984 -0.00694519
+ 2.97e+10Hz 0.00664379 -0.00697364
+ 2.98e+10Hz 0.00663774 -0.00700211
+ 2.99e+10Hz 0.00663167 -0.00703059
+ 3e+10Hz 0.00662559 -0.0070591
+ 3.01e+10Hz 0.0066195 -0.00708762
+ 3.02e+10Hz 0.0066134 -0.00711617
+ 3.03e+10Hz 0.00660728 -0.00714473
+ 3.04e+10Hz 0.00660115 -0.00717332
+ 3.05e+10Hz 0.00659499 -0.00720193
+ 3.06e+10Hz 0.00658882 -0.00723057
+ 3.07e+10Hz 0.00658263 -0.00725924
+ 3.08e+10Hz 0.00657642 -0.00728793
+ 3.09e+10Hz 0.00657018 -0.00731664
+ 3.1e+10Hz 0.00656392 -0.00734539
+ 3.11e+10Hz 0.00655764 -0.00737417
+ 3.12e+10Hz 0.00655133 -0.00740297
+ 3.13e+10Hz 0.00654499 -0.00743181
+ 3.14e+10Hz 0.00653862 -0.00746067
+ 3.15e+10Hz 0.00653223 -0.00748957
+ 3.16e+10Hz 0.0065258 -0.00751851
+ 3.17e+10Hz 0.00651933 -0.00754747
+ 3.18e+10Hz 0.00651284 -0.00757647
+ 3.19e+10Hz 0.0065063 -0.0076055
+ 3.2e+10Hz 0.00649973 -0.00763456
+ 3.21e+10Hz 0.00649312 -0.00766366
+ 3.22e+10Hz 0.00648647 -0.0076928
+ 3.23e+10Hz 0.00647977 -0.00772197
+ 3.24e+10Hz 0.00647304 -0.00775117
+ 3.25e+10Hz 0.00646626 -0.00778041
+ 3.26e+10Hz 0.00645943 -0.00780968
+ 3.27e+10Hz 0.00645255 -0.00783899
+ 3.28e+10Hz 0.00644563 -0.00786834
+ 3.29e+10Hz 0.00643865 -0.00789772
+ 3.3e+10Hz 0.00643162 -0.00792713
+ 3.31e+10Hz 0.00642454 -0.00795658
+ 3.32e+10Hz 0.00641741 -0.00798607
+ 3.33e+10Hz 0.00641021 -0.00801559
+ 3.34e+10Hz 0.00640296 -0.00804514
+ 3.35e+10Hz 0.00639565 -0.00807473
+ 3.36e+10Hz 0.00638828 -0.00810435
+ 3.37e+10Hz 0.00638085 -0.00813401
+ 3.38e+10Hz 0.00637336 -0.0081637
+ 3.39e+10Hz 0.00636579 -0.00819342
+ 3.4e+10Hz 0.00635817 -0.00822317
+ 3.41e+10Hz 0.00635047 -0.00825296
+ 3.42e+10Hz 0.00634271 -0.00828277
+ 3.43e+10Hz 0.00633488 -0.00831262
+ 3.44e+10Hz 0.00632698 -0.00834249
+ 3.45e+10Hz 0.006319 -0.00837239
+ 3.46e+10Hz 0.00631095 -0.00840233
+ 3.47e+10Hz 0.00630283 -0.00843229
+ 3.48e+10Hz 0.00629463 -0.00846227
+ 3.49e+10Hz 0.00628635 -0.00849228
+ 3.5e+10Hz 0.006278 -0.00852232
+ 3.51e+10Hz 0.00626956 -0.00855238
+ 3.52e+10Hz 0.00626105 -0.00858247
+ 3.53e+10Hz 0.00625245 -0.00861258
+ 3.54e+10Hz 0.00624377 -0.0086427
+ 3.55e+10Hz 0.00623501 -0.00867285
+ 3.56e+10Hz 0.00622617 -0.00870302
+ 3.57e+10Hz 0.00621724 -0.00873321
+ 3.58e+10Hz 0.00620822 -0.00876341
+ 3.59e+10Hz 0.00619912 -0.00879363
+ 3.6e+10Hz 0.00618992 -0.00882387
+ 3.61e+10Hz 0.00618064 -0.00885412
+ 3.62e+10Hz 0.00617128 -0.00888438
+ 3.63e+10Hz 0.00616182 -0.00891465
+ 3.64e+10Hz 0.00615227 -0.00894494
+ 3.65e+10Hz 0.00614262 -0.00897523
+ 3.66e+10Hz 0.00613289 -0.00900553
+ 3.67e+10Hz 0.00612307 -0.00903584
+ 3.68e+10Hz 0.00611315 -0.00906616
+ 3.69e+10Hz 0.00610313 -0.00909648
+ 3.7e+10Hz 0.00609303 -0.0091268
+ 3.71e+10Hz 0.00608282 -0.00915712
+ 3.72e+10Hz 0.00607253 -0.00918745
+ 3.73e+10Hz 0.00606213 -0.00921777
+ 3.74e+10Hz 0.00605165 -0.00924809
+ 3.75e+10Hz 0.00604106 -0.00927841
+ 3.76e+10Hz 0.00603038 -0.00930872
+ 3.77e+10Hz 0.0060196 -0.00933903
+ 3.78e+10Hz 0.00600873 -0.00936933
+ 3.79e+10Hz 0.00599776 -0.00939962
+ 3.8e+10Hz 0.00598669 -0.0094299
+ 3.81e+10Hz 0.00597552 -0.00946017
+ 3.82e+10Hz 0.00596426 -0.00949043
+ 3.83e+10Hz 0.0059529 -0.00952067
+ 3.84e+10Hz 0.00594144 -0.0095509
+ 3.85e+10Hz 0.00592989 -0.00958111
+ 3.86e+10Hz 0.00591823 -0.00961131
+ 3.87e+10Hz 0.00590648 -0.00964148
+ 3.88e+10Hz 0.00589464 -0.00967163
+ 3.89e+10Hz 0.00588269 -0.00970177
+ 3.9e+10Hz 0.00587065 -0.00973187
+ 3.91e+10Hz 0.00585851 -0.00976196
+ 3.92e+10Hz 0.00584628 -0.00979201
+ 3.93e+10Hz 0.00583395 -0.00982204
+ 3.94e+10Hz 0.00582152 -0.00985205
+ 3.95e+10Hz 0.005809 -0.00988202
+ 3.96e+10Hz 0.00579639 -0.00991196
+ 3.97e+10Hz 0.00578368 -0.00994187
+ 3.98e+10Hz 0.00577088 -0.00997175
+ 3.99e+10Hz 0.00575798 -0.0100016
+ 4e+10Hz 0.00574499 -0.0100314
+ 4.01e+10Hz 0.00573191 -0.0100612
+ 4.02e+10Hz 0.00571873 -0.0100909
+ 4.03e+10Hz 0.00570547 -0.0101206
+ 4.04e+10Hz 0.00569211 -0.0101502
+ 4.05e+10Hz 0.00567866 -0.0101798
+ 4.06e+10Hz 0.00566513 -0.0102094
+ 4.07e+10Hz 0.0056515 -0.0102389
+ 4.08e+10Hz 0.00563779 -0.0102684
+ 4.09e+10Hz 0.00562399 -0.0102979
+ 4.1e+10Hz 0.00561011 -0.0103272
+ 4.11e+10Hz 0.00559614 -0.0103566
+ 4.12e+10Hz 0.00558208 -0.0103859
+ 4.13e+10Hz 0.00556794 -0.0104151
+ 4.14e+10Hz 0.00555372 -0.0104443
+ 4.15e+10Hz 0.00553941 -0.0104734
+ 4.16e+10Hz 0.00552503 -0.0105025
+ 4.17e+10Hz 0.00551056 -0.0105316
+ 4.18e+10Hz 0.00549601 -0.0105605
+ 4.19e+10Hz 0.00548139 -0.0105895
+ 4.2e+10Hz 0.00546669 -0.0106183
+ 4.21e+10Hz 0.00545191 -0.0106472
+ 4.22e+10Hz 0.00543705 -0.0106759
+ 4.23e+10Hz 0.00542212 -0.0107046
+ 4.24e+10Hz 0.00540712 -0.0107333
+ 4.25e+10Hz 0.00539205 -0.0107619
+ 4.26e+10Hz 0.0053769 -0.0107904
+ 4.27e+10Hz 0.00536168 -0.0108189
+ 4.28e+10Hz 0.0053464 -0.0108473
+ 4.29e+10Hz 0.00533104 -0.0108756
+ 4.3e+10Hz 0.00531562 -0.0109039
+ 4.31e+10Hz 0.00530013 -0.0109321
+ 4.32e+10Hz 0.00528458 -0.0109603
+ 4.33e+10Hz 0.00526896 -0.0109884
+ 4.34e+10Hz 0.00525328 -0.0110164
+ 4.35e+10Hz 0.00523754 -0.0110444
+ 4.36e+10Hz 0.00522174 -0.0110723
+ 4.37e+10Hz 0.00520587 -0.0111001
+ 4.38e+10Hz 0.00518995 -0.0111279
+ 4.39e+10Hz 0.00517397 -0.0111556
+ 4.4e+10Hz 0.00515794 -0.0111833
+ 4.41e+10Hz 0.00514185 -0.0112109
+ 4.42e+10Hz 0.0051257 -0.0112384
+ 4.43e+10Hz 0.00510951 -0.0112659
+ 4.44e+10Hz 0.00509326 -0.0112933
+ 4.45e+10Hz 0.00507696 -0.0113206
+ 4.46e+10Hz 0.00506061 -0.0113479
+ 4.47e+10Hz 0.00504421 -0.0113751
+ 4.48e+10Hz 0.00502776 -0.0114022
+ 4.49e+10Hz 0.00501127 -0.0114293
+ 4.5e+10Hz 0.00499473 -0.0114563
+ 4.51e+10Hz 0.00497815 -0.0114833
+ 4.52e+10Hz 0.00496152 -0.0115102
+ 4.53e+10Hz 0.00494485 -0.011537
+ 4.54e+10Hz 0.00492814 -0.0115637
+ 4.55e+10Hz 0.00491139 -0.0115904
+ 4.56e+10Hz 0.0048946 -0.0116171
+ 4.57e+10Hz 0.00487777 -0.0116436
+ 4.58e+10Hz 0.00486091 -0.0116701
+ 4.59e+10Hz 0.004844 -0.0116966
+ 4.6e+10Hz 0.00482706 -0.0117229
+ 4.61e+10Hz 0.00481009 -0.0117493
+ 4.62e+10Hz 0.00479308 -0.0117755
+ 4.63e+10Hz 0.00477604 -0.0118017
+ 4.64e+10Hz 0.00475897 -0.0118279
+ 4.65e+10Hz 0.00474187 -0.0118539
+ 4.66e+10Hz 0.00472473 -0.01188
+ 4.67e+10Hz 0.00470757 -0.0119059
+ 4.68e+10Hz 0.00469037 -0.0119318
+ 4.69e+10Hz 0.00467315 -0.0119577
+ 4.7e+10Hz 0.0046559 -0.0119834
+ 4.71e+10Hz 0.00463863 -0.0120092
+ 4.72e+10Hz 0.00462133 -0.0120349
+ 4.73e+10Hz 0.004604 -0.0120605
+ 4.74e+10Hz 0.00458665 -0.012086
+ 4.75e+10Hz 0.00456928 -0.0121115
+ 4.76e+10Hz 0.00455188 -0.012137
+ 4.77e+10Hz 0.00453446 -0.0121624
+ 4.78e+10Hz 0.00451701 -0.0121878
+ 4.79e+10Hz 0.00449955 -0.0122131
+ 4.8e+10Hz 0.00448206 -0.0122383
+ 4.81e+10Hz 0.00446456 -0.0122635
+ 4.82e+10Hz 0.00444703 -0.0122887
+ 4.83e+10Hz 0.00442948 -0.0123138
+ 4.84e+10Hz 0.00441192 -0.0123388
+ 4.85e+10Hz 0.00439433 -0.0123638
+ 4.86e+10Hz 0.00437673 -0.0123888
+ 4.87e+10Hz 0.00435911 -0.0124137
+ 4.88e+10Hz 0.00434147 -0.0124386
+ 4.89e+10Hz 0.00432381 -0.0124634
+ 4.9e+10Hz 0.00430614 -0.0124882
+ 4.91e+10Hz 0.00428845 -0.0125129
+ 4.92e+10Hz 0.00427074 -0.0125376
+ 4.93e+10Hz 0.00425302 -0.0125623
+ 4.94e+10Hz 0.00423528 -0.0125869
+ 4.95e+10Hz 0.00421752 -0.0126114
+ 4.96e+10Hz 0.00419975 -0.012636
+ 4.97e+10Hz 0.00418197 -0.0126605
+ 4.98e+10Hz 0.00416416 -0.0126849
+ 4.99e+10Hz 0.00414634 -0.0127094
+ 5e+10Hz 0.00412851 -0.0127337
+ 5.01e+10Hz 0.00411066 -0.0127581
+ 5.02e+10Hz 0.00409279 -0.0127824
+ 5.03e+10Hz 0.00407491 -0.0128067
+ 5.04e+10Hz 0.00405702 -0.0128309
+ 5.05e+10Hz 0.00403911 -0.0128552
+ 5.06e+10Hz 0.00402118 -0.0128793
+ 5.07e+10Hz 0.00400323 -0.0129035
+ 5.08e+10Hz 0.00398527 -0.0129276
+ 5.09e+10Hz 0.0039673 -0.0129517
+ 5.1e+10Hz 0.0039493 -0.0129758
+ 5.11e+10Hz 0.00393129 -0.0129998
+ 5.12e+10Hz 0.00391327 -0.0130238
+ 5.13e+10Hz 0.00389523 -0.0130478
+ 5.14e+10Hz 0.00387717 -0.0130718
+ 5.15e+10Hz 0.00385909 -0.0130957
+ 5.16e+10Hz 0.00384099 -0.0131196
+ 5.17e+10Hz 0.00382288 -0.0131435
+ 5.18e+10Hz 0.00380475 -0.0131673
+ 5.19e+10Hz 0.00378659 -0.0131912
+ 5.2e+10Hz 0.00376842 -0.013215
+ 5.21e+10Hz 0.00375023 -0.0132388
+ 5.22e+10Hz 0.00373202 -0.0132625
+ 5.23e+10Hz 0.00371379 -0.0132863
+ 5.24e+10Hz 0.00369554 -0.01331
+ 5.25e+10Hz 0.00367727 -0.0133337
+ 5.26e+10Hz 0.00365898 -0.0133574
+ 5.27e+10Hz 0.00364066 -0.013381
+ 5.28e+10Hz 0.00362232 -0.0134047
+ 5.29e+10Hz 0.00360396 -0.0134283
+ 5.3e+10Hz 0.00358558 -0.0134519
+ 5.31e+10Hz 0.00356717 -0.0134755
+ 5.32e+10Hz 0.00354873 -0.0134991
+ 5.33e+10Hz 0.00353027 -0.0135226
+ 5.34e+10Hz 0.00351179 -0.0135462
+ 5.35e+10Hz 0.00349328 -0.0135697
+ 5.36e+10Hz 0.00347474 -0.0135932
+ 5.37e+10Hz 0.00345617 -0.0136167
+ 5.38e+10Hz 0.00343758 -0.0136402
+ 5.39e+10Hz 0.00341896 -0.0136636
+ 5.4e+10Hz 0.00340031 -0.0136871
+ 5.41e+10Hz 0.00338162 -0.0137105
+ 5.42e+10Hz 0.00336291 -0.0137339
+ 5.43e+10Hz 0.00334417 -0.0137573
+ 5.44e+10Hz 0.0033254 -0.0137807
+ 5.45e+10Hz 0.00330659 -0.0138041
+ 5.46e+10Hz 0.00328775 -0.0138274
+ 5.47e+10Hz 0.00326888 -0.0138507
+ 5.48e+10Hz 0.00324997 -0.0138741
+ 5.49e+10Hz 0.00323103 -0.0138974
+ 5.5e+10Hz 0.00321206 -0.0139207
+ 5.51e+10Hz 0.00319305 -0.013944
+ 5.52e+10Hz 0.003174 -0.0139672
+ 5.53e+10Hz 0.00315491 -0.0139905
+ 5.54e+10Hz 0.00313579 -0.0140137
+ 5.55e+10Hz 0.00311663 -0.0140369
+ 5.56e+10Hz 0.00309743 -0.0140601
+ 5.57e+10Hz 0.00307819 -0.0140833
+ 5.58e+10Hz 0.00305891 -0.0141065
+ 5.59e+10Hz 0.00303959 -0.0141296
+ 5.6e+10Hz 0.00302023 -0.0141528
+ 5.61e+10Hz 0.00300083 -0.0141759
+ 5.62e+10Hz 0.00298138 -0.014199
+ 5.63e+10Hz 0.0029619 -0.0142221
+ 5.64e+10Hz 0.00294236 -0.0142452
+ 5.65e+10Hz 0.00292279 -0.0142682
+ 5.66e+10Hz 0.00290317 -0.0142913
+ 5.67e+10Hz 0.0028835 -0.0143143
+ 5.68e+10Hz 0.00286379 -0.0143373
+ 5.69e+10Hz 0.00284404 -0.0143603
+ 5.7e+10Hz 0.00282424 -0.0143832
+ 5.71e+10Hz 0.00280439 -0.0144062
+ 5.72e+10Hz 0.00278449 -0.0144291
+ 5.73e+10Hz 0.00276454 -0.014452
+ 5.74e+10Hz 0.00274455 -0.0144749
+ 5.75e+10Hz 0.00272451 -0.0144978
+ 5.76e+10Hz 0.00270442 -0.0145206
+ 5.77e+10Hz 0.00268427 -0.0145434
+ 5.78e+10Hz 0.00266408 -0.0145662
+ 5.79e+10Hz 0.00264384 -0.014589
+ 5.8e+10Hz 0.00262355 -0.0146117
+ 5.81e+10Hz 0.0026032 -0.0146345
+ 5.82e+10Hz 0.00258281 -0.0146571
+ 5.83e+10Hz 0.00256236 -0.0146798
+ 5.84e+10Hz 0.00254186 -0.0147025
+ 5.85e+10Hz 0.00252131 -0.0147251
+ 5.86e+10Hz 0.00250071 -0.0147477
+ 5.87e+10Hz 0.00248005 -0.0147702
+ 5.88e+10Hz 0.00245934 -0.0147928
+ 5.89e+10Hz 0.00243858 -0.0148153
+ 5.9e+10Hz 0.00241776 -0.0148378
+ 5.91e+10Hz 0.00239689 -0.0148602
+ 5.92e+10Hz 0.00237597 -0.0148826
+ 5.93e+10Hz 0.00235499 -0.014905
+ 5.94e+10Hz 0.00233395 -0.0149274
+ 5.95e+10Hz 0.00231287 -0.0149497
+ 5.96e+10Hz 0.00229172 -0.014972
+ 5.97e+10Hz 0.00227053 -0.0149942
+ 5.98e+10Hz 0.00224928 -0.0150164
+ 5.99e+10Hz 0.00222797 -0.0150386
+ 6e+10Hz 0.00220661 -0.0150607
+ 6.01e+10Hz 0.0021852 -0.0150829
+ 6.02e+10Hz 0.00216373 -0.0151049
+ 6.03e+10Hz 0.0021422 -0.015127
+ 6.04e+10Hz 0.00212063 -0.0151489
+ 6.05e+10Hz 0.00209899 -0.0151709
+ 6.06e+10Hz 0.00207731 -0.0151928
+ 6.07e+10Hz 0.00205556 -0.0152147
+ 6.08e+10Hz 0.00203377 -0.0152365
+ 6.09e+10Hz 0.00201192 -0.0152583
+ 6.1e+10Hz 0.00199002 -0.01528
+ 6.11e+10Hz 0.00196806 -0.0153017
+ 6.12e+10Hz 0.00194605 -0.0153234
+ 6.13e+10Hz 0.00192398 -0.015345
+ 6.14e+10Hz 0.00190187 -0.0153665
+ 6.15e+10Hz 0.0018797 -0.015388
+ 6.16e+10Hz 0.00185747 -0.0154095
+ 6.17e+10Hz 0.0018352 -0.0154309
+ 6.18e+10Hz 0.00181287 -0.0154523
+ 6.19e+10Hz 0.00179049 -0.0154736
+ 6.2e+10Hz 0.00176806 -0.0154949
+ 6.21e+10Hz 0.00174558 -0.0155161
+ 6.22e+10Hz 0.00172305 -0.0155373
+ 6.23e+10Hz 0.00170047 -0.0155584
+ 6.24e+10Hz 0.00167783 -0.0155795
+ 6.25e+10Hz 0.00165515 -0.0156005
+ 6.26e+10Hz 0.00163242 -0.0156214
+ 6.27e+10Hz 0.00160964 -0.0156423
+ 6.28e+10Hz 0.00158682 -0.0156632
+ 6.29e+10Hz 0.00156394 -0.015684
+ 6.3e+10Hz 0.00154102 -0.0157047
+ 6.31e+10Hz 0.00151805 -0.0157254
+ 6.32e+10Hz 0.00149503 -0.015746
+ 6.33e+10Hz 0.00147197 -0.0157666
+ 6.34e+10Hz 0.00144886 -0.0157871
+ 6.35e+10Hz 0.00142571 -0.0158076
+ 6.36e+10Hz 0.00140252 -0.015828
+ 6.37e+10Hz 0.00137928 -0.0158483
+ 6.38e+10Hz 0.001356 -0.0158686
+ 6.39e+10Hz 0.00133267 -0.0158888
+ 6.4e+10Hz 0.0013093 -0.015909
+ 6.41e+10Hz 0.0012859 -0.0159291
+ 6.42e+10Hz 0.00126245 -0.0159491
+ 6.43e+10Hz 0.00123896 -0.0159691
+ 6.44e+10Hz 0.00121543 -0.015989
+ 6.45e+10Hz 0.00119186 -0.0160089
+ 6.46e+10Hz 0.00116826 -0.0160287
+ 6.47e+10Hz 0.00114461 -0.0160484
+ 6.48e+10Hz 0.00112093 -0.016068
+ 6.49e+10Hz 0.00109722 -0.0160876
+ 6.5e+10Hz 0.00107346 -0.0161072
+ 6.51e+10Hz 0.00104968 -0.0161267
+ 6.52e+10Hz 0.00102586 -0.0161461
+ 6.53e+10Hz 0.001002 -0.0161654
+ 6.54e+10Hz 0.000978114 -0.0161847
+ 6.55e+10Hz 0.000954194 -0.0162039
+ 6.56e+10Hz 0.000930242 -0.0162231
+ 6.57e+10Hz 0.000906259 -0.0162422
+ 6.58e+10Hz 0.000882246 -0.0162612
+ 6.59e+10Hz 0.000858204 -0.0162802
+ 6.6e+10Hz 0.000834133 -0.0162991
+ 6.61e+10Hz 0.000810033 -0.0163179
+ 6.62e+10Hz 0.000785906 -0.0163367
+ 6.63e+10Hz 0.000761752 -0.0163554
+ 6.64e+10Hz 0.000737572 -0.016374
+ 6.65e+10Hz 0.000713366 -0.0163926
+ 6.66e+10Hz 0.000689136 -0.0164111
+ 6.67e+10Hz 0.000664881 -0.0164295
+ 6.68e+10Hz 0.000640603 -0.0164479
+ 6.69e+10Hz 0.000616302 -0.0164662
+ 6.7e+10Hz 0.000591979 -0.0164845
+ 6.71e+10Hz 0.000567634 -0.0165026
+ 6.72e+10Hz 0.000543269 -0.0165208
+ 6.73e+10Hz 0.000518883 -0.0165388
+ 6.74e+10Hz 0.000494478 -0.0165568
+ 6.75e+10Hz 0.000470054 -0.0165747
+ 6.76e+10Hz 0.000445611 -0.0165926
+ 6.77e+10Hz 0.000421151 -0.0166104
+ 6.78e+10Hz 0.000396674 -0.0166281
+ 6.79e+10Hz 0.00037218 -0.0166458
+ 6.8e+10Hz 0.00034767 -0.0166634
+ 6.81e+10Hz 0.000323145 -0.016681
+ 6.82e+10Hz 0.000298606 -0.0166985
+ 6.83e+10Hz 0.000274052 -0.0167159
+ 6.84e+10Hz 0.000249484 -0.0167332
+ 6.85e+10Hz 0.000224904 -0.0167505
+ 6.86e+10Hz 0.00020031 -0.0167678
+ 6.87e+10Hz 0.000175705 -0.016785
+ 6.88e+10Hz 0.000151089 -0.0168021
+ 6.89e+10Hz 0.000126461 -0.0168191
+ 6.9e+10Hz 0.000101823 -0.0168361
+ 6.91e+10Hz 7.71752e-05 -0.0168531
+ 6.92e+10Hz 5.25176e-05 -0.01687
+ 6.93e+10Hz 2.7851e-05 -0.0168868
+ 6.94e+10Hz 3.17567e-06 -0.0169035
+ 6.95e+10Hz -2.15078e-05 -0.0169202
+ 6.96e+10Hz -4.61991e-05 -0.0169369
+ 6.97e+10Hz -7.08978e-05 -0.0169535
+ 6.98e+10Hz -9.56035e-05 -0.01697
+ 6.99e+10Hz -0.000120316 -0.0169865
+ 7e+10Hz -0.000145034 -0.0170029
+ 7.01e+10Hz -0.000169759 -0.0170193
+ 7.02e+10Hz -0.000194489 -0.0170356
+ 7.03e+10Hz -0.000219224 -0.0170519
+ 7.04e+10Hz -0.000243964 -0.0170681
+ 7.05e+10Hz -0.000268709 -0.0170842
+ 7.06e+10Hz -0.000293458 -0.0171003
+ 7.07e+10Hz -0.000318212 -0.0171163
+ 7.08e+10Hz -0.000342969 -0.0171323
+ 7.09e+10Hz -0.00036773 -0.0171483
+ 7.1e+10Hz -0.000392494 -0.0171642
+ 7.11e+10Hz -0.000417262 -0.01718
+ 7.12e+10Hz -0.000442032 -0.0171958
+ 7.13e+10Hz -0.000466806 -0.0172116
+ 7.14e+10Hz -0.000491582 -0.0172272
+ 7.15e+10Hz -0.000516361 -0.0172429
+ 7.16e+10Hz -0.000541142 -0.0172585
+ 7.17e+10Hz -0.000565925 -0.017274
+ 7.18e+10Hz -0.000590711 -0.0172895
+ 7.19e+10Hz -0.000615499 -0.017305
+ 7.2e+10Hz -0.000640289 -0.0173204
+ 7.21e+10Hz -0.000665081 -0.0173358
+ 7.22e+10Hz -0.000689875 -0.0173511
+ 7.23e+10Hz -0.000714671 -0.0173664
+ 7.24e+10Hz -0.000739469 -0.0173816
+ 7.25e+10Hz -0.000764269 -0.0173968
+ 7.26e+10Hz -0.000789071 -0.0174119
+ 7.27e+10Hz -0.000813875 -0.017427
+ 7.28e+10Hz -0.000838681 -0.0174421
+ 7.29e+10Hz -0.00086349 -0.0174571
+ 7.3e+10Hz -0.0008883 -0.0174721
+ 7.31e+10Hz -0.000913113 -0.017487
+ 7.32e+10Hz -0.000937929 -0.0175019
+ 7.33e+10Hz -0.000962747 -0.0175168
+ 7.34e+10Hz -0.000987567 -0.0175316
+ 7.35e+10Hz -0.00101239 -0.0175464
+ 7.36e+10Hz -0.00103722 -0.0175611
+ 7.37e+10Hz -0.00106205 -0.0175758
+ 7.38e+10Hz -0.00108688 -0.0175905
+ 7.39e+10Hz -0.00111172 -0.0176051
+ 7.4e+10Hz -0.00113656 -0.0176197
+ 7.41e+10Hz -0.0011614 -0.0176343
+ 7.42e+10Hz -0.00118625 -0.0176488
+ 7.43e+10Hz -0.0012111 -0.0176633
+ 7.44e+10Hz -0.00123596 -0.0176778
+ 7.45e+10Hz -0.00126082 -0.0176922
+ 7.46e+10Hz -0.00128569 -0.0177066
+ 7.47e+10Hz -0.00131056 -0.0177209
+ 7.48e+10Hz -0.00133544 -0.0177352
+ 7.49e+10Hz -0.00136033 -0.0177495
+ 7.5e+10Hz -0.00138522 -0.0177638
+ 7.51e+10Hz -0.00141012 -0.017778
+ 7.52e+10Hz -0.00143503 -0.0177921
+ 7.53e+10Hz -0.00145994 -0.0178063
+ 7.54e+10Hz -0.00148486 -0.0178204
+ 7.55e+10Hz -0.00150979 -0.0178345
+ 7.56e+10Hz -0.00153472 -0.0178486
+ 7.57e+10Hz -0.00155967 -0.0178626
+ 7.58e+10Hz -0.00158463 -0.0178766
+ 7.59e+10Hz -0.00160959 -0.0178905
+ 7.6e+10Hz -0.00163456 -0.0179045
+ 7.61e+10Hz -0.00165955 -0.0179184
+ 7.62e+10Hz -0.00168454 -0.0179322
+ 7.63e+10Hz -0.00170955 -0.0179461
+ 7.64e+10Hz -0.00173457 -0.0179599
+ 7.65e+10Hz -0.0017596 -0.0179737
+ 7.66e+10Hz -0.00178464 -0.0179874
+ 7.67e+10Hz -0.00180969 -0.0180011
+ 7.68e+10Hz -0.00183476 -0.0180148
+ 7.69e+10Hz -0.00185984 -0.0180285
+ 7.7e+10Hz -0.00188493 -0.0180421
+ 7.71e+10Hz -0.00191004 -0.0180557
+ 7.72e+10Hz -0.00193516 -0.0180693
+ 7.73e+10Hz -0.0019603 -0.0180828
+ 7.74e+10Hz -0.00198546 -0.0180963
+ 7.75e+10Hz -0.00201062 -0.0181098
+ 7.76e+10Hz -0.00203581 -0.0181232
+ 7.77e+10Hz -0.00206101 -0.0181366
+ 7.78e+10Hz -0.00208623 -0.01815
+ 7.79e+10Hz -0.00211147 -0.0181634
+ 7.8e+10Hz -0.00213672 -0.0181767
+ 7.81e+10Hz -0.00216199 -0.01819
+ 7.82e+10Hz -0.00218728 -0.0182033
+ 7.83e+10Hz -0.00221259 -0.0182165
+ 7.84e+10Hz -0.00223792 -0.0182297
+ 7.85e+10Hz -0.00226327 -0.0182429
+ 7.86e+10Hz -0.00228864 -0.018256
+ 7.87e+10Hz -0.00231403 -0.0182691
+ 7.88e+10Hz -0.00233944 -0.0182822
+ 7.89e+10Hz -0.00236487 -0.0182952
+ 7.9e+10Hz -0.00239032 -0.0183083
+ 7.91e+10Hz -0.0024158 -0.0183212
+ 7.92e+10Hz -0.00244129 -0.0183342
+ 7.93e+10Hz -0.00246681 -0.0183471
+ 7.94e+10Hz -0.00249235 -0.01836
+ 7.95e+10Hz -0.00251792 -0.0183728
+ 7.96e+10Hz -0.00254351 -0.0183856
+ 7.97e+10Hz -0.00256912 -0.0183984
+ 7.98e+10Hz -0.00259475 -0.0184112
+ 7.99e+10Hz -0.00262041 -0.0184239
+ 8e+10Hz -0.0026461 -0.0184366
+ 8.01e+10Hz -0.00267181 -0.0184492
+ 8.02e+10Hz -0.00269754 -0.0184618
+ 8.03e+10Hz -0.0027233 -0.0184744
+ 8.04e+10Hz -0.00274908 -0.0184869
+ 8.05e+10Hz -0.00277489 -0.0184994
+ 8.06e+10Hz -0.00280073 -0.0185119
+ 8.07e+10Hz -0.00282659 -0.0185243
+ 8.08e+10Hz -0.00285248 -0.0185367
+ 8.09e+10Hz -0.0028784 -0.018549
+ 8.1e+10Hz -0.00290434 -0.0185613
+ 8.11e+10Hz -0.00293031 -0.0185736
+ 8.12e+10Hz -0.0029563 -0.0185858
+ 8.13e+10Hz -0.00298233 -0.018598
+ 8.14e+10Hz -0.00300838 -0.0186101
+ 8.15e+10Hz -0.00303445 -0.0186222
+ 8.16e+10Hz -0.00306056 -0.0186343
+ 8.17e+10Hz -0.00308669 -0.0186463
+ 8.18e+10Hz -0.00311285 -0.0186583
+ 8.19e+10Hz -0.00313904 -0.0186702
+ 8.2e+10Hz -0.00316525 -0.0186821
+ 8.21e+10Hz -0.00319149 -0.018694
+ 8.22e+10Hz -0.00321776 -0.0187058
+ 8.23e+10Hz -0.00324406 -0.0187175
+ 8.24e+10Hz -0.00327039 -0.0187293
+ 8.25e+10Hz -0.00329674 -0.0187409
+ 8.26e+10Hz -0.00332312 -0.0187525
+ 8.27e+10Hz -0.00334953 -0.0187641
+ 8.28e+10Hz -0.00337596 -0.0187756
+ 8.29e+10Hz -0.00340242 -0.0187871
+ 8.3e+10Hz -0.00342892 -0.0187986
+ 8.31e+10Hz -0.00345543 -0.0188099
+ 8.32e+10Hz -0.00348198 -0.0188213
+ 8.33e+10Hz -0.00350855 -0.0188326
+ 8.34e+10Hz -0.00353515 -0.0188438
+ 8.35e+10Hz -0.00356177 -0.018855
+ 8.36e+10Hz -0.00358843 -0.0188661
+ 8.37e+10Hz -0.0036151 -0.0188772
+ 8.38e+10Hz -0.00364181 -0.0188882
+ 8.39e+10Hz -0.00366854 -0.0188992
+ 8.4e+10Hz -0.0036953 -0.0189101
+ 8.41e+10Hz -0.00372208 -0.018921
+ 8.42e+10Hz -0.00374888 -0.0189318
+ 8.43e+10Hz -0.00377572 -0.0189426
+ 8.44e+10Hz -0.00380258 -0.0189533
+ 8.45e+10Hz -0.00382946 -0.0189639
+ 8.46e+10Hz -0.00385636 -0.0189745
+ 8.47e+10Hz -0.00388329 -0.0189851
+ 8.48e+10Hz -0.00391025 -0.0189956
+ 8.49e+10Hz -0.00393723 -0.019006
+ 8.5e+10Hz -0.00396423 -0.0190164
+ 8.51e+10Hz -0.00399125 -0.0190267
+ 8.52e+10Hz -0.0040183 -0.0190369
+ 8.53e+10Hz -0.00404537 -0.0190471
+ 8.54e+10Hz -0.00407246 -0.0190573
+ 8.55e+10Hz -0.00409957 -0.0190674
+ 8.56e+10Hz -0.0041267 -0.0190774
+ 8.57e+10Hz -0.00415385 -0.0190873
+ 8.58e+10Hz -0.00418103 -0.0190972
+ 8.59e+10Hz -0.00420822 -0.0191071
+ 8.6e+10Hz -0.00423543 -0.0191168
+ 8.61e+10Hz -0.00426266 -0.0191266
+ 8.62e+10Hz -0.00428991 -0.0191362
+ 8.63e+10Hz -0.00431718 -0.0191458
+ 8.64e+10Hz -0.00434447 -0.0191554
+ 8.65e+10Hz -0.00437177 -0.0191648
+ 8.66e+10Hz -0.00439909 -0.0191742
+ 8.67e+10Hz -0.00442643 -0.0191836
+ 8.68e+10Hz -0.00445378 -0.0191929
+ 8.69e+10Hz -0.00448115 -0.0192021
+ 8.7e+10Hz -0.00450853 -0.0192112
+ 8.71e+10Hz -0.00453593 -0.0192203
+ 8.72e+10Hz -0.00456334 -0.0192293
+ 8.73e+10Hz -0.00459076 -0.0192383
+ 8.74e+10Hz -0.0046182 -0.0192472
+ 8.75e+10Hz -0.00464565 -0.019256
+ 8.76e+10Hz -0.00467311 -0.0192648
+ 8.77e+10Hz -0.00470059 -0.0192735
+ 8.78e+10Hz -0.00472807 -0.0192822
+ 8.79e+10Hz -0.00475556 -0.0192907
+ 8.8e+10Hz -0.00478307 -0.0192992
+ 8.81e+10Hz -0.00481058 -0.0193077
+ 8.82e+10Hz -0.00483811 -0.0193161
+ 8.83e+10Hz -0.00486564 -0.0193244
+ 8.84e+10Hz -0.00489318 -0.0193326
+ 8.85e+10Hz -0.00492072 -0.0193408
+ 8.86e+10Hz -0.00494828 -0.0193489
+ 8.87e+10Hz -0.00497583 -0.019357
+ 8.88e+10Hz -0.0050034 -0.0193649
+ 8.89e+10Hz -0.00503097 -0.0193729
+ 8.9e+10Hz -0.00505855 -0.0193807
+ 8.91e+10Hz -0.00508613 -0.0193885
+ 8.92e+10Hz -0.00511371 -0.0193962
+ 8.93e+10Hz -0.0051413 -0.0194039
+ 8.94e+10Hz -0.00516888 -0.0194115
+ 8.95e+10Hz -0.00519648 -0.019419
+ 8.96e+10Hz -0.00522407 -0.0194265
+ 8.97e+10Hz -0.00525166 -0.0194338
+ 8.98e+10Hz -0.00527926 -0.0194412
+ 8.99e+10Hz -0.00530685 -0.0194484
+ 9e+10Hz -0.00533445 -0.0194556
+ 9.01e+10Hz -0.00536204 -0.0194628
+ 9.02e+10Hz -0.00538963 -0.0194698
+ 9.03e+10Hz -0.00541723 -0.0194768
+ 9.04e+10Hz -0.00544481 -0.0194838
+ 9.05e+10Hz -0.0054724 -0.0194907
+ 9.06e+10Hz -0.00549998 -0.0194975
+ 9.07e+10Hz -0.00552756 -0.0195042
+ 9.08e+10Hz -0.00555514 -0.0195109
+ 9.09e+10Hz -0.00558271 -0.0195175
+ 9.1e+10Hz -0.00561028 -0.0195241
+ 9.11e+10Hz -0.00563784 -0.0195306
+ 9.12e+10Hz -0.00566539 -0.019537
+ 9.13e+10Hz -0.00569294 -0.0195433
+ 9.14e+10Hz -0.00572048 -0.0195497
+ 9.15e+10Hz -0.00574802 -0.0195559
+ 9.16e+10Hz -0.00577554 -0.0195621
+ 9.17e+10Hz -0.00580306 -0.0195682
+ 9.18e+10Hz -0.00583058 -0.0195742
+ 9.19e+10Hz -0.00585808 -0.0195802
+ 9.2e+10Hz -0.00588557 -0.0195862
+ 9.21e+10Hz -0.00591306 -0.019592
+ 9.22e+10Hz -0.00594053 -0.0195979
+ 9.23e+10Hz -0.005968 -0.0196036
+ 9.24e+10Hz -0.00599545 -0.0196093
+ 9.25e+10Hz -0.0060229 -0.0196149
+ 9.26e+10Hz -0.00605033 -0.0196205
+ 9.27e+10Hz -0.00607776 -0.019626
+ 9.28e+10Hz -0.00610517 -0.0196315
+ 9.29e+10Hz -0.00613257 -0.0196369
+ 9.3e+10Hz -0.00615996 -0.0196422
+ 9.31e+10Hz -0.00618733 -0.0196475
+ 9.32e+10Hz -0.0062147 -0.0196527
+ 9.33e+10Hz -0.00624205 -0.0196579
+ 9.34e+10Hz -0.00626938 -0.019663
+ 9.35e+10Hz -0.00629671 -0.0196681
+ 9.36e+10Hz -0.00632402 -0.0196731
+ 9.37e+10Hz -0.00635132 -0.019678
+ 9.38e+10Hz -0.0063786 -0.0196829
+ 9.39e+10Hz -0.00640587 -0.0196877
+ 9.4e+10Hz -0.00643313 -0.0196925
+ 9.41e+10Hz -0.00646037 -0.0196972
+ 9.42e+10Hz -0.0064876 -0.0197019
+ 9.43e+10Hz -0.00651481 -0.0197065
+ 9.44e+10Hz -0.00654201 -0.0197111
+ 9.45e+10Hz -0.00656919 -0.0197156
+ 9.46e+10Hz -0.00659636 -0.0197201
+ 9.47e+10Hz -0.00662351 -0.0197245
+ 9.48e+10Hz -0.00665065 -0.0197288
+ 9.49e+10Hz -0.00667778 -0.0197331
+ 9.5e+10Hz -0.00670488 -0.0197374
+ 9.51e+10Hz -0.00673198 -0.0197416
+ 9.52e+10Hz -0.00675905 -0.0197457
+ 9.53e+10Hz -0.00678612 -0.0197499
+ 9.54e+10Hz -0.00681316 -0.0197539
+ 9.55e+10Hz -0.0068402 -0.0197579
+ 9.56e+10Hz -0.00686721 -0.0197619
+ 9.57e+10Hz -0.00689421 -0.0197658
+ 9.58e+10Hz -0.0069212 -0.0197696
+ 9.59e+10Hz -0.00694817 -0.0197734
+ 9.6e+10Hz -0.00697512 -0.0197772
+ 9.61e+10Hz -0.00700206 -0.0197809
+ 9.62e+10Hz -0.00702899 -0.0197846
+ 9.63e+10Hz -0.00705589 -0.0197882
+ 9.64e+10Hz -0.00708279 -0.0197918
+ 9.65e+10Hz -0.00710967 -0.0197953
+ 9.66e+10Hz -0.00713653 -0.0197988
+ 9.67e+10Hz -0.00716338 -0.0198023
+ 9.68e+10Hz -0.00719021 -0.0198056
+ 9.69e+10Hz -0.00721703 -0.019809
+ 9.7e+10Hz -0.00724383 -0.0198123
+ 9.71e+10Hz -0.00727062 -0.0198156
+ 9.72e+10Hz -0.0072974 -0.0198188
+ 9.73e+10Hz -0.00732416 -0.0198219
+ 9.74e+10Hz -0.0073509 -0.0198251
+ 9.75e+10Hz -0.00737763 -0.0198281
+ 9.76e+10Hz -0.00740435 -0.0198312
+ 9.77e+10Hz -0.00743105 -0.0198342
+ 9.78e+10Hz -0.00745774 -0.0198371
+ 9.79e+10Hz -0.00748442 -0.01984
+ 9.8e+10Hz -0.00751108 -0.0198429
+ 9.81e+10Hz -0.00753773 -0.0198457
+ 9.82e+10Hz -0.00756437 -0.0198485
+ 9.83e+10Hz -0.00759099 -0.0198513
+ 9.84e+10Hz -0.0076176 -0.0198539
+ 9.85e+10Hz -0.0076442 -0.0198566
+ 9.86e+10Hz -0.00767078 -0.0198592
+ 9.87e+10Hz -0.00769736 -0.0198618
+ 9.88e+10Hz -0.00772392 -0.0198643
+ 9.89e+10Hz -0.00775047 -0.0198668
+ 9.9e+10Hz -0.007777 -0.0198693
+ 9.91e+10Hz -0.00780353 -0.0198717
+ 9.92e+10Hz -0.00783004 -0.019874
+ 9.93e+10Hz -0.00785654 -0.0198763
+ 9.94e+10Hz -0.00788303 -0.0198786
+ 9.95e+10Hz -0.00790951 -0.0198809
+ 9.96e+10Hz -0.00793598 -0.0198831
+ 9.97e+10Hz -0.00796244 -0.0198852
+ 9.98e+10Hz -0.00798889 -0.0198873
+ 9.99e+10Hz -0.00801533 -0.0198894
+ 1e+11Hz -0.00804175 -0.0198914
+ 1.001e+11Hz -0.00806817 -0.0198934
+ 1.002e+11Hz -0.00809458 -0.0198954
+ 1.003e+11Hz -0.00812098 -0.0198973
+ 1.004e+11Hz -0.00814737 -0.0198992
+ 1.005e+11Hz -0.00817375 -0.019901
+ 1.006e+11Hz -0.00820012 -0.0199028
+ 1.007e+11Hz -0.00822648 -0.0199045
+ 1.008e+11Hz -0.00825283 -0.0199063
+ 1.009e+11Hz -0.00827917 -0.0199079
+ 1.01e+11Hz -0.00830551 -0.0199095
+ 1.011e+11Hz -0.00833184 -0.0199111
+ 1.012e+11Hz -0.00835816 -0.0199127
+ 1.013e+11Hz -0.00838447 -0.0199142
+ 1.014e+11Hz -0.00841077 -0.0199156
+ 1.015e+11Hz -0.00843707 -0.019917
+ 1.016e+11Hz -0.00846336 -0.0199184
+ 1.017e+11Hz -0.00848964 -0.0199197
+ 1.018e+11Hz -0.00851591 -0.019921
+ 1.019e+11Hz -0.00854217 -0.0199223
+ 1.02e+11Hz -0.00856843 -0.0199235
+ 1.021e+11Hz -0.00859468 -0.0199246
+ 1.022e+11Hz -0.00862093 -0.0199257
+ 1.023e+11Hz -0.00864717 -0.0199268
+ 1.024e+11Hz -0.0086734 -0.0199278
+ 1.025e+11Hz -0.00869962 -0.0199288
+ 1.026e+11Hz -0.00872584 -0.0199298
+ 1.027e+11Hz -0.00875205 -0.0199307
+ 1.028e+11Hz -0.00877825 -0.0199315
+ 1.029e+11Hz -0.00880445 -0.0199323
+ 1.03e+11Hz -0.00883064 -0.0199331
+ 1.031e+11Hz -0.00885682 -0.0199338
+ 1.032e+11Hz -0.008883 -0.0199345
+ 1.033e+11Hz -0.00890917 -0.0199351
+ 1.034e+11Hz -0.00893534 -0.0199357
+ 1.035e+11Hz -0.00896149 -0.0199363
+ 1.036e+11Hz -0.00898764 -0.0199368
+ 1.037e+11Hz -0.00901379 -0.0199372
+ 1.038e+11Hz -0.00903993 -0.0199376
+ 1.039e+11Hz -0.00906606 -0.019938
+ 1.04e+11Hz -0.00909218 -0.0199383
+ 1.041e+11Hz -0.0091183 -0.0199385
+ 1.042e+11Hz -0.00914441 -0.0199388
+ 1.043e+11Hz -0.00917052 -0.0199389
+ 1.044e+11Hz -0.00919662 -0.019939
+ 1.045e+11Hz -0.00922271 -0.0199391
+ 1.046e+11Hz -0.00924879 -0.0199391
+ 1.047e+11Hz -0.00927487 -0.0199391
+ 1.048e+11Hz -0.00930094 -0.019939
+ 1.049e+11Hz -0.009327 -0.0199389
+ 1.05e+11Hz -0.00935305 -0.0199388
+ 1.051e+11Hz -0.0093791 -0.0199385
+ 1.052e+11Hz -0.00940514 -0.0199383
+ 1.053e+11Hz -0.00943117 -0.019938
+ 1.054e+11Hz -0.00945719 -0.0199376
+ 1.055e+11Hz -0.00948321 -0.0199372
+ 1.056e+11Hz -0.00950921 -0.0199367
+ 1.057e+11Hz -0.00953521 -0.0199362
+ 1.058e+11Hz -0.0095612 -0.0199356
+ 1.059e+11Hz -0.00958718 -0.019935
+ 1.06e+11Hz -0.00961315 -0.0199343
+ 1.061e+11Hz -0.00963911 -0.0199336
+ 1.062e+11Hz -0.00966506 -0.0199328
+ 1.063e+11Hz -0.009691 -0.019932
+ 1.064e+11Hz -0.00971693 -0.0199311
+ 1.065e+11Hz -0.00974285 -0.0199302
+ 1.066e+11Hz -0.00976876 -0.0199292
+ 1.067e+11Hz -0.00979465 -0.0199281
+ 1.068e+11Hz -0.00982054 -0.019927
+ 1.069e+11Hz -0.00984641 -0.0199259
+ 1.07e+11Hz -0.00987228 -0.0199247
+ 1.071e+11Hz -0.00989813 -0.0199234
+ 1.072e+11Hz -0.00992397 -0.0199221
+ 1.073e+11Hz -0.00994979 -0.0199208
+ 1.074e+11Hz -0.0099756 -0.0199194
+ 1.075e+11Hz -0.0100014 -0.0199179
+ 1.076e+11Hz -0.0100272 -0.0199164
+ 1.077e+11Hz -0.010053 -0.0199148
+ 1.078e+11Hz -0.0100787 -0.0199132
+ 1.079e+11Hz -0.0101045 -0.0199115
+ 1.08e+11Hz -0.0101302 -0.0199097
+ 1.081e+11Hz -0.0101559 -0.0199079
+ 1.082e+11Hz -0.0101816 -0.0199061
+ 1.083e+11Hz -0.0102073 -0.0199042
+ 1.084e+11Hz -0.0102329 -0.0199022
+ 1.085e+11Hz -0.0102586 -0.0199002
+ 1.086e+11Hz -0.0102842 -0.0198981
+ 1.087e+11Hz -0.0103098 -0.019896
+ 1.088e+11Hz -0.0103354 -0.0198938
+ 1.089e+11Hz -0.010361 -0.0198916
+ 1.09e+11Hz -0.0103865 -0.0198893
+ 1.091e+11Hz -0.0104121 -0.0198869
+ 1.092e+11Hz -0.0104376 -0.0198845
+ 1.093e+11Hz -0.0104631 -0.0198821
+ 1.094e+11Hz -0.0104886 -0.0198796
+ 1.095e+11Hz -0.010514 -0.019877
+ 1.096e+11Hz -0.0105394 -0.0198744
+ 1.097e+11Hz -0.0105648 -0.0198717
+ 1.098e+11Hz -0.0105902 -0.0198689
+ 1.099e+11Hz -0.0106156 -0.0198661
+ 1.1e+11Hz -0.0106409 -0.0198633
+ 1.101e+11Hz -0.0106663 -0.0198604
+ 1.102e+11Hz -0.0106916 -0.0198574
+ 1.103e+11Hz -0.0107168 -0.0198544
+ 1.104e+11Hz -0.0107421 -0.0198513
+ 1.105e+11Hz -0.0107673 -0.0198482
+ 1.106e+11Hz -0.0107925 -0.019845
+ 1.107e+11Hz -0.0108177 -0.0198418
+ 1.108e+11Hz -0.0108428 -0.0198385
+ 1.109e+11Hz -0.0108679 -0.0198351
+ 1.11e+11Hz -0.010893 -0.0198317
+ 1.111e+11Hz -0.0109181 -0.0198283
+ 1.112e+11Hz -0.0109431 -0.0198248
+ 1.113e+11Hz -0.0109681 -0.0198212
+ 1.114e+11Hz -0.0109931 -0.0198176
+ 1.115e+11Hz -0.0110181 -0.0198139
+ 1.116e+11Hz -0.011043 -0.0198102
+ 1.117e+11Hz -0.0110679 -0.0198064
+ 1.118e+11Hz -0.0110927 -0.0198026
+ 1.119e+11Hz -0.0111176 -0.0197987
+ 1.12e+11Hz -0.0111424 -0.0197947
+ 1.121e+11Hz -0.0111671 -0.0197908
+ 1.122e+11Hz -0.0111919 -0.0197867
+ 1.123e+11Hz -0.0112166 -0.0197826
+ 1.124e+11Hz -0.0112412 -0.0197785
+ 1.125e+11Hz -0.0112659 -0.0197743
+ 1.126e+11Hz -0.0112905 -0.01977
+ 1.127e+11Hz -0.011315 -0.0197657
+ 1.128e+11Hz -0.0113396 -0.0197614
+ 1.129e+11Hz -0.0113641 -0.019757
+ 1.13e+11Hz -0.0113886 -0.0197525
+ 1.131e+11Hz -0.011413 -0.019748
+ 1.132e+11Hz -0.0114374 -0.0197435
+ 1.133e+11Hz -0.0114618 -0.0197389
+ 1.134e+11Hz -0.0114861 -0.0197342
+ 1.135e+11Hz -0.0115104 -0.0197295
+ 1.136e+11Hz -0.0115346 -0.0197248
+ 1.137e+11Hz -0.0115588 -0.01972
+ 1.138e+11Hz -0.011583 -0.0197151
+ 1.139e+11Hz -0.0116072 -0.0197102
+ 1.14e+11Hz -0.0116313 -0.0197053
+ 1.141e+11Hz -0.0116553 -0.0197003
+ 1.142e+11Hz -0.0116794 -0.0196953
+ 1.143e+11Hz -0.0117034 -0.0196902
+ 1.144e+11Hz -0.0117273 -0.0196851
+ 1.145e+11Hz -0.0117512 -0.0196799
+ 1.146e+11Hz -0.0117751 -0.0196747
+ 1.147e+11Hz -0.011799 -0.0196695
+ 1.148e+11Hz -0.0118228 -0.0196642
+ 1.149e+11Hz -0.0118465 -0.0196588
+ 1.15e+11Hz -0.0118702 -0.0196534
+ 1.151e+11Hz -0.0118939 -0.019648
+ 1.152e+11Hz -0.0119176 -0.0196425
+ 1.153e+11Hz -0.0119412 -0.019637
+ 1.154e+11Hz -0.0119647 -0.0196315
+ 1.155e+11Hz -0.0119883 -0.0196259
+ 1.156e+11Hz -0.0120117 -0.0196202
+ 1.157e+11Hz -0.0120352 -0.0196146
+ 1.158e+11Hz -0.0120586 -0.0196088
+ 1.159e+11Hz -0.0120819 -0.0196031
+ 1.16e+11Hz -0.0121053 -0.0195973
+ 1.161e+11Hz -0.0121285 -0.0195914
+ 1.162e+11Hz -0.0121518 -0.0195856
+ 1.163e+11Hz -0.012175 -0.0195797
+ 1.164e+11Hz -0.0121981 -0.0195737
+ 1.165e+11Hz -0.0122212 -0.0195677
+ 1.166e+11Hz -0.0122443 -0.0195617
+ 1.167e+11Hz -0.0122673 -0.0195556
+ 1.168e+11Hz -0.0122903 -0.0195495
+ 1.169e+11Hz -0.0123133 -0.0195434
+ 1.17e+11Hz -0.0123362 -0.0195372
+ 1.171e+11Hz -0.012359 -0.019531
+ 1.172e+11Hz -0.0123819 -0.0195248
+ 1.173e+11Hz -0.0124047 -0.0195185
+ 1.174e+11Hz -0.0124274 -0.0195122
+ 1.175e+11Hz -0.0124501 -0.0195059
+ 1.176e+11Hz -0.0124728 -0.0194995
+ 1.177e+11Hz -0.0124954 -0.0194931
+ 1.178e+11Hz -0.012518 -0.0194866
+ 1.179e+11Hz -0.0125405 -0.0194802
+ 1.18e+11Hz -0.012563 -0.0194737
+ 1.181e+11Hz -0.0125854 -0.0194671
+ 1.182e+11Hz -0.0126079 -0.0194606
+ 1.183e+11Hz -0.0126302 -0.019454
+ 1.184e+11Hz -0.0126526 -0.0194473
+ 1.185e+11Hz -0.0126749 -0.0194407
+ 1.186e+11Hz -0.0126971 -0.019434
+ 1.187e+11Hz -0.0127193 -0.0194273
+ 1.188e+11Hz -0.0127415 -0.0194205
+ 1.189e+11Hz -0.0127636 -0.0194137
+ 1.19e+11Hz -0.0127857 -0.0194069
+ 1.191e+11Hz -0.0128078 -0.0194001
+ 1.192e+11Hz -0.0128298 -0.0193932
+ 1.193e+11Hz -0.0128518 -0.0193863
+ 1.194e+11Hz -0.0128737 -0.0193794
+ 1.195e+11Hz -0.0128956 -0.0193725
+ 1.196e+11Hz -0.0129175 -0.0193655
+ 1.197e+11Hz -0.0129393 -0.0193585
+ 1.198e+11Hz -0.0129611 -0.0193515
+ 1.199e+11Hz -0.0129828 -0.0193444
+ 1.2e+11Hz -0.0130045 -0.0193373
+ 1.201e+11Hz -0.0130262 -0.0193302
+ 1.202e+11Hz -0.0130478 -0.0193231
+ 1.203e+11Hz -0.0130694 -0.0193159
+ 1.204e+11Hz -0.0130909 -0.0193088
+ 1.205e+11Hz -0.0131125 -0.0193016
+ 1.206e+11Hz -0.0131339 -0.0192943
+ 1.207e+11Hz -0.0131554 -0.0192871
+ 1.208e+11Hz -0.0131768 -0.0192798
+ 1.209e+11Hz -0.0131982 -0.0192725
+ 1.21e+11Hz -0.0132195 -0.0192651
+ 1.211e+11Hz -0.0132408 -0.0192578
+ 1.212e+11Hz -0.013262 -0.0192504
+ 1.213e+11Hz -0.0132833 -0.019243
+ 1.214e+11Hz -0.0133045 -0.0192356
+ 1.215e+11Hz -0.0133256 -0.0192281
+ 1.216e+11Hz -0.0133467 -0.0192206
+ 1.217e+11Hz -0.0133678 -0.0192131
+ 1.218e+11Hz -0.0133889 -0.0192056
+ 1.219e+11Hz -0.0134099 -0.0191981
+ 1.22e+11Hz -0.0134309 -0.0191905
+ 1.221e+11Hz -0.0134518 -0.0191829
+ 1.222e+11Hz -0.0134727 -0.0191753
+ 1.223e+11Hz -0.0134936 -0.0191676
+ 1.224e+11Hz -0.0135144 -0.01916
+ 1.225e+11Hz -0.0135353 -0.0191523
+ 1.226e+11Hz -0.013556 -0.0191446
+ 1.227e+11Hz -0.0135768 -0.0191369
+ 1.228e+11Hz -0.0135975 -0.0191291
+ 1.229e+11Hz -0.0136182 -0.0191213
+ 1.23e+11Hz -0.0136388 -0.0191135
+ 1.231e+11Hz -0.0136594 -0.0191057
+ 1.232e+11Hz -0.01368 -0.0190978
+ 1.233e+11Hz -0.0137006 -0.0190899
+ 1.234e+11Hz -0.0137211 -0.0190821
+ 1.235e+11Hz -0.0137416 -0.0190741
+ 1.236e+11Hz -0.013762 -0.0190662
+ 1.237e+11Hz -0.0137825 -0.0190582
+ 1.238e+11Hz -0.0138028 -0.0190502
+ 1.239e+11Hz -0.0138232 -0.0190422
+ 1.24e+11Hz -0.0138435 -0.0190342
+ 1.241e+11Hz -0.0138638 -0.0190261
+ 1.242e+11Hz -0.0138841 -0.019018
+ 1.243e+11Hz -0.0139043 -0.0190099
+ 1.244e+11Hz -0.0139246 -0.0190018
+ 1.245e+11Hz -0.0139447 -0.0189936
+ 1.246e+11Hz -0.0139649 -0.0189854
+ 1.247e+11Hz -0.013985 -0.0189772
+ 1.248e+11Hz -0.0140051 -0.018969
+ 1.249e+11Hz -0.0140251 -0.0189607
+ 1.25e+11Hz -0.0140452 -0.0189524
+ 1.251e+11Hz -0.0140652 -0.0189441
+ 1.252e+11Hz -0.0140851 -0.0189358
+ 1.253e+11Hz -0.0141051 -0.0189274
+ 1.254e+11Hz -0.014125 -0.018919
+ 1.255e+11Hz -0.0141448 -0.0189106
+ 1.256e+11Hz -0.0141647 -0.0189022
+ 1.257e+11Hz -0.0141845 -0.0188937
+ 1.258e+11Hz -0.0142043 -0.0188852
+ 1.259e+11Hz -0.0142241 -0.0188767
+ 1.26e+11Hz -0.0142438 -0.0188681
+ 1.261e+11Hz -0.0142635 -0.0188596
+ 1.262e+11Hz -0.0142831 -0.018851
+ 1.263e+11Hz -0.0143028 -0.0188423
+ 1.264e+11Hz -0.0143224 -0.0188337
+ 1.265e+11Hz -0.014342 -0.018825
+ 1.266e+11Hz -0.0143615 -0.0188163
+ 1.267e+11Hz -0.014381 -0.0188076
+ 1.268e+11Hz -0.0144005 -0.0187988
+ 1.269e+11Hz -0.01442 -0.01879
+ 1.27e+11Hz -0.0144394 -0.0187812
+ 1.271e+11Hz -0.0144588 -0.0187724
+ 1.272e+11Hz -0.0144781 -0.0187635
+ 1.273e+11Hz -0.0144975 -0.0187546
+ 1.274e+11Hz -0.0145168 -0.0187456
+ 1.275e+11Hz -0.014536 -0.0187367
+ 1.276e+11Hz -0.0145553 -0.0187277
+ 1.277e+11Hz -0.0145745 -0.0187187
+ 1.278e+11Hz -0.0145937 -0.0187096
+ 1.279e+11Hz -0.0146128 -0.0187005
+ 1.28e+11Hz -0.0146319 -0.0186914
+ 1.281e+11Hz -0.014651 -0.0186823
+ 1.282e+11Hz -0.01467 -0.0186731
+ 1.283e+11Hz -0.014689 -0.0186639
+ 1.284e+11Hz -0.014708 -0.0186547
+ 1.285e+11Hz -0.014727 -0.0186454
+ 1.286e+11Hz -0.0147459 -0.0186362
+ 1.287e+11Hz -0.0147648 -0.0186268
+ 1.288e+11Hz -0.0147836 -0.0186175
+ 1.289e+11Hz -0.0148024 -0.0186081
+ 1.29e+11Hz -0.0148212 -0.0185987
+ 1.291e+11Hz -0.0148399 -0.0185892
+ 1.292e+11Hz -0.0148587 -0.0185798
+ 1.293e+11Hz -0.0148773 -0.0185703
+ 1.294e+11Hz -0.014896 -0.0185607
+ 1.295e+11Hz -0.0149146 -0.0185512
+ 1.296e+11Hz -0.0149331 -0.0185416
+ 1.297e+11Hz -0.0149517 -0.0185319
+ 1.298e+11Hz -0.0149701 -0.0185223
+ 1.299e+11Hz -0.0149886 -0.0185126
+ 1.3e+11Hz -0.015007 -0.0185028
+ 1.301e+11Hz -0.0150254 -0.0184931
+ 1.302e+11Hz -0.0150437 -0.0184833
+ 1.303e+11Hz -0.015062 -0.0184735
+ 1.304e+11Hz -0.0150803 -0.0184636
+ 1.305e+11Hz -0.0150985 -0.0184537
+ 1.306e+11Hz -0.0151167 -0.0184438
+ 1.307e+11Hz -0.0151349 -0.0184339
+ 1.308e+11Hz -0.015153 -0.0184239
+ 1.309e+11Hz -0.015171 -0.0184139
+ 1.31e+11Hz -0.0151891 -0.0184039
+ 1.311e+11Hz -0.0152071 -0.0183938
+ 1.312e+11Hz -0.015225 -0.0183837
+ 1.313e+11Hz -0.0152429 -0.0183735
+ 1.314e+11Hz -0.0152608 -0.0183634
+ 1.315e+11Hz -0.0152786 -0.0183532
+ 1.316e+11Hz -0.0152963 -0.0183429
+ 1.317e+11Hz -0.0153141 -0.0183327
+ 1.318e+11Hz -0.0153318 -0.0183224
+ 1.319e+11Hz -0.0153494 -0.0183121
+ 1.32e+11Hz -0.015367 -0.0183017
+ 1.321e+11Hz -0.0153846 -0.0182913
+ 1.322e+11Hz -0.0154021 -0.0182809
+ 1.323e+11Hz -0.0154195 -0.0182705
+ 1.324e+11Hz -0.0154369 -0.01826
+ 1.325e+11Hz -0.0154543 -0.0182495
+ 1.326e+11Hz -0.0154716 -0.018239
+ 1.327e+11Hz -0.0154889 -0.0182284
+ 1.328e+11Hz -0.0155061 -0.0182178
+ 1.329e+11Hz -0.0155233 -0.0182072
+ 1.33e+11Hz -0.0155404 -0.0181966
+ 1.331e+11Hz -0.0155575 -0.0181859
+ 1.332e+11Hz -0.0155745 -0.0181752
+ 1.333e+11Hz -0.0155915 -0.0181645
+ 1.334e+11Hz -0.0156085 -0.0181537
+ 1.335e+11Hz -0.0156253 -0.0181429
+ 1.336e+11Hz -0.0156422 -0.0181321
+ 1.337e+11Hz -0.0156589 -0.0181212
+ 1.338e+11Hz -0.0156757 -0.0181104
+ 1.339e+11Hz -0.0156923 -0.0180995
+ 1.34e+11Hz -0.015709 -0.0180886
+ 1.341e+11Hz -0.0157255 -0.0180776
+ 1.342e+11Hz -0.0157421 -0.0180666
+ 1.343e+11Hz -0.0157585 -0.0180556
+ 1.344e+11Hz -0.0157749 -0.0180446
+ 1.345e+11Hz -0.0157913 -0.0180336
+ 1.346e+11Hz -0.0158076 -0.0180225
+ 1.347e+11Hz -0.0158238 -0.0180114
+ 1.348e+11Hz -0.01584 -0.0180003
+ 1.349e+11Hz -0.0158562 -0.0179892
+ 1.35e+11Hz -0.0158723 -0.017978
+ 1.351e+11Hz -0.0158883 -0.0179668
+ 1.352e+11Hz -0.0159043 -0.0179556
+ 1.353e+11Hz -0.0159202 -0.0179444
+ 1.354e+11Hz -0.015936 -0.0179332
+ 1.355e+11Hz -0.0159518 -0.0179219
+ 1.356e+11Hz -0.0159676 -0.0179106
+ 1.357e+11Hz -0.0159833 -0.0178993
+ 1.358e+11Hz -0.0159989 -0.017888
+ 1.359e+11Hz -0.0160145 -0.0178766
+ 1.36e+11Hz -0.01603 -0.0178653
+ 1.361e+11Hz -0.0160454 -0.0178539
+ 1.362e+11Hz -0.0160608 -0.0178425
+ 1.363e+11Hz -0.0160761 -0.0178311
+ 1.364e+11Hz -0.0160914 -0.0178197
+ 1.365e+11Hz -0.0161066 -0.0178082
+ 1.366e+11Hz -0.0161218 -0.0177968
+ 1.367e+11Hz -0.0161369 -0.0177853
+ 1.368e+11Hz -0.0161519 -0.0177738
+ 1.369e+11Hz -0.0161669 -0.0177623
+ 1.37e+11Hz -0.0161818 -0.0177508
+ 1.371e+11Hz -0.0161967 -0.0177393
+ 1.372e+11Hz -0.0162115 -0.0177278
+ 1.373e+11Hz -0.0162262 -0.0177162
+ 1.374e+11Hz -0.0162409 -0.0177047
+ 1.375e+11Hz -0.0162555 -0.0176931
+ 1.376e+11Hz -0.0162701 -0.0176816
+ 1.377e+11Hz -0.0162845 -0.01767
+ 1.378e+11Hz -0.016299 -0.0176584
+ 1.379e+11Hz -0.0163133 -0.0176468
+ 1.38e+11Hz -0.0163277 -0.0176352
+ 1.381e+11Hz -0.0163419 -0.0176236
+ 1.382e+11Hz -0.0163561 -0.0176119
+ 1.383e+11Hz -0.0163702 -0.0176003
+ 1.384e+11Hz -0.0163843 -0.0175887
+ 1.385e+11Hz -0.0163983 -0.0175771
+ 1.386e+11Hz -0.0164122 -0.0175654
+ 1.387e+11Hz -0.0164261 -0.0175538
+ 1.388e+11Hz -0.0164399 -0.0175421
+ 1.389e+11Hz -0.0164537 -0.0175305
+ 1.39e+11Hz -0.0164674 -0.0175188
+ 1.391e+11Hz -0.016481 -0.0175072
+ 1.392e+11Hz -0.0164946 -0.0174955
+ 1.393e+11Hz -0.0165081 -0.0174839
+ 1.394e+11Hz -0.0165215 -0.0174722
+ 1.395e+11Hz -0.0165349 -0.0174606
+ 1.396e+11Hz -0.0165482 -0.0174489
+ 1.397e+11Hz -0.0165615 -0.0174373
+ 1.398e+11Hz -0.0165747 -0.0174256
+ 1.399e+11Hz -0.0165879 -0.017414
+ 1.4e+11Hz -0.0166009 -0.0174024
+ 1.401e+11Hz -0.016614 -0.0173907
+ 1.402e+11Hz -0.0166269 -0.0173791
+ 1.403e+11Hz -0.0166398 -0.0173675
+ 1.404e+11Hz -0.0166527 -0.0173559
+ 1.405e+11Hz -0.0166655 -0.0173443
+ 1.406e+11Hz -0.0166782 -0.0173327
+ 1.407e+11Hz -0.0166908 -0.0173211
+ 1.408e+11Hz -0.0167035 -0.0173095
+ 1.409e+11Hz -0.016716 -0.0172979
+ 1.41e+11Hz -0.0167285 -0.0172863
+ 1.411e+11Hz -0.0167409 -0.0172748
+ 1.412e+11Hz -0.0167533 -0.0172632
+ 1.413e+11Hz -0.0167656 -0.0172517
+ 1.414e+11Hz -0.0167779 -0.0172402
+ 1.415e+11Hz -0.01679 -0.0172286
+ 1.416e+11Hz -0.0168022 -0.0172171
+ 1.417e+11Hz -0.0168143 -0.0172056
+ 1.418e+11Hz -0.0168263 -0.0171942
+ 1.419e+11Hz -0.0168383 -0.0171827
+ 1.42e+11Hz -0.0168502 -0.0171712
+ 1.421e+11Hz -0.016862 -0.0171598
+ 1.422e+11Hz -0.0168738 -0.0171484
+ 1.423e+11Hz -0.0168856 -0.017137
+ 1.424e+11Hz -0.0168973 -0.0171256
+ 1.425e+11Hz -0.0169089 -0.0171142
+ 1.426e+11Hz -0.0169205 -0.0171028
+ 1.427e+11Hz -0.016932 -0.0170915
+ 1.428e+11Hz -0.0169435 -0.0170801
+ 1.429e+11Hz -0.0169549 -0.0170688
+ 1.43e+11Hz -0.0169662 -0.0170575
+ 1.431e+11Hz -0.0169775 -0.0170463
+ 1.432e+11Hz -0.0169888 -0.017035
+ 1.433e+11Hz -0.017 -0.0170238
+ 1.434e+11Hz -0.0170112 -0.0170125
+ 1.435e+11Hz -0.0170223 -0.0170013
+ 1.436e+11Hz -0.0170333 -0.0169902
+ 1.437e+11Hz -0.0170443 -0.016979
+ 1.438e+11Hz -0.0170553 -0.0169679
+ 1.439e+11Hz -0.0170661 -0.0169567
+ 1.44e+11Hz -0.017077 -0.0169456
+ 1.441e+11Hz -0.0170878 -0.0169346
+ 1.442e+11Hz -0.0170985 -0.0169235
+ 1.443e+11Hz -0.0171092 -0.0169125
+ 1.444e+11Hz -0.0171199 -0.0169015
+ 1.445e+11Hz -0.0171305 -0.0168905
+ 1.446e+11Hz -0.017141 -0.0168795
+ 1.447e+11Hz -0.0171515 -0.0168686
+ 1.448e+11Hz -0.017162 -0.0168576
+ 1.449e+11Hz -0.0171724 -0.0168468
+ 1.45e+11Hz -0.0171828 -0.0168359
+ 1.451e+11Hz -0.0171931 -0.016825
+ 1.452e+11Hz -0.0172033 -0.0168142
+ 1.453e+11Hz -0.0172136 -0.0168034
+ 1.454e+11Hz -0.0172238 -0.0167926
+ 1.455e+11Hz -0.0172339 -0.0167819
+ 1.456e+11Hz -0.017244 -0.0167712
+ 1.457e+11Hz -0.017254 -0.0167605
+ 1.458e+11Hz -0.017264 -0.0167498
+ 1.459e+11Hz -0.017274 -0.0167391
+ 1.46e+11Hz -0.0172839 -0.0167285
+ 1.461e+11Hz -0.0172938 -0.0167179
+ 1.462e+11Hz -0.0173036 -0.0167073
+ 1.463e+11Hz -0.0173134 -0.0166968
+ 1.464e+11Hz -0.0173231 -0.0166863
+ 1.465e+11Hz -0.0173328 -0.0166758
+ 1.466e+11Hz -0.0173425 -0.0166653
+ 1.467e+11Hz -0.0173521 -0.0166549
+ 1.468e+11Hz -0.0173617 -0.0166445
+ 1.469e+11Hz -0.0173712 -0.0166341
+ 1.47e+11Hz -0.0173807 -0.0166237
+ 1.471e+11Hz -0.0173902 -0.0166134
+ 1.472e+11Hz -0.0173996 -0.0166031
+ 1.473e+11Hz -0.017409 -0.0165928
+ 1.474e+11Hz -0.0174183 -0.0165826
+ 1.475e+11Hz -0.0174276 -0.0165723
+ 1.476e+11Hz -0.0174369 -0.0165622
+ 1.477e+11Hz -0.0174461 -0.016552
+ 1.478e+11Hz -0.0174553 -0.0165419
+ 1.479e+11Hz -0.0174644 -0.0165317
+ 1.48e+11Hz -0.0174736 -0.0165217
+ 1.481e+11Hz -0.0174826 -0.0165116
+ 1.482e+11Hz -0.0174917 -0.0165016
+ 1.483e+11Hz -0.0175007 -0.0164916
+ 1.484e+11Hz -0.0175096 -0.0164816
+ 1.485e+11Hz -0.0175186 -0.0164717
+ 1.486e+11Hz -0.0175275 -0.0164618
+ 1.487e+11Hz -0.0175363 -0.0164519
+ 1.488e+11Hz -0.0175451 -0.0164421
+ 1.489e+11Hz -0.0175539 -0.0164322
+ 1.49e+11Hz -0.0175627 -0.0164224
+ 1.491e+11Hz -0.0175714 -0.0164127
+ 1.492e+11Hz -0.0175801 -0.016403
+ 1.493e+11Hz -0.0175887 -0.0163932
+ 1.494e+11Hz -0.0175973 -0.0163836
+ 1.495e+11Hz -0.0176059 -0.0163739
+ 1.496e+11Hz -0.0176144 -0.0163643
+ 1.497e+11Hz -0.0176229 -0.0163547
+ 1.498e+11Hz -0.0176314 -0.0163452
+ 1.499e+11Hz -0.0176399 -0.0163356
+ 1.5e+11Hz -0.0176483 -0.0163261
+ 1.501e+11Hz -0.0176566 -0.0163167
+ 1.502e+11Hz -0.017665 -0.0163072
+ 1.503e+11Hz -0.0176733 -0.0162978
+ 1.504e+11Hz -0.0176816 -0.0162885
+ 1.505e+11Hz -0.0176898 -0.0162791
+ 1.506e+11Hz -0.017698 -0.0162698
+ 1.507e+11Hz -0.0177062 -0.0162605
+ 1.508e+11Hz -0.0177144 -0.0162513
+ 1.509e+11Hz -0.0177225 -0.016242
+ 1.51e+11Hz -0.0177305 -0.0162329
+ 1.511e+11Hz -0.0177386 -0.0162237
+ 1.512e+11Hz -0.0177466 -0.0162146
+ 1.513e+11Hz -0.0177546 -0.0162055
+ 1.514e+11Hz -0.0177626 -0.0161964
+ 1.515e+11Hz -0.0177705 -0.0161874
+ 1.516e+11Hz -0.0177784 -0.0161784
+ 1.517e+11Hz -0.0177862 -0.0161694
+ 1.518e+11Hz -0.0177941 -0.0161605
+ 1.519e+11Hz -0.0178019 -0.0161516
+ 1.52e+11Hz -0.0178096 -0.0161427
+ 1.521e+11Hz -0.0178174 -0.0161338
+ 1.522e+11Hz -0.0178251 -0.016125
+ 1.523e+11Hz -0.0178327 -0.0161163
+ 1.524e+11Hz -0.0178404 -0.0161075
+ 1.525e+11Hz -0.017848 -0.0160988
+ 1.526e+11Hz -0.0178556 -0.0160901
+ 1.527e+11Hz -0.0178631 -0.0160815
+ 1.528e+11Hz -0.0178707 -0.0160729
+ 1.529e+11Hz -0.0178781 -0.0160643
+ 1.53e+11Hz -0.0178856 -0.0160558
+ 1.531e+11Hz -0.017893 -0.0160473
+ 1.532e+11Hz -0.0179004 -0.0160388
+ 1.533e+11Hz -0.0179078 -0.0160304
+ 1.534e+11Hz -0.0179152 -0.016022
+ 1.535e+11Hz -0.0179225 -0.0160137
+ 1.536e+11Hz -0.0179298 -0.0160053
+ 1.537e+11Hz -0.017937 -0.0159971
+ 1.538e+11Hz -0.0179442 -0.0159888
+ 1.539e+11Hz -0.0179514 -0.0159806
+ 1.54e+11Hz -0.0179586 -0.0159724
+ 1.541e+11Hz -0.0179657 -0.0159643
+ 1.542e+11Hz -0.0179728 -0.0159562
+ 1.543e+11Hz -0.0179799 -0.0159481
+ 1.544e+11Hz -0.017987 -0.0159401
+ 1.545e+11Hz -0.017994 -0.0159321
+ 1.546e+11Hz -0.018001 -0.0159242
+ 1.547e+11Hz -0.018008 -0.0159163
+ 1.548e+11Hz -0.0180149 -0.0159084
+ 1.549e+11Hz -0.0180218 -0.0159006
+ 1.55e+11Hz -0.0180287 -0.0158928
+ 1.551e+11Hz -0.0180355 -0.0158851
+ 1.552e+11Hz -0.0180424 -0.0158774
+ 1.553e+11Hz -0.0180492 -0.0158697
+ 1.554e+11Hz -0.0180559 -0.0158621
+ 1.555e+11Hz -0.0180627 -0.0158546
+ 1.556e+11Hz -0.0180694 -0.015847
+ 1.557e+11Hz -0.0180761 -0.0158396
+ 1.558e+11Hz -0.0180828 -0.0158321
+ 1.559e+11Hz -0.0180894 -0.0158247
+ 1.56e+11Hz -0.018096 -0.0158174
+ 1.561e+11Hz -0.0181026 -0.0158101
+ 1.562e+11Hz -0.0181092 -0.0158028
+ 1.563e+11Hz -0.0181157 -0.0157956
+ 1.564e+11Hz -0.0181222 -0.0157885
+ 1.565e+11Hz -0.0181287 -0.0157814
+ 1.566e+11Hz -0.0181352 -0.0157743
+ 1.567e+11Hz -0.0181416 -0.0157673
+ 1.568e+11Hz -0.018148 -0.0157603
+ 1.569e+11Hz -0.0181544 -0.0157534
+ 1.57e+11Hz -0.0181608 -0.0157465
+ 1.571e+11Hz -0.0181672 -0.0157397
+ 1.572e+11Hz -0.0181735 -0.0157329
+ 1.573e+11Hz -0.0181798 -0.0157262
+ 1.574e+11Hz -0.0181861 -0.0157196
+ 1.575e+11Hz -0.0181924 -0.0157129
+ 1.576e+11Hz -0.0181986 -0.0157064
+ 1.577e+11Hz -0.0182048 -0.0156999
+ 1.578e+11Hz -0.018211 -0.0156934
+ 1.579e+11Hz -0.0182172 -0.015687
+ 1.58e+11Hz -0.0182234 -0.0156807
+ 1.581e+11Hz -0.0182295 -0.0156744
+ 1.582e+11Hz -0.0182357 -0.0156682
+ 1.583e+11Hz -0.0182418 -0.015662
+ 1.584e+11Hz -0.0182479 -0.0156559
+ 1.585e+11Hz -0.018254 -0.0156498
+ 1.586e+11Hz -0.01826 -0.0156438
+ 1.587e+11Hz -0.0182661 -0.0156379
+ 1.588e+11Hz -0.0182721 -0.015632
+ 1.589e+11Hz -0.0182781 -0.0156262
+ 1.59e+11Hz -0.0182842 -0.0156204
+ 1.591e+11Hz -0.0182901 -0.0156147
+ 1.592e+11Hz -0.0182961 -0.0156091
+ 1.593e+11Hz -0.0183021 -0.0156035
+ 1.594e+11Hz -0.0183081 -0.015598
+ 1.595e+11Hz -0.018314 -0.0155925
+ 1.596e+11Hz -0.01832 -0.0155871
+ 1.597e+11Hz -0.0183259 -0.0155818
+ 1.598e+11Hz -0.0183318 -0.0155765
+ 1.599e+11Hz -0.0183378 -0.0155713
+ 1.6e+11Hz -0.0183437 -0.0155662
+ 1.601e+11Hz -0.0183496 -0.0155611
+ 1.602e+11Hz -0.0183555 -0.0155561
+ 1.603e+11Hz -0.0183614 -0.0155512
+ 1.604e+11Hz -0.0183673 -0.0155463
+ 1.605e+11Hz -0.0183732 -0.0155415
+ 1.606e+11Hz -0.0183791 -0.0155368
+ 1.607e+11Hz -0.018385 -0.0155321
+ 1.608e+11Hz -0.0183909 -0.0155275
+ 1.609e+11Hz -0.0183967 -0.0155229
+ 1.61e+11Hz -0.0184026 -0.0155185
+ 1.611e+11Hz -0.0184085 -0.0155141
+ 1.612e+11Hz -0.0184144 -0.0155098
+ 1.613e+11Hz -0.0184204 -0.0155055
+ 1.614e+11Hz -0.0184263 -0.0155013
+ 1.615e+11Hz -0.0184322 -0.0154972
+ 1.616e+11Hz -0.0184381 -0.0154932
+ 1.617e+11Hz -0.0184441 -0.0154892
+ 1.618e+11Hz -0.01845 -0.0154853
+ 1.619e+11Hz -0.018456 -0.0154814
+ 1.62e+11Hz -0.0184619 -0.0154777
+ 1.621e+11Hz -0.0184679 -0.015474
+ 1.622e+11Hz -0.0184739 -0.0154704
+ 1.623e+11Hz -0.0184799 -0.0154668
+ 1.624e+11Hz -0.0184859 -0.0154634
+ 1.625e+11Hz -0.018492 -0.01546
+ 1.626e+11Hz -0.018498 -0.0154567
+ 1.627e+11Hz -0.0185041 -0.0154534
+ 1.628e+11Hz -0.0185102 -0.0154502
+ 1.629e+11Hz -0.0185164 -0.0154471
+ 1.63e+11Hz -0.0185225 -0.0154441
+ 1.631e+11Hz -0.0185287 -0.0154411
+ 1.632e+11Hz -0.0185349 -0.0154383
+ 1.633e+11Hz -0.0185411 -0.0154354
+ 1.634e+11Hz -0.0185473 -0.0154327
+ 1.635e+11Hz -0.0185536 -0.01543
+ 1.636e+11Hz -0.0185599 -0.0154275
+ 1.637e+11Hz -0.0185663 -0.0154249
+ 1.638e+11Hz -0.0185726 -0.0154225
+ 1.639e+11Hz -0.018579 -0.0154201
+ 1.64e+11Hz -0.0185855 -0.0154178
+ 1.641e+11Hz -0.018592 -0.0154156
+ 1.642e+11Hz -0.0185985 -0.0154135
+ 1.643e+11Hz -0.018605 -0.0154114
+ 1.644e+11Hz -0.0186116 -0.0154094
+ 1.645e+11Hz -0.0186183 -0.0154075
+ 1.646e+11Hz -0.0186249 -0.0154056
+ 1.647e+11Hz -0.0186316 -0.0154038
+ 1.648e+11Hz -0.0186384 -0.0154021
+ 1.649e+11Hz -0.0186452 -0.0154005
+ 1.65e+11Hz -0.0186521 -0.0153989
+ 1.651e+11Hz -0.018659 -0.0153974
+ 1.652e+11Hz -0.0186659 -0.0153959
+ 1.653e+11Hz -0.0186729 -0.0153946
+ 1.654e+11Hz -0.01868 -0.0153933
+ 1.655e+11Hz -0.0186871 -0.0153921
+ 1.656e+11Hz -0.0186943 -0.0153909
+ 1.657e+11Hz -0.0187015 -0.0153898
+ 1.658e+11Hz -0.0187088 -0.0153888
+ 1.659e+11Hz -0.0187161 -0.0153878
+ 1.66e+11Hz -0.0187235 -0.015387
+ 1.661e+11Hz -0.018731 -0.0153861
+ 1.662e+11Hz -0.0187385 -0.0153854
+ 1.663e+11Hz -0.0187461 -0.0153847
+ 1.664e+11Hz -0.0187538 -0.0153841
+ 1.665e+11Hz -0.0187615 -0.0153835
+ 1.666e+11Hz -0.0187693 -0.015383
+ 1.667e+11Hz -0.0187771 -0.0153826
+ 1.668e+11Hz -0.0187851 -0.0153822
+ 1.669e+11Hz -0.0187931 -0.0153819
+ 1.67e+11Hz -0.0188011 -0.0153816
+ 1.671e+11Hz -0.0188093 -0.0153814
+ 1.672e+11Hz -0.0188175 -0.0153813
+ 1.673e+11Hz -0.0188258 -0.0153812
+ 1.674e+11Hz -0.0188342 -0.0153812
+ 1.675e+11Hz -0.0188426 -0.0153812
+ 1.676e+11Hz -0.0188512 -0.0153813
+ 1.677e+11Hz -0.0188598 -0.0153814
+ 1.678e+11Hz -0.0188685 -0.0153816
+ 1.679e+11Hz -0.0188773 -0.0153818
+ 1.68e+11Hz -0.0188861 -0.0153821
+ 1.681e+11Hz -0.0188951 -0.0153825
+ 1.682e+11Hz -0.0189041 -0.0153828
+ 1.683e+11Hz -0.0189132 -0.0153833
+ 1.684e+11Hz -0.0189225 -0.0153837
+ 1.685e+11Hz -0.0189318 -0.0153843
+ 1.686e+11Hz -0.0189412 -0.0153848
+ 1.687e+11Hz -0.0189506 -0.0153854
+ 1.688e+11Hz -0.0189602 -0.0153861
+ 1.689e+11Hz -0.0189699 -0.0153868
+ 1.69e+11Hz -0.0189797 -0.0153875
+ 1.691e+11Hz -0.0189895 -0.0153883
+ 1.692e+11Hz -0.0189995 -0.0153891
+ 1.693e+11Hz -0.0190095 -0.0153899
+ 1.694e+11Hz -0.0190197 -0.0153908
+ 1.695e+11Hz -0.01903 -0.0153917
+ 1.696e+11Hz -0.0190403 -0.0153926
+ 1.697e+11Hz -0.0190508 -0.0153936
+ 1.698e+11Hz -0.0190613 -0.0153946
+ 1.699e+11Hz -0.019072 -0.0153956
+ 1.7e+11Hz -0.0190828 -0.0153966
+ 1.701e+11Hz -0.0190936 -0.0153977
+ 1.702e+11Hz -0.0191046 -0.0153988
+ 1.703e+11Hz -0.0191157 -0.0153999
+ 1.704e+11Hz -0.0191269 -0.015401
+ 1.705e+11Hz -0.0191382 -0.0154022
+ 1.706e+11Hz -0.0191496 -0.0154034
+ 1.707e+11Hz -0.0191611 -0.0154045
+ 1.708e+11Hz -0.0191727 -0.0154057
+ 1.709e+11Hz -0.0191844 -0.0154069
+ 1.71e+11Hz -0.0191963 -0.0154081
+ 1.711e+11Hz -0.0192082 -0.0154094
+ 1.712e+11Hz -0.0192203 -0.0154106
+ 1.713e+11Hz -0.0192325 -0.0154118
+ 1.714e+11Hz -0.0192447 -0.0154131
+ 1.715e+11Hz -0.0192571 -0.0154143
+ 1.716e+11Hz -0.0192696 -0.0154155
+ 1.717e+11Hz -0.0192823 -0.0154168
+ 1.718e+11Hz -0.019295 -0.015418
+ 1.719e+11Hz -0.0193079 -0.0154192
+ 1.72e+11Hz -0.0193208 -0.0154205
+ 1.721e+11Hz -0.0193339 -0.0154217
+ 1.722e+11Hz -0.0193471 -0.0154229
+ 1.723e+11Hz -0.0193604 -0.0154241
+ 1.724e+11Hz -0.0193738 -0.0154252
+ 1.725e+11Hz -0.0193874 -0.0154264
+ 1.726e+11Hz -0.019401 -0.0154276
+ 1.727e+11Hz -0.0194148 -0.0154287
+ 1.728e+11Hz -0.0194287 -0.0154298
+ 1.729e+11Hz -0.0194427 -0.0154309
+ 1.73e+11Hz -0.0194568 -0.0154319
+ 1.731e+11Hz -0.019471 -0.015433
+ 1.732e+11Hz -0.0194854 -0.015434
+ 1.733e+11Hz -0.0194999 -0.015435
+ 1.734e+11Hz -0.0195144 -0.0154359
+ 1.735e+11Hz -0.0195291 -0.0154368
+ 1.736e+11Hz -0.0195439 -0.0154377
+ 1.737e+11Hz -0.0195589 -0.0154386
+ 1.738e+11Hz -0.0195739 -0.0154394
+ 1.739e+11Hz -0.019589 -0.0154402
+ 1.74e+11Hz -0.0196043 -0.0154409
+ 1.741e+11Hz -0.0196197 -0.0154416
+ 1.742e+11Hz -0.0196352 -0.0154422
+ 1.743e+11Hz -0.0196508 -0.0154428
+ 1.744e+11Hz -0.0196665 -0.0154434
+ 1.745e+11Hz -0.0196823 -0.0154439
+ 1.746e+11Hz -0.0196983 -0.0154443
+ 1.747e+11Hz -0.0197143 -0.0154447
+ 1.748e+11Hz -0.0197305 -0.015445
+ 1.749e+11Hz -0.0197468 -0.0154453
+ 1.75e+11Hz -0.0197632 -0.0154455
+ 1.751e+11Hz -0.0197797 -0.0154457
+ 1.752e+11Hz -0.0197963 -0.0154458
+ 1.753e+11Hz -0.019813 -0.0154459
+ 1.754e+11Hz -0.0198298 -0.0154458
+ 1.755e+11Hz -0.0198467 -0.0154457
+ 1.756e+11Hz -0.0198637 -0.0154456
+ 1.757e+11Hz -0.0198809 -0.0154453
+ 1.758e+11Hz -0.0198981 -0.015445
+ 1.759e+11Hz -0.0199154 -0.0154447
+ 1.76e+11Hz -0.0199329 -0.0154442
+ 1.761e+11Hz -0.0199504 -0.0154437
+ 1.762e+11Hz -0.0199681 -0.0154431
+ 1.763e+11Hz -0.0199858 -0.0154424
+ 1.764e+11Hz -0.0200037 -0.0154416
+ 1.765e+11Hz -0.0200216 -0.0154408
+ 1.766e+11Hz -0.0200397 -0.0154399
+ 1.767e+11Hz -0.0200578 -0.0154389
+ 1.768e+11Hz -0.020076 -0.0154378
+ 1.769e+11Hz -0.0200943 -0.0154366
+ 1.77e+11Hz -0.0201128 -0.0154353
+ 1.771e+11Hz -0.0201313 -0.0154339
+ 1.772e+11Hz -0.0201499 -0.0154325
+ 1.773e+11Hz -0.0201685 -0.0154309
+ 1.774e+11Hz -0.0201873 -0.0154293
+ 1.775e+11Hz -0.0202062 -0.0154275
+ 1.776e+11Hz -0.0202251 -0.0154257
+ 1.777e+11Hz -0.0202442 -0.0154237
+ 1.778e+11Hz -0.0202633 -0.0154217
+ 1.779e+11Hz -0.0202825 -0.0154196
+ 1.78e+11Hz -0.0203018 -0.0154173
+ 1.781e+11Hz -0.0203211 -0.015415
+ 1.782e+11Hz -0.0203406 -0.0154125
+ 1.783e+11Hz -0.0203601 -0.01541
+ 1.784e+11Hz -0.0203797 -0.0154073
+ 1.785e+11Hz -0.0203993 -0.0154045
+ 1.786e+11Hz -0.0204191 -0.0154016
+ 1.787e+11Hz -0.0204389 -0.0153986
+ 1.788e+11Hz -0.0204588 -0.0153955
+ 1.789e+11Hz -0.0204787 -0.0153923
+ 1.79e+11Hz -0.0204987 -0.015389
+ 1.791e+11Hz -0.0205188 -0.0153855
+ 1.792e+11Hz -0.0205389 -0.015382
+ 1.793e+11Hz -0.0205592 -0.0153783
+ 1.794e+11Hz -0.0205794 -0.0153745
+ 1.795e+11Hz -0.0205997 -0.0153706
+ 1.796e+11Hz -0.0206201 -0.0153666
+ 1.797e+11Hz -0.0206406 -0.0153624
+ 1.798e+11Hz -0.0206611 -0.0153581
+ 1.799e+11Hz -0.0206816 -0.0153538
+ 1.8e+11Hz -0.0207022 -0.0153492
+ 1.801e+11Hz -0.0207229 -0.0153446
+ 1.802e+11Hz -0.0207436 -0.0153399
+ 1.803e+11Hz -0.0207643 -0.015335
+ 1.804e+11Hz -0.0207851 -0.01533
+ 1.805e+11Hz -0.020806 -0.0153248
+ 1.806e+11Hz -0.0208269 -0.0153196
+ 1.807e+11Hz -0.0208478 -0.0153142
+ 1.808e+11Hz -0.0208688 -0.0153087
+ 1.809e+11Hz -0.0208898 -0.015303
+ 1.81e+11Hz -0.0209108 -0.0152973
+ 1.811e+11Hz -0.0209319 -0.0152914
+ 1.812e+11Hz -0.020953 -0.0152854
+ 1.813e+11Hz -0.0209741 -0.0152792
+ 1.814e+11Hz -0.0209953 -0.0152729
+ 1.815e+11Hz -0.0210165 -0.0152665
+ 1.816e+11Hz -0.0210377 -0.01526
+ 1.817e+11Hz -0.0210589 -0.0152533
+ 1.818e+11Hz -0.0210802 -0.0152465
+ 1.819e+11Hz -0.0211015 -0.0152396
+ 1.82e+11Hz -0.0211228 -0.0152325
+ 1.821e+11Hz -0.0211441 -0.0152253
+ 1.822e+11Hz -0.0211655 -0.015218
+ 1.823e+11Hz -0.0211868 -0.0152105
+ 1.824e+11Hz -0.0212082 -0.0152029
+ 1.825e+11Hz -0.0212296 -0.0151952
+ 1.826e+11Hz -0.021251 -0.0151874
+ 1.827e+11Hz -0.0212724 -0.0151794
+ 1.828e+11Hz -0.0212938 -0.0151713
+ 1.829e+11Hz -0.0213152 -0.015163
+ 1.83e+11Hz -0.0213367 -0.0151546
+ 1.831e+11Hz -0.0213581 -0.0151461
+ 1.832e+11Hz -0.0213795 -0.0151375
+ 1.833e+11Hz -0.0214009 -0.0151287
+ 1.834e+11Hz -0.0214223 -0.0151198
+ 1.835e+11Hz -0.0214438 -0.0151107
+ 1.836e+11Hz -0.0214652 -0.0151016
+ 1.837e+11Hz -0.0214866 -0.0150923
+ 1.838e+11Hz -0.021508 -0.0150828
+ 1.839e+11Hz -0.0215293 -0.0150733
+ 1.84e+11Hz -0.0215507 -0.0150636
+ 1.841e+11Hz -0.0215721 -0.0150538
+ 1.842e+11Hz -0.0215934 -0.0150438
+ 1.843e+11Hz -0.0216147 -0.0150337
+ 1.844e+11Hz -0.021636 -0.0150235
+ 1.845e+11Hz -0.0216573 -0.0150132
+ 1.846e+11Hz -0.0216786 -0.0150027
+ 1.847e+11Hz -0.0216998 -0.0149921
+ 1.848e+11Hz -0.021721 -0.0149814
+ 1.849e+11Hz -0.0217422 -0.0149705
+ 1.85e+11Hz -0.0217634 -0.0149595
+ 1.851e+11Hz -0.0217845 -0.0149484
+ 1.852e+11Hz -0.0218057 -0.0149372
+ 1.853e+11Hz -0.0218267 -0.0149258
+ 1.854e+11Hz -0.0218478 -0.0149144
+ 1.855e+11Hz -0.0218688 -0.0149028
+ 1.856e+11Hz -0.0218898 -0.014891
+ 1.857e+11Hz -0.0219107 -0.0148792
+ 1.858e+11Hz -0.0219316 -0.0148672
+ 1.859e+11Hz -0.0219525 -0.0148551
+ 1.86e+11Hz -0.0219733 -0.0148429
+ 1.861e+11Hz -0.0219941 -0.0148306
+ 1.862e+11Hz -0.0220148 -0.0148181
+ 1.863e+11Hz -0.0220355 -0.0148055
+ 1.864e+11Hz -0.0220561 -0.0147928
+ 1.865e+11Hz -0.0220767 -0.01478
+ 1.866e+11Hz -0.0220973 -0.0147671
+ 1.867e+11Hz -0.0221178 -0.014754
+ 1.868e+11Hz -0.0221382 -0.0147409
+ 1.869e+11Hz -0.0221586 -0.0147276
+ 1.87e+11Hz -0.022179 -0.0147142
+ 1.871e+11Hz -0.0221993 -0.0147007
+ 1.872e+11Hz -0.0222195 -0.0146871
+ 1.873e+11Hz -0.0222397 -0.0146734
+ 1.874e+11Hz -0.0222598 -0.0146595
+ 1.875e+11Hz -0.0222799 -0.0146456
+ 1.876e+11Hz -0.0222999 -0.0146315
+ 1.877e+11Hz -0.0223198 -0.0146174
+ 1.878e+11Hz -0.0223397 -0.0146031
+ 1.879e+11Hz -0.0223595 -0.0145887
+ 1.88e+11Hz -0.0223793 -0.0145742
+ 1.881e+11Hz -0.022399 -0.0145597
+ 1.882e+11Hz -0.0224186 -0.014545
+ 1.883e+11Hz -0.0224381 -0.0145302
+ 1.884e+11Hz -0.0224576 -0.0145153
+ 1.885e+11Hz -0.022477 -0.0145003
+ 1.886e+11Hz -0.0224964 -0.0144852
+ 1.887e+11Hz -0.0225157 -0.01447
+ 1.888e+11Hz -0.0225349 -0.0144547
+ 1.889e+11Hz -0.022554 -0.0144393
+ 1.89e+11Hz -0.0225731 -0.0144238
+ 1.891e+11Hz -0.0225921 -0.0144082
+ 1.892e+11Hz -0.022611 -0.0143926
+ 1.893e+11Hz -0.0226298 -0.0143768
+ 1.894e+11Hz -0.0226486 -0.0143609
+ 1.895e+11Hz -0.0226673 -0.014345
+ 1.896e+11Hz -0.0226859 -0.0143289
+ 1.897e+11Hz -0.0227044 -0.0143128
+ 1.898e+11Hz -0.0227228 -0.0142966
+ 1.899e+11Hz -0.0227412 -0.0142803
+ 1.9e+11Hz -0.0227595 -0.0142639
+ 1.901e+11Hz -0.0227777 -0.0142474
+ 1.902e+11Hz -0.0227958 -0.0142308
+ 1.903e+11Hz -0.0228138 -0.0142142
+ 1.904e+11Hz -0.0228318 -0.0141975
+ 1.905e+11Hz -0.0228496 -0.0141807
+ 1.906e+11Hz -0.0228674 -0.0141638
+ 1.907e+11Hz -0.0228851 -0.0141468
+ 1.908e+11Hz -0.0229027 -0.0141298
+ 1.909e+11Hz -0.0229203 -0.0141127
+ 1.91e+11Hz -0.0229377 -0.0140955
+ 1.911e+11Hz -0.022955 -0.0140782
+ 1.912e+11Hz -0.0229723 -0.0140609
+ 1.913e+11Hz -0.0229894 -0.0140434
+ 1.914e+11Hz -0.0230065 -0.014026
+ 1.915e+11Hz -0.0230235 -0.0140084
+ 1.916e+11Hz -0.0230404 -0.0139908
+ 1.917e+11Hz -0.0230572 -0.0139731
+ 1.918e+11Hz -0.0230739 -0.0139553
+ 1.919e+11Hz -0.0230905 -0.0139375
+ 1.92e+11Hz -0.0231071 -0.0139196
+ 1.921e+11Hz -0.0231235 -0.0139017
+ 1.922e+11Hz -0.0231398 -0.0138837
+ 1.923e+11Hz -0.0231561 -0.0138656
+ 1.924e+11Hz -0.0231722 -0.0138475
+ 1.925e+11Hz -0.0231883 -0.0138293
+ 1.926e+11Hz -0.0232042 -0.013811
+ 1.927e+11Hz -0.0232201 -0.0137927
+ 1.928e+11Hz -0.0232359 -0.0137744
+ 1.929e+11Hz -0.0232516 -0.013756
+ 1.93e+11Hz -0.0232671 -0.0137375
+ 1.931e+11Hz -0.0232826 -0.013719
+ 1.932e+11Hz -0.023298 -0.0137004
+ 1.933e+11Hz -0.0233133 -0.0136818
+ 1.934e+11Hz -0.0233285 -0.0136631
+ 1.935e+11Hz -0.0233435 -0.0136444
+ 1.936e+11Hz -0.0233585 -0.0136257
+ 1.937e+11Hz -0.0233734 -0.0136069
+ 1.938e+11Hz -0.0233882 -0.013588
+ 1.939e+11Hz -0.0234029 -0.0135691
+ 1.94e+11Hz -0.0234175 -0.0135502
+ 1.941e+11Hz -0.023432 -0.0135312
+ 1.942e+11Hz -0.0234464 -0.0135122
+ 1.943e+11Hz -0.0234607 -0.0134932
+ 1.944e+11Hz -0.0234749 -0.0134741
+ 1.945e+11Hz -0.023489 -0.013455
+ 1.946e+11Hz -0.023503 -0.0134358
+ 1.947e+11Hz -0.0235169 -0.0134167
+ 1.948e+11Hz -0.0235307 -0.0133974
+ 1.949e+11Hz -0.0235444 -0.0133782
+ 1.95e+11Hz -0.023558 -0.0133589
+ 1.951e+11Hz -0.0235714 -0.0133396
+ 1.952e+11Hz -0.0235848 -0.0133203
+ 1.953e+11Hz -0.0235981 -0.0133009
+ 1.954e+11Hz -0.0236113 -0.0132815
+ 1.955e+11Hz -0.0236244 -0.0132621
+ 1.956e+11Hz -0.0236374 -0.0132427
+ 1.957e+11Hz -0.0236503 -0.0132232
+ 1.958e+11Hz -0.0236631 -0.0132038
+ 1.959e+11Hz -0.0236758 -0.0131843
+ 1.96e+11Hz -0.0236884 -0.0131648
+ 1.961e+11Hz -0.0237009 -0.0131453
+ 1.962e+11Hz -0.0237132 -0.0131257
+ 1.963e+11Hz -0.0237255 -0.0131062
+ 1.964e+11Hz -0.0237377 -0.0130866
+ 1.965e+11Hz -0.0237498 -0.013067
+ 1.966e+11Hz -0.0237618 -0.0130474
+ 1.967e+11Hz -0.0237737 -0.0130278
+ 1.968e+11Hz -0.0237855 -0.0130082
+ 1.969e+11Hz -0.0237972 -0.0129886
+ 1.97e+11Hz -0.0238088 -0.012969
+ 1.971e+11Hz -0.0238202 -0.0129494
+ 1.972e+11Hz -0.0238316 -0.0129297
+ 1.973e+11Hz -0.0238429 -0.0129101
+ 1.974e+11Hz -0.0238541 -0.0128905
+ 1.975e+11Hz -0.0238652 -0.0128709
+ 1.976e+11Hz -0.0238762 -0.0128512
+ 1.977e+11Hz -0.0238871 -0.0128316
+ 1.978e+11Hz -0.0238979 -0.012812
+ 1.979e+11Hz -0.0239087 -0.0127924
+ 1.98e+11Hz -0.0239193 -0.0127728
+ 1.981e+11Hz -0.0239298 -0.0127532
+ 1.982e+11Hz -0.0239402 -0.0127336
+ 1.983e+11Hz -0.0239505 -0.012714
+ 1.984e+11Hz -0.0239608 -0.0126944
+ 1.985e+11Hz -0.0239709 -0.0126749
+ 1.986e+11Hz -0.023981 -0.0126553
+ 1.987e+11Hz -0.0239909 -0.0126358
+ 1.988e+11Hz -0.0240008 -0.0126163
+ 1.989e+11Hz -0.0240105 -0.0125968
+ 1.99e+11Hz -0.0240202 -0.0125773
+ 1.991e+11Hz -0.0240298 -0.0125579
+ 1.992e+11Hz -0.0240393 -0.0125385
+ 1.993e+11Hz -0.0240487 -0.012519
+ 1.994e+11Hz -0.024058 -0.0124997
+ 1.995e+11Hz -0.0240672 -0.0124803
+ 1.996e+11Hz -0.0240764 -0.0124609
+ 1.997e+11Hz -0.0240854 -0.0124416
+ 1.998e+11Hz -0.0240944 -0.0124224
+ 1.999e+11Hz -0.0241033 -0.0124031
+ 2e+11Hz -0.0241121 -0.0123839
+ 2.001e+11Hz -0.0241208 -0.0123647
+ 2.002e+11Hz -0.0241294 -0.0123455
+ 2.003e+11Hz -0.0241379 -0.0123264
+ 2.004e+11Hz -0.0241464 -0.0123073
+ 2.005e+11Hz -0.0241548 -0.0122883
+ 2.006e+11Hz -0.0241631 -0.0122693
+ 2.007e+11Hz -0.0241713 -0.0122503
+ 2.008e+11Hz -0.0241794 -0.0122313
+ 2.009e+11Hz -0.0241875 -0.0122124
+ 2.01e+11Hz -0.0241955 -0.0121936
+ 2.011e+11Hz -0.0242034 -0.0121748
+ 2.012e+11Hz -0.0242112 -0.012156
+ 2.013e+11Hz -0.024219 -0.0121373
+ 2.014e+11Hz -0.0242267 -0.0121186
+ 2.015e+11Hz -0.0242343 -0.0121
+ 2.016e+11Hz -0.0242418 -0.0120814
+ 2.017e+11Hz -0.0242493 -0.0120629
+ 2.018e+11Hz -0.0242567 -0.0120444
+ 2.019e+11Hz -0.024264 -0.012026
+ 2.02e+11Hz -0.0242713 -0.0120076
+ 2.021e+11Hz -0.0242785 -0.0119893
+ 2.022e+11Hz -0.0242856 -0.011971
+ 2.023e+11Hz -0.0242927 -0.0119528
+ 2.024e+11Hz -0.0242997 -0.0119347
+ 2.025e+11Hz -0.0243067 -0.0119166
+ 2.026e+11Hz -0.0243136 -0.0118985
+ 2.027e+11Hz -0.0243204 -0.0118805
+ 2.028e+11Hz -0.0243272 -0.0118626
+ 2.029e+11Hz -0.0243339 -0.0118448
+ 2.03e+11Hz -0.0243406 -0.011827
+ 2.031e+11Hz -0.0243472 -0.0118093
+ 2.032e+11Hz -0.0243538 -0.0117916
+ 2.033e+11Hz -0.0243603 -0.011774
+ 2.034e+11Hz -0.0243668 -0.0117564
+ 2.035e+11Hz -0.0243732 -0.011739
+ 2.036e+11Hz -0.0243796 -0.0117216
+ 2.037e+11Hz -0.0243859 -0.0117042
+ 2.038e+11Hz -0.0243922 -0.011687
+ 2.039e+11Hz -0.0243984 -0.0116698
+ 2.04e+11Hz -0.0244046 -0.0116526
+ 2.041e+11Hz -0.0244108 -0.0116356
+ 2.042e+11Hz -0.024417 -0.0116186
+ 2.043e+11Hz -0.0244231 -0.0116017
+ 2.044e+11Hz -0.0244291 -0.0115848
+ 2.045e+11Hz -0.0244352 -0.0115681
+ 2.046e+11Hz -0.0244412 -0.0115514
+ 2.047e+11Hz -0.0244472 -0.0115348
+ 2.048e+11Hz -0.0244531 -0.0115182
+ 2.049e+11Hz -0.0244591 -0.0115017
+ 2.05e+11Hz -0.024465 -0.0114853
+ 2.051e+11Hz -0.0244709 -0.011469
+ 2.052e+11Hz -0.0244767 -0.0114528
+ 2.053e+11Hz -0.0244826 -0.0114366
+ 2.054e+11Hz -0.0244884 -0.0114205
+ 2.055e+11Hz -0.0244943 -0.0114045
+ 2.056e+11Hz -0.0245001 -0.0113886
+ 2.057e+11Hz -0.0245059 -0.0113727
+ 2.058e+11Hz -0.0245117 -0.0113569
+ 2.059e+11Hz -0.0245175 -0.0113412
+ 2.06e+11Hz -0.0245233 -0.0113256
+ 2.061e+11Hz -0.0245291 -0.0113101
+ 2.062e+11Hz -0.0245349 -0.0112946
+ 2.063e+11Hz -0.0245407 -0.0112792
+ 2.064e+11Hz -0.0245465 -0.0112639
+ 2.065e+11Hz -0.0245523 -0.0112487
+ 2.066e+11Hz -0.0245581 -0.0112335
+ 2.067e+11Hz -0.0245639 -0.0112184
+ 2.068e+11Hz -0.0245698 -0.0112034
+ 2.069e+11Hz -0.0245756 -0.0111885
+ 2.07e+11Hz -0.0245815 -0.0111737
+ 2.071e+11Hz -0.0245874 -0.0111589
+ 2.072e+11Hz -0.0245933 -0.0111442
+ 2.073e+11Hz -0.0245993 -0.0111296
+ 2.074e+11Hz -0.0246052 -0.0111151
+ 2.075e+11Hz -0.0246112 -0.0111006
+ 2.076e+11Hz -0.0246172 -0.0110862
+ 2.077e+11Hz -0.0246233 -0.0110719
+ 2.078e+11Hz -0.0246294 -0.0110577
+ 2.079e+11Hz -0.0246355 -0.0110435
+ 2.08e+11Hz -0.0246417 -0.0110294
+ 2.081e+11Hz -0.0246479 -0.0110154
+ 2.082e+11Hz -0.0246541 -0.0110014
+ 2.083e+11Hz -0.0246604 -0.0109876
+ 2.084e+11Hz -0.0246667 -0.0109738
+ 2.085e+11Hz -0.0246731 -0.01096
+ 2.086e+11Hz -0.0246795 -0.0109464
+ 2.087e+11Hz -0.024686 -0.0109328
+ 2.088e+11Hz -0.0246926 -0.0109192
+ 2.089e+11Hz -0.0246992 -0.0109058
+ 2.09e+11Hz -0.0247058 -0.0108923
+ 2.091e+11Hz -0.0247125 -0.010879
+ 2.092e+11Hz -0.0247193 -0.0108657
+ 2.093e+11Hz -0.0247262 -0.0108525
+ 2.094e+11Hz -0.0247331 -0.0108393
+ 2.095e+11Hz -0.0247401 -0.0108262
+ 2.096e+11Hz -0.0247471 -0.0108132
+ 2.097e+11Hz -0.0247543 -0.0108002
+ 2.098e+11Hz -0.0247615 -0.0107873
+ 2.099e+11Hz -0.0247688 -0.0107744
+ 2.1e+11Hz -0.0247761 -0.0107615
+ 2.101e+11Hz -0.0247836 -0.0107488
+ 2.102e+11Hz -0.0247911 -0.010736
+ 2.103e+11Hz -0.0247988 -0.0107233
+ 2.104e+11Hz -0.0248065 -0.0107107
+ 2.105e+11Hz -0.0248143 -0.0106981
+ 2.106e+11Hz -0.0248222 -0.0106855
+ 2.107e+11Hz -0.0248301 -0.010673
+ 2.108e+11Hz -0.0248382 -0.0106605
+ 2.109e+11Hz -0.0248464 -0.010648
+ 2.11e+11Hz -0.0248547 -0.0106356
+ 2.111e+11Hz -0.0248631 -0.0106232
+ 2.112e+11Hz -0.0248715 -0.0106109
+ 2.113e+11Hz -0.0248801 -0.0105985
+ 2.114e+11Hz -0.0248888 -0.0105862
+ 2.115e+11Hz -0.0248976 -0.0105739
+ 2.116e+11Hz -0.0249065 -0.0105616
+ 2.117e+11Hz -0.0249155 -0.0105494
+ 2.118e+11Hz -0.0249247 -0.0105372
+ 2.119e+11Hz -0.0249339 -0.0105249
+ 2.12e+11Hz -0.0249433 -0.0105127
+ 2.121e+11Hz -0.0249527 -0.0105005
+ 2.122e+11Hz -0.0249623 -0.0104883
+ 2.123e+11Hz -0.024972 -0.0104761
+ 2.124e+11Hz -0.0249819 -0.0104639
+ 2.125e+11Hz -0.0249918 -0.0104517
+ 2.126e+11Hz -0.0250019 -0.0104395
+ 2.127e+11Hz -0.0250121 -0.0104273
+ 2.128e+11Hz -0.0250225 -0.010415
+ 2.129e+11Hz -0.0250329 -0.0104028
+ 2.13e+11Hz -0.0250435 -0.0103905
+ 2.131e+11Hz -0.0250542 -0.0103783
+ 2.132e+11Hz -0.0250651 -0.010366
+ 2.133e+11Hz -0.025076 -0.0103536
+ 2.134e+11Hz -0.0250871 -0.0103413
+ 2.135e+11Hz -0.0250984 -0.0103289
+ 2.136e+11Hz -0.0251098 -0.0103165
+ 2.137e+11Hz -0.0251213 -0.010304
+ 2.138e+11Hz -0.0251329 -0.0102915
+ 2.139e+11Hz -0.0251447 -0.010279
+ 2.14e+11Hz -0.0251566 -0.0102664
+ 2.141e+11Hz -0.0251687 -0.0102538
+ 2.142e+11Hz -0.0251808 -0.0102411
+ 2.143e+11Hz -0.0251932 -0.0102283
+ 2.144e+11Hz -0.0252056 -0.0102155
+ 2.145e+11Hz -0.0252182 -0.0102026
+ 2.146e+11Hz -0.025231 -0.0101897
+ 2.147e+11Hz -0.0252438 -0.0101767
+ 2.148e+11Hz -0.0252569 -0.0101636
+ 2.149e+11Hz -0.02527 -0.0101504
+ 2.15e+11Hz -0.0252833 -0.0101372
+ 2.151e+11Hz -0.0252967 -0.0101239
+ 2.152e+11Hz -0.0253103 -0.0101105
+ 2.153e+11Hz -0.025324 -0.010097
+ 2.154e+11Hz -0.0253378 -0.0100834
+ 2.155e+11Hz -0.0253518 -0.0100697
+ 2.156e+11Hz -0.0253659 -0.0100559
+ 2.157e+11Hz -0.0253802 -0.010042
+ 2.158e+11Hz -0.0253946 -0.010028
+ 2.159e+11Hz -0.0254091 -0.0100139
+ 2.16e+11Hz -0.0254238 -0.00999965
+ 2.161e+11Hz -0.0254385 -0.0099853
+ 2.162e+11Hz -0.0254535 -0.00997083
+ 2.163e+11Hz -0.0254685 -0.00995624
+ 2.164e+11Hz -0.0254837 -0.00994151
+ 2.165e+11Hz -0.025499 -0.00992666
+ 2.166e+11Hz -0.0255145 -0.00991166
+ 2.167e+11Hz -0.02553 -0.00989653
+ 2.168e+11Hz -0.0255457 -0.00988125
+ 2.169e+11Hz -0.0255615 -0.00986583
+ 2.17e+11Hz -0.0255775 -0.00985026
+ 2.171e+11Hz -0.0255935 -0.00983453
+ 2.172e+11Hz -0.0256097 -0.00981864
+ 2.173e+11Hz -0.025626 -0.0098026
+ 2.174e+11Hz -0.0256424 -0.00978639
+ 2.175e+11Hz -0.025659 -0.00977001
+ 2.176e+11Hz -0.0256756 -0.00975347
+ 2.177e+11Hz -0.0256924 -0.00973675
+ 2.178e+11Hz -0.0257093 -0.00971985
+ 2.179e+11Hz -0.0257262 -0.00970276
+ 2.18e+11Hz -0.0257433 -0.0096855
+ 2.181e+11Hz -0.0257605 -0.00966805
+ 2.182e+11Hz -0.0257778 -0.0096504
+ 2.183e+11Hz -0.0257952 -0.00963256
+ 2.184e+11Hz -0.0258126 -0.00961452
+ 2.185e+11Hz -0.0258302 -0.00959629
+ 2.186e+11Hz -0.0258479 -0.00957785
+ 2.187e+11Hz -0.0258656 -0.0095592
+ 2.188e+11Hz -0.0258834 -0.00954034
+ 2.189e+11Hz -0.0259014 -0.00952126
+ 2.19e+11Hz -0.0259194 -0.00950197
+ 2.191e+11Hz -0.0259374 -0.00948247
+ 2.192e+11Hz -0.0259556 -0.00946273
+ 2.193e+11Hz -0.0259738 -0.00944278
+ 2.194e+11Hz -0.0259921 -0.00942259
+ 2.195e+11Hz -0.0260104 -0.00940218
+ 2.196e+11Hz -0.0260288 -0.00938153
+ 2.197e+11Hz -0.0260473 -0.00936064
+ 2.198e+11Hz -0.0260658 -0.00933951
+ 2.199e+11Hz -0.0260844 -0.00931815
+ 2.2e+11Hz -0.026103 -0.00929654
+ 2.201e+11Hz -0.0261217 -0.00927468
+ 2.202e+11Hz -0.0261404 -0.00925257
+ 2.203e+11Hz -0.0261591 -0.00923021
+ 2.204e+11Hz -0.0261779 -0.00920759
+ 2.205e+11Hz -0.0261967 -0.00918472
+ 2.206e+11Hz -0.0262156 -0.00916159
+ 2.207e+11Hz -0.0262344 -0.0091382
+ 2.208e+11Hz -0.0262533 -0.00911455
+ 2.209e+11Hz -0.0262722 -0.00909063
+ 2.21e+11Hz -0.0262911 -0.00906644
+ 2.211e+11Hz -0.0263099 -0.00904199
+ 2.212e+11Hz -0.0263288 -0.00901726
+ 2.213e+11Hz -0.0263477 -0.00899226
+ 2.214e+11Hz -0.0263666 -0.00896699
+ 2.215e+11Hz -0.0263855 -0.00894144
+ 2.216e+11Hz -0.0264044 -0.00891561
+ 2.217e+11Hz -0.0264232 -0.00888951
+ 2.218e+11Hz -0.026442 -0.00886312
+ 2.219e+11Hz -0.0264608 -0.00883645
+ 2.22e+11Hz -0.0264796 -0.0088095
+ 2.221e+11Hz -0.0264983 -0.00878227
+ 2.222e+11Hz -0.0265169 -0.00875475
+ 2.223e+11Hz -0.0265356 -0.00872694
+ 2.224e+11Hz -0.0265541 -0.00869884
+ 2.225e+11Hz -0.0265727 -0.00867046
+ 2.226e+11Hz -0.0265911 -0.00864179
+ 2.227e+11Hz -0.0266095 -0.00861283
+ 2.228e+11Hz -0.0266278 -0.00858358
+ 2.229e+11Hz -0.026646 -0.00855404
+ 2.23e+11Hz -0.0266642 -0.0085242
+ 2.231e+11Hz -0.0266823 -0.00849408
+ 2.232e+11Hz -0.0267003 -0.00846366
+ 2.233e+11Hz -0.0267181 -0.00843296
+ 2.234e+11Hz -0.0267359 -0.00840196
+ 2.235e+11Hz -0.0267536 -0.00837066
+ 2.236e+11Hz -0.0267712 -0.00833908
+ 2.237e+11Hz -0.0267886 -0.0083072
+ 2.238e+11Hz -0.026806 -0.00827504
+ 2.239e+11Hz -0.0268232 -0.00824258
+ 2.24e+11Hz -0.0268402 -0.00820983
+ 2.241e+11Hz -0.0268572 -0.00817679
+ 2.242e+11Hz -0.026874 -0.00814346
+ 2.243e+11Hz -0.0268906 -0.00810984
+ 2.244e+11Hz -0.0269071 -0.00807593
+ 2.245e+11Hz -0.0269235 -0.00804174
+ 2.246e+11Hz -0.0269397 -0.00800726
+ 2.247e+11Hz -0.0269557 -0.0079725
+ 2.248e+11Hz -0.0269716 -0.00793745
+ 2.249e+11Hz -0.0269872 -0.00790212
+ 2.25e+11Hz -0.0270027 -0.00786651
+ 2.251e+11Hz -0.027018 -0.00783062
+ 2.252e+11Hz -0.0270332 -0.00779445
+ 2.253e+11Hz -0.0270481 -0.007758
+ 2.254e+11Hz -0.0270628 -0.00772128
+ 2.255e+11Hz -0.0270773 -0.00768429
+ 2.256e+11Hz -0.0270917 -0.00764702
+ 2.257e+11Hz -0.0271058 -0.00760949
+ 2.258e+11Hz -0.0271196 -0.00757169
+ 2.259e+11Hz -0.0271333 -0.00753363
+ 2.26e+11Hz -0.0271467 -0.0074953
+ 2.261e+11Hz -0.0271599 -0.00745671
+ 2.262e+11Hz -0.0271729 -0.00741787
+ 2.263e+11Hz -0.0271856 -0.00737877
+ 2.264e+11Hz -0.0271981 -0.00733942
+ 2.265e+11Hz -0.0272103 -0.00729982
+ 2.266e+11Hz -0.0272222 -0.00725997
+ 2.267e+11Hz -0.0272339 -0.00721988
+ 2.268e+11Hz -0.0272453 -0.00717955
+ 2.269e+11Hz -0.0272565 -0.00713898
+ 2.27e+11Hz -0.0272674 -0.00709817
+ 2.271e+11Hz -0.027278 -0.00705714
+ 2.272e+11Hz -0.0272883 -0.00701587
+ 2.273e+11Hz -0.0272984 -0.00697438
+ 2.274e+11Hz -0.0273081 -0.00693267
+ 2.275e+11Hz -0.0273176 -0.00689075
+ 2.276e+11Hz -0.0273267 -0.00684861
+ 2.277e+11Hz -0.0273356 -0.00680626
+ 2.278e+11Hz -0.0273441 -0.0067637
+ 2.279e+11Hz -0.0273523 -0.00672094
+ 2.28e+11Hz -0.0273602 -0.00667798
+ 2.281e+11Hz -0.0273678 -0.00663483
+ 2.282e+11Hz -0.0273751 -0.00659148
+ 2.283e+11Hz -0.0273821 -0.00654795
+ 2.284e+11Hz -0.0273887 -0.00650424
+ 2.285e+11Hz -0.027395 -0.00646035
+ 2.286e+11Hz -0.0274009 -0.00641629
+ 2.287e+11Hz -0.0274065 -0.00637206
+ 2.288e+11Hz -0.0274118 -0.00632767
+ 2.289e+11Hz -0.0274167 -0.00628311
+ 2.29e+11Hz -0.0274213 -0.0062384
+ 2.291e+11Hz -0.0274255 -0.00619354
+ 2.292e+11Hz -0.0274294 -0.00614853
+ 2.293e+11Hz -0.0274329 -0.00610338
+ 2.294e+11Hz -0.0274361 -0.0060581
+ 2.295e+11Hz -0.0274388 -0.00601268
+ 2.296e+11Hz -0.0274413 -0.00596714
+ 2.297e+11Hz -0.0274433 -0.00592148
+ 2.298e+11Hz -0.027445 -0.0058757
+ 2.299e+11Hz -0.0274463 -0.00582981
+ 2.3e+11Hz -0.0274472 -0.00578382
+ 2.301e+11Hz -0.0274478 -0.00573772
+ 2.302e+11Hz -0.027448 -0.00569153
+ 2.303e+11Hz -0.0274478 -0.00564524
+ 2.304e+11Hz -0.0274472 -0.00559888
+ 2.305e+11Hz -0.0274462 -0.00555243
+ 2.306e+11Hz -0.0274449 -0.00550591
+ 2.307e+11Hz -0.0274431 -0.00545932
+ 2.308e+11Hz -0.027441 -0.00541266
+ 2.309e+11Hz -0.0274384 -0.00536595
+ 2.31e+11Hz -0.0274355 -0.00531919
+ 2.311e+11Hz -0.0274322 -0.00527237
+ 2.312e+11Hz -0.0274285 -0.00522552
+ 2.313e+11Hz -0.0274244 -0.00517863
+ 2.314e+11Hz -0.0274199 -0.00513171
+ 2.315e+11Hz -0.027415 -0.00508477
+ 2.316e+11Hz -0.0274097 -0.00503781
+ 2.317e+11Hz -0.027404 -0.00499083
+ 2.318e+11Hz -0.0273979 -0.00494384
+ 2.319e+11Hz -0.0273914 -0.00489686
+ 2.32e+11Hz -0.0273845 -0.00484988
+ 2.321e+11Hz -0.0273773 -0.0048029
+ 2.322e+11Hz -0.0273696 -0.00475594
+ 2.323e+11Hz -0.0273615 -0.004709
+ 2.324e+11Hz -0.027353 -0.00466209
+ 2.325e+11Hz -0.0273441 -0.00461521
+ 2.326e+11Hz -0.0273348 -0.00456836
+ 2.327e+11Hz -0.0273251 -0.00452156
+ 2.328e+11Hz -0.027315 -0.00447481
+ 2.329e+11Hz -0.0273045 -0.00442811
+ 2.33e+11Hz -0.0272936 -0.00438147
+ 2.331e+11Hz -0.0272824 -0.0043349
+ 2.332e+11Hz -0.0272707 -0.0042884
+ 2.333e+11Hz -0.0272586 -0.00424197
+ 2.334e+11Hz -0.0272461 -0.00419563
+ 2.335e+11Hz -0.0272333 -0.00414937
+ 2.336e+11Hz -0.02722 -0.00410321
+ 2.337e+11Hz -0.0272064 -0.00405715
+ 2.338e+11Hz -0.0271923 -0.00401119
+ 2.339e+11Hz -0.0271779 -0.00396534
+ 2.34e+11Hz -0.0271631 -0.0039196
+ 2.341e+11Hz -0.0271479 -0.00387399
+ 2.342e+11Hz -0.0271324 -0.0038285
+ 2.343e+11Hz -0.0271164 -0.00378314
+ 2.344e+11Hz -0.0271001 -0.00373791
+ 2.345e+11Hz -0.0270834 -0.00369283
+ 2.346e+11Hz -0.0270663 -0.00364789
+ 2.347e+11Hz -0.0270489 -0.00360311
+ 2.348e+11Hz -0.027031 -0.00355848
+ 2.349e+11Hz -0.0270129 -0.00351401
+ 2.35e+11Hz -0.0269943 -0.00346971
+ 2.351e+11Hz -0.0269754 -0.00342559
+ 2.352e+11Hz -0.0269561 -0.00338163
+ 2.353e+11Hz -0.0269365 -0.00333786
+ 2.354e+11Hz -0.0269165 -0.00329428
+ 2.355e+11Hz -0.0268962 -0.00325088
+ 2.356e+11Hz -0.0268755 -0.00320768
+ 2.357e+11Hz -0.0268545 -0.00316468
+ 2.358e+11Hz -0.0268331 -0.00312188
+ 2.359e+11Hz -0.0268114 -0.0030793
+ 2.36e+11Hz -0.0267894 -0.00303692
+ 2.361e+11Hz -0.026767 -0.00299476
+ 2.362e+11Hz -0.0267443 -0.00295283
+ 2.363e+11Hz -0.0267213 -0.00291112
+ 2.364e+11Hz -0.026698 -0.00286964
+ 2.365e+11Hz -0.0266743 -0.00282839
+ 2.366e+11Hz -0.0266503 -0.00278739
+ 2.367e+11Hz -0.0266261 -0.00274662
+ 2.368e+11Hz -0.0266015 -0.0027061
+ 2.369e+11Hz -0.0265766 -0.00266583
+ 2.37e+11Hz -0.0265514 -0.00262581
+ 2.371e+11Hz -0.0265259 -0.00258605
+ 2.372e+11Hz -0.0265002 -0.00254655
+ 2.373e+11Hz -0.0264741 -0.00250732
+ 2.374e+11Hz -0.0264478 -0.00246835
+ 2.375e+11Hz -0.0264212 -0.00242965
+ 2.376e+11Hz -0.0263943 -0.00239123
+ 2.377e+11Hz -0.0263671 -0.00235308
+ 2.378e+11Hz -0.0263397 -0.00231521
+ 2.379e+11Hz -0.026312 -0.00227762
+ 2.38e+11Hz -0.0262841 -0.00224033
+ 2.381e+11Hz -0.0262559 -0.00220331
+ 2.382e+11Hz -0.0262275 -0.00216659
+ 2.383e+11Hz -0.0261988 -0.00213017
+ 2.384e+11Hz -0.0261699 -0.00209404
+ 2.385e+11Hz -0.0261408 -0.00205821
+ 2.386e+11Hz -0.0261114 -0.00202268
+ 2.387e+11Hz -0.0260818 -0.00198746
+ 2.388e+11Hz -0.026052 -0.00195254
+ 2.389e+11Hz -0.0260219 -0.00191792
+ 2.39e+11Hz -0.0259917 -0.00188362
+ 2.391e+11Hz -0.0259613 -0.00184963
+ 2.392e+11Hz -0.0259306 -0.00181595
+ 2.393e+11Hz -0.0258998 -0.00178259
+ 2.394e+11Hz -0.0258687 -0.00174955
+ 2.395e+11Hz -0.0258375 -0.00171682
+ 2.396e+11Hz -0.0258061 -0.00168442
+ 2.397e+11Hz -0.0257746 -0.00165234
+ 2.398e+11Hz -0.0257428 -0.00162058
+ 2.399e+11Hz -0.0257109 -0.00158914
+ 2.4e+11Hz -0.0256788 -0.00155803
+ 2.401e+11Hz -0.0256466 -0.00152724
+ 2.402e+11Hz -0.0256142 -0.00149679
+ 2.403e+11Hz -0.0255817 -0.00146666
+ 2.404e+11Hz -0.025549 -0.00143686
+ 2.405e+11Hz -0.0255162 -0.00140739
+ 2.406e+11Hz -0.0254833 -0.00137825
+ 2.407e+11Hz -0.0254502 -0.00134944
+ 2.408e+11Hz -0.025417 -0.00132096
+ 2.409e+11Hz -0.0253837 -0.00129281
+ 2.41e+11Hz -0.0253503 -0.001265
+ 2.411e+11Hz -0.0253168 -0.00123752
+ 2.412e+11Hz -0.0252831 -0.00121037
+ 2.413e+11Hz -0.0252494 -0.00118355
+ 2.414e+11Hz -0.0252156 -0.00115707
+ 2.415e+11Hz -0.0251817 -0.00113092
+ 2.416e+11Hz -0.0251477 -0.0011051
+ 2.417e+11Hz -0.0251136 -0.00107961
+ 2.418e+11Hz -0.0250794 -0.00105445
+ 2.419e+11Hz -0.0250452 -0.00102962
+ 2.42e+11Hz -0.0250109 -0.00100513
+ 2.421e+11Hz -0.0249766 -0.000980965
+ 2.422e+11Hz -0.0249422 -0.000957129
+ 2.423e+11Hz -0.0249077 -0.000933622
+ 2.424e+11Hz -0.0248732 -0.000910443
+ 2.425e+11Hz -0.0248386 -0.00088759
+ 2.426e+11Hz -0.024804 -0.000865064
+ 2.427e+11Hz -0.0247694 -0.000842863
+ 2.428e+11Hz -0.0247347 -0.000820986
+ 2.429e+11Hz -0.0247001 -0.000799432
+ 2.43e+11Hz -0.0246653 -0.000778199
+ 2.431e+11Hz -0.0246306 -0.000757287
+ 2.432e+11Hz -0.0245959 -0.000736694
+ 2.433e+11Hz -0.0245611 -0.000716418
+ 2.434e+11Hz -0.0245264 -0.000696459
+ 2.435e+11Hz -0.0244916 -0.000676815
+ 2.436e+11Hz -0.0244568 -0.000657484
+ 2.437e+11Hz -0.0244221 -0.000638464
+ 2.438e+11Hz -0.0243873 -0.000619755
+ 2.439e+11Hz -0.0243526 -0.000601353
+ 2.44e+11Hz -0.0243179 -0.000583258
+ 2.441e+11Hz -0.0242832 -0.000565468
+ 2.442e+11Hz -0.0242485 -0.000547981
+ 2.443e+11Hz -0.0242139 -0.000530794
+ 2.444e+11Hz -0.0241793 -0.000513906
+ 2.445e+11Hz -0.0241447 -0.000497316
+ 2.446e+11Hz -0.0241101 -0.00048102
+ 2.447e+11Hz -0.0240756 -0.000465017
+ 2.448e+11Hz -0.0240412 -0.000449304
+ 2.449e+11Hz -0.0240068 -0.00043388
+ 2.45e+11Hz -0.0239724 -0.000418742
+ 2.451e+11Hz -0.0239381 -0.000403888
+ 2.452e+11Hz -0.0239039 -0.000389316
+ 2.453e+11Hz -0.0238697 -0.000375023
+ 2.454e+11Hz -0.0238356 -0.000361008
+ 2.455e+11Hz -0.0238015 -0.000347267
+ 2.456e+11Hz -0.0237676 -0.000333798
+ 2.457e+11Hz -0.0237337 -0.0003206
+ 2.458e+11Hz -0.0236998 -0.000307669
+ 2.459e+11Hz -0.0236661 -0.000295002
+ 2.46e+11Hz -0.0236324 -0.000282599
+ 2.461e+11Hz -0.0235988 -0.000270455
+ 2.462e+11Hz -0.0235653 -0.000258569
+ 2.463e+11Hz -0.0235319 -0.000246937
+ 2.464e+11Hz -0.0234985 -0.000235558
+ 2.465e+11Hz -0.0234653 -0.000224429
+ 2.466e+11Hz -0.0234321 -0.000213547
+ 2.467e+11Hz -0.0233991 -0.000202909
+ 2.468e+11Hz -0.0233662 -0.000192513
+ 2.469e+11Hz -0.0233333 -0.000182357
+ 2.47e+11Hz -0.0233006 -0.000172437
+ 2.471e+11Hz -0.0232679 -0.000162751
+ 2.472e+11Hz -0.0232354 -0.000153296
+ 2.473e+11Hz -0.023203 -0.00014407
+ 2.474e+11Hz -0.0231706 -0.00013507
+ 2.475e+11Hz -0.0231384 -0.000126293
+ 2.476e+11Hz -0.0231063 -0.000117737
+ 2.477e+11Hz -0.0230744 -0.000109399
+ 2.478e+11Hz -0.0230425 -0.000101277
+ 2.479e+11Hz -0.0230108 -9.33669e-05
+ 2.48e+11Hz -0.0229792 -8.5667e-05
+ 2.481e+11Hz -0.0229477 -7.81745e-05
+ 2.482e+11Hz -0.0229163 -7.08868e-05
+ 2.483e+11Hz -0.022885 -6.38012e-05
+ 2.484e+11Hz -0.0228539 -5.6915e-05
+ 2.485e+11Hz -0.0228229 -5.02257e-05
+ 2.486e+11Hz -0.0227921 -4.37307e-05
+ 2.487e+11Hz -0.0227613 -3.74273e-05
+ 2.488e+11Hz -0.0227307 -3.13131e-05
+ 2.489e+11Hz -0.0227002 -2.53853e-05
+ 2.49e+11Hz -0.0226699 -1.96415e-05
+ 2.491e+11Hz -0.0226397 -1.4079e-05
+ 2.492e+11Hz -0.0226096 -8.69551e-06
+ 2.493e+11Hz -0.0225796 -3.48836e-06
+ 2.494e+11Hz -0.0225498 1.5449e-06
+ 2.495e+11Hz -0.0225202 6.40676e-06
+ 2.496e+11Hz -0.0224906 1.10997e-05
+ 2.497e+11Hz -0.0224612 1.5626e-05
+ 2.498e+11Hz -0.022432 1.99883e-05
+ 2.499e+11Hz -0.0224029 2.41889e-05
+ 2.5e+11Hz -0.0223739 2.82301e-05
+ 2.501e+11Hz -0.022345 3.21144e-05
+ 2.502e+11Hz -0.0223163 3.5844e-05
+ 2.503e+11Hz -0.0222878 3.94213e-05
+ 2.504e+11Hz -0.0222594 4.28485e-05
+ 2.505e+11Hz -0.0222311 4.61279e-05
+ 2.506e+11Hz -0.022203 4.92618e-05
+ 2.507e+11Hz -0.022175 5.22523e-05
+ 2.508e+11Hz -0.0221471 5.51017e-05
+ 2.509e+11Hz -0.0221194 5.78121e-05
+ 2.51e+11Hz -0.0220919 6.03856e-05
+ 2.511e+11Hz -0.0220645 6.28245e-05
+ 2.512e+11Hz -0.0220372 6.51306e-05
+ 2.513e+11Hz -0.0220101 6.73063e-05
+ 2.514e+11Hz -0.0219831 6.93533e-05
+ 2.515e+11Hz -0.0219563 7.12739e-05
+ 2.516e+11Hz -0.0219296 7.307e-05
+ 2.517e+11Hz -0.0219031 7.47435e-05
+ 2.518e+11Hz -0.0218767 7.62963e-05
+ 2.519e+11Hz -0.0218505 7.77305e-05
+ 2.52e+11Hz -0.0218244 7.90478e-05
+ 2.521e+11Hz -0.0217984 8.02503e-05
+ 2.522e+11Hz -0.0217726 8.13396e-05
+ 2.523e+11Hz -0.021747 8.23176e-05
+ 2.524e+11Hz -0.0217215 8.31861e-05
+ 2.525e+11Hz -0.0216961 8.39469e-05
+ 2.526e+11Hz -0.0216709 8.46017e-05
+ 2.527e+11Hz -0.0216458 8.51522e-05
+ 2.528e+11Hz -0.0216209 8.56002e-05
+ 2.529e+11Hz -0.0215961 8.59473e-05
+ 2.53e+11Hz -0.0215715 8.61952e-05
+ 2.531e+11Hz -0.021547 8.63456e-05
+ 2.532e+11Hz -0.0215227 8.63999e-05
+ 2.533e+11Hz -0.0214985 8.63598e-05
+ 2.534e+11Hz -0.0214745 8.6227e-05
+ 2.535e+11Hz -0.0214506 8.60029e-05
+ 2.536e+11Hz -0.0214269 8.56891e-05
+ 2.537e+11Hz -0.0214033 8.52871e-05
+ 2.538e+11Hz -0.0213798 8.47985e-05
+ 2.539e+11Hz -0.0213565 8.42246e-05
+ 2.54e+11Hz -0.0213334 8.3567e-05
+ 2.541e+11Hz -0.0213104 8.28271e-05
+ 2.542e+11Hz -0.0212875 8.20064e-05
+ 2.543e+11Hz -0.0212648 8.11063e-05
+ 2.544e+11Hz -0.0212423 8.01282e-05
+ 2.545e+11Hz -0.0212199 7.90735e-05
+ 2.546e+11Hz -0.0211976 7.79437e-05
+ 2.547e+11Hz -0.0211755 7.674e-05
+ 2.548e+11Hz -0.0211536 7.54639e-05
+ 2.549e+11Hz -0.0211318 7.41168e-05
+ 2.55e+11Hz -0.0211101 7.26999e-05
+ 2.551e+11Hz -0.0210886 7.12146e-05
+ 2.552e+11Hz -0.0210673 6.96624e-05
+ 2.553e+11Hz -0.0210461 6.80445e-05
+ 2.554e+11Hz -0.021025 6.63622e-05
+ 2.555e+11Hz -0.0210041 6.4617e-05
+ 2.556e+11Hz -0.0209833 6.28101e-05
+ 2.557e+11Hz -0.0209627 6.09428e-05
+ 2.558e+11Hz -0.0209423 5.90166e-05
+ 2.559e+11Hz -0.020922 5.70326e-05
+ 2.56e+11Hz -0.0209018 5.49924e-05
+ 2.561e+11Hz -0.0208818 5.28972e-05
+ 2.562e+11Hz -0.020862 5.07483e-05
+ 2.563e+11Hz -0.0208423 4.85471e-05
+ 2.564e+11Hz -0.0208228 4.62949e-05
+ 2.565e+11Hz -0.0208034 4.39932e-05
+ 2.566e+11Hz -0.0207841 4.16432e-05
+ 2.567e+11Hz -0.0207651 3.92464e-05
+ 2.568e+11Hz -0.0207461 3.68041e-05
+ 2.569e+11Hz -0.0207274 3.43178e-05
+ 2.57e+11Hz -0.0207088 3.17889e-05
+ 2.571e+11Hz -0.0206903 2.92187e-05
+ 2.572e+11Hz -0.020672 2.66087e-05
+ 2.573e+11Hz -0.0206538 2.39604e-05
+ 2.574e+11Hz -0.0206359 2.12753e-05
+ 2.575e+11Hz -0.020618 1.85547e-05
+ 2.576e+11Hz -0.0206004 1.58003e-05
+ 2.577e+11Hz -0.0205828 1.30135e-05
+ 2.578e+11Hz -0.0205655 1.0196e-05
+ 2.579e+11Hz -0.0205483 7.34912e-06
+ 2.58e+11Hz -0.0205312 4.47462e-06
+ 2.581e+11Hz -0.0205144 1.57405e-06
+ 2.582e+11Hz -0.0204976 -1.35096e-06
+ 2.583e+11Hz -0.0204811 -4.29876e-06
+ 2.584e+11Hz -0.0204647 -7.26767e-06
+ 2.585e+11Hz -0.0204485 -1.0256e-05
+ 2.586e+11Hz -0.0204324 -1.3262e-05
+ 2.587e+11Hz -0.0204165 -1.6284e-05
+ 2.588e+11Hz -0.0204007 -1.93201e-05
+ 2.589e+11Hz -0.0203852 -2.23686e-05
+ 2.59e+11Hz -0.0203697 -2.54275e-05
+ 2.591e+11Hz -0.0203545 -2.84952e-05
+ 2.592e+11Hz -0.0203394 -3.15696e-05
+ 2.593e+11Hz -0.0203245 -3.46488e-05
+ 2.594e+11Hz -0.0203097 -3.77309e-05
+ 2.595e+11Hz -0.0202951 -4.08139e-05
+ 2.596e+11Hz -0.0202807 -4.38958e-05
+ 2.597e+11Hz -0.0202665 -4.69745e-05
+ 2.598e+11Hz -0.0202524 -5.00479e-05
+ 2.599e+11Hz -0.0202385 -5.3114e-05
+ 2.6e+11Hz -0.0202247 -5.61705e-05
+ 2.601e+11Hz -0.0202112 -5.92153e-05
+ 2.602e+11Hz -0.0201977 -6.22462e-05
+ 2.603e+11Hz -0.0201845 -6.5261e-05
+ 2.604e+11Hz -0.0201714 -6.82573e-05
+ 2.605e+11Hz -0.0201585 -7.12328e-05
+ 2.606e+11Hz -0.0201458 -7.41852e-05
+ 2.607e+11Hz -0.0201333 -7.71121e-05
+ 2.608e+11Hz -0.0201209 -8.00111e-05
+ 2.609e+11Hz -0.0201087 -8.28796e-05
+ 2.61e+11Hz -0.0200966 -8.57153e-05
+ 2.611e+11Hz -0.0200848 -8.85157e-05
+ 2.612e+11Hz -0.0200731 -9.1278e-05
+ 2.613e+11Hz -0.0200616 -9.39998e-05
+ 2.614e+11Hz -0.0200502 -9.66785e-05
+ 2.615e+11Hz -0.020039 -9.93113e-05
+ 2.616e+11Hz -0.020028 -0.000101896
+ 2.617e+11Hz -0.0200172 -0.000104429
+ 2.618e+11Hz -0.0200065 -0.000106908
+ 2.619e+11Hz -0.019996 -0.00010933
+ 2.62e+11Hz -0.0199857 -0.000111693
+ 2.621e+11Hz -0.0199756 -0.000113993
+ 2.622e+11Hz -0.0199656 -0.000116228
+ 2.623e+11Hz -0.0199558 -0.000118394
+ 2.624e+11Hz -0.0199462 -0.00012049
+ 2.625e+11Hz -0.0199367 -0.000122511
+ 2.626e+11Hz -0.0199274 -0.000124455
+ 2.627e+11Hz -0.0199183 -0.000126319
+ 2.628e+11Hz -0.0199094 -0.0001281
+ 2.629e+11Hz -0.0199006 -0.000129794
+ 2.63e+11Hz -0.019892 -0.000131399
+ 2.631e+11Hz -0.0198835 -0.000132912
+ 2.632e+11Hz -0.0198753 -0.000134329
+ 2.633e+11Hz -0.0198672 -0.000135647
+ 2.634e+11Hz -0.0198592 -0.000136863
+ 2.635e+11Hz -0.0198514 -0.000137973
+ 2.636e+11Hz -0.0198438 -0.000138976
+ 2.637e+11Hz -0.0198364 -0.000139866
+ 2.638e+11Hz -0.0198291 -0.000140642
+ 2.639e+11Hz -0.0198219 -0.0001413
+ 2.64e+11Hz -0.0198149 -0.000141836
+ 2.641e+11Hz -0.0198081 -0.000142247
+ 2.642e+11Hz -0.0198015 -0.00014253
+ 2.643e+11Hz -0.019795 -0.000142682
+ 2.644e+11Hz -0.0197886 -0.000142699
+ 2.645e+11Hz -0.0197824 -0.000142578
+ 2.646e+11Hz -0.0197764 -0.000142315
+ 2.647e+11Hz -0.0197705 -0.000141908
+ 2.648e+11Hz -0.0197647 -0.000141353
+ 2.649e+11Hz -0.0197591 -0.000140646
+ 2.65e+11Hz -0.0197536 -0.000139785
+ 2.651e+11Hz -0.0197483 -0.000138766
+ 2.652e+11Hz -0.0197431 -0.000137585
+ 2.653e+11Hz -0.0197381 -0.00013624
+ 2.654e+11Hz -0.0197332 -0.000134726
+ 2.655e+11Hz -0.0197284 -0.000133042
+ 2.656e+11Hz -0.0197237 -0.000131182
+ 2.657e+11Hz -0.0197192 -0.000129145
+ 2.658e+11Hz -0.0197148 -0.000126927
+ 2.659e+11Hz -0.0197105 -0.000124524
+ 2.66e+11Hz -0.0197064 -0.000121934
+ 2.661e+11Hz -0.0197023 -0.000119153
+ 2.662e+11Hz -0.0196984 -0.000116178
+ 2.663e+11Hz -0.0196946 -0.000113006
+ 2.664e+11Hz -0.0196909 -0.000109633
+ 2.665e+11Hz -0.0196873 -0.000106058
+ 2.666e+11Hz -0.0196838 -0.000102276
+ 2.667e+11Hz -0.0196804 -9.82843e-05
+ 2.668e+11Hz -0.0196771 -9.40805e-05
+ 2.669e+11Hz -0.0196739 -8.96614e-05
+ 2.67e+11Hz -0.0196708 -8.5024e-05
+ 2.671e+11Hz -0.0196678 -8.01655e-05
+ 2.672e+11Hz -0.0196648 -7.5083e-05
+ 2.673e+11Hz -0.019662 -6.97738e-05
+ 2.674e+11Hz -0.0196592 -6.42351e-05
+ 2.675e+11Hz -0.0196564 -5.84643e-05
+ 2.676e+11Hz -0.0196538 -5.24586e-05
+ 2.677e+11Hz -0.0196512 -4.62156e-05
+ 2.678e+11Hz -0.0196486 -3.97327e-05
+ 2.679e+11Hz -0.0196462 -3.30074e-05
+ 2.68e+11Hz -0.0196437 -2.60373e-05
+ 2.681e+11Hz -0.0196413 -1.88202e-05
+ 2.682e+11Hz -0.019639 -1.13536e-05
+ 2.683e+11Hz -0.0196367 -3.63541e-06
+ 2.684e+11Hz -0.0196344 4.33653e-06
+ 2.685e+11Hz -0.0196322 1.25643e-05
+ 2.686e+11Hz -0.01963 2.10499e-05
+ 2.687e+11Hz -0.0196278 2.97953e-05
+ 2.688e+11Hz -0.0196256 3.88023e-05
+ 2.689e+11Hz -0.0196234 4.80727e-05
+ 2.69e+11Hz -0.0196212 5.76082e-05
+ 2.691e+11Hz -0.0196191 6.74105e-05
+ 2.692e+11Hz -0.0196169 7.74809e-05
+ 2.693e+11Hz -0.0196147 8.78211e-05
+ 2.694e+11Hz -0.0196125 9.84323e-05
+ 2.695e+11Hz -0.0196103 0.000109316
+ 2.696e+11Hz -0.019608 0.000120473
+ 2.697e+11Hz -0.0196058 0.000131905
+ 2.698e+11Hz -0.0196035 0.000143612
+ 2.699e+11Hz -0.0196011 0.000155596
+ 2.7e+11Hz -0.0195987 0.000167857
+ 2.701e+11Hz -0.0195962 0.000180396
+ 2.702e+11Hz -0.0195937 0.000193214
+ 2.703e+11Hz -0.0195912 0.00020631
+ 2.704e+11Hz -0.0195885 0.000219687
+ 2.705e+11Hz -0.0195858 0.000233343
+ 2.706e+11Hz -0.019583 0.000247279
+ 2.707e+11Hz -0.0195801 0.000261495
+ 2.708e+11Hz -0.0195771 0.000275991
+ 2.709e+11Hz -0.0195741 0.000290768
+ 2.71e+11Hz -0.0195709 0.000305823
+ 2.711e+11Hz -0.0195676 0.000321159
+ 2.712e+11Hz -0.0195642 0.000336773
+ 2.713e+11Hz -0.0195607 0.000352665
+ 2.714e+11Hz -0.019557 0.000368835
+ 2.715e+11Hz -0.0195532 0.000385281
+ 2.716e+11Hz -0.0195493 0.000402004
+ 2.717e+11Hz -0.0195453 0.000419001
+ 2.718e+11Hz -0.019541 0.000436272
+ 2.719e+11Hz -0.0195367 0.000453815
+ 2.72e+11Hz -0.0195321 0.000471629
+ 2.721e+11Hz -0.0195274 0.000489712
+ 2.722e+11Hz -0.0195226 0.000508063
+ 2.723e+11Hz -0.0195175 0.00052668
+ 2.724e+11Hz -0.0195123 0.000545561
+ 2.725e+11Hz -0.0195069 0.000564704
+ 2.726e+11Hz -0.0195012 0.000584106
+ 2.727e+11Hz -0.0194954 0.000603767
+ 2.728e+11Hz -0.0194894 0.000623682
+ 2.729e+11Hz -0.0194831 0.000643851
+ 2.73e+11Hz -0.0194766 0.000664269
+ 2.731e+11Hz -0.0194699 0.000684935
+ 2.732e+11Hz -0.019463 0.000705845
+ 2.733e+11Hz -0.0194558 0.000726996
+ 2.734e+11Hz -0.0194484 0.000748386
+ 2.735e+11Hz -0.0194408 0.000770011
+ 2.736e+11Hz -0.0194329 0.000791868
+ 2.737e+11Hz -0.0194247 0.000813953
+ 2.738e+11Hz -0.0194162 0.000836262
+ 2.739e+11Hz -0.0194075 0.000858792
+ 2.74e+11Hz -0.0193985 0.000881539
+ 2.741e+11Hz -0.0193893 0.000904499
+ 2.742e+11Hz -0.0193797 0.000927668
+ 2.743e+11Hz -0.0193699 0.000951042
+ 2.744e+11Hz -0.0193597 0.000974616
+ 2.745e+11Hz -0.0193493 0.000998386
+ 2.746e+11Hz -0.0193385 0.00102235
+ 2.747e+11Hz -0.0193275 0.0010465
+ 2.748e+11Hz -0.0193161 0.00107083
+ 2.749e+11Hz -0.0193044 0.00109533
+ 2.75e+11Hz -0.0192923 0.00112001
+ 2.751e+11Hz -0.01928 0.00114486
+ 2.752e+11Hz -0.0192673 0.00116986
+ 2.753e+11Hz -0.0192542 0.00119503
+ 2.754e+11Hz -0.0192409 0.00122034
+ 2.755e+11Hz -0.0192271 0.0012458
+ 2.756e+11Hz -0.019213 0.0012714
+ 2.757e+11Hz -0.0191986 0.00129713
+ 2.758e+11Hz -0.0191838 0.00132299
+ 2.759e+11Hz -0.0191686 0.00134898
+ 2.76e+11Hz -0.0191531 0.00137508
+ 2.761e+11Hz -0.0191372 0.00140129
+ 2.762e+11Hz -0.0191209 0.0014276
+ 2.763e+11Hz -0.0191042 0.00145401
+ 2.764e+11Hz -0.0190872 0.00148051
+ 2.765e+11Hz -0.0190698 0.0015071
+ 2.766e+11Hz -0.0190519 0.00153376
+ 2.767e+11Hz -0.0190337 0.0015605
+ 2.768e+11Hz -0.0190151 0.0015873
+ 2.769e+11Hz -0.0189961 0.00161415
+ 2.77e+11Hz -0.0189767 0.00164106
+ 2.771e+11Hz -0.0189569 0.00166802
+ 2.772e+11Hz -0.0189367 0.001695
+ 2.773e+11Hz -0.0189161 0.00172202
+ 2.774e+11Hz -0.018895 0.00174907
+ 2.775e+11Hz -0.0188736 0.00177613
+ 2.776e+11Hz -0.0188518 0.00180319
+ 2.777e+11Hz -0.0188295 0.00183026
+ 2.778e+11Hz -0.0188068 0.00185732
+ 2.779e+11Hz -0.0187837 0.00188437
+ 2.78e+11Hz -0.0187602 0.0019114
+ 2.781e+11Hz -0.0187363 0.0019384
+ 2.782e+11Hz -0.0187119 0.00196536
+ 2.783e+11Hz -0.0186871 0.00199228
+ 2.784e+11Hz -0.0186619 0.00201915
+ 2.785e+11Hz -0.0186363 0.00204596
+ 2.786e+11Hz -0.0186103 0.0020727
+ 2.787e+11Hz -0.0185838 0.00209937
+ 2.788e+11Hz -0.0185569 0.00212596
+ 2.789e+11Hz -0.0185296 0.00215246
+ 2.79e+11Hz -0.0185019 0.00217886
+ 2.791e+11Hz -0.0184737 0.00220516
+ 2.792e+11Hz -0.0184451 0.00223134
+ 2.793e+11Hz -0.0184161 0.00225741
+ 2.794e+11Hz -0.0183867 0.00228334
+ 2.795e+11Hz -0.0183569 0.00230914
+ 2.796e+11Hz -0.0183266 0.0023348
+ 2.797e+11Hz -0.018296 0.00236031
+ 2.798e+11Hz -0.0182649 0.00238565
+ 2.799e+11Hz -0.0182334 0.00241084
+ 2.8e+11Hz -0.0182015 0.00243584
+ 2.801e+11Hz -0.0181691 0.00246067
+ 2.802e+11Hz -0.0181364 0.0024853
+ 2.803e+11Hz -0.0181033 0.00250974
+ 2.804e+11Hz -0.0180698 0.00253398
+ 2.805e+11Hz -0.0180358 0.002558
+ 2.806e+11Hz -0.0180015 0.00258181
+ 2.807e+11Hz -0.0179668 0.00260538
+ 2.808e+11Hz -0.0179317 0.00262873
+ 2.809e+11Hz -0.0178962 0.00265183
+ 2.81e+11Hz -0.0178603 0.00267468
+ 2.811e+11Hz -0.017824 0.00269728
+ 2.812e+11Hz -0.0177874 0.00271962
+ 2.813e+11Hz -0.0177504 0.00274168
+ 2.814e+11Hz -0.017713 0.00276347
+ 2.815e+11Hz -0.0176752 0.00278497
+ 2.816e+11Hz -0.0176371 0.00280619
+ 2.817e+11Hz -0.0175986 0.0028271
+ 2.818e+11Hz -0.0175598 0.00284772
+ 2.819e+11Hz -0.0175207 0.00286802
+ 2.82e+11Hz -0.0174811 0.002888
+ 2.821e+11Hz -0.0174413 0.00290766
+ 2.822e+11Hz -0.0174011 0.00292699
+ 2.823e+11Hz -0.0173606 0.00294599
+ 2.824e+11Hz -0.0173198 0.00296464
+ 2.825e+11Hz -0.0172786 0.00298294
+ 2.826e+11Hz -0.0172372 0.00300089
+ 2.827e+11Hz -0.0171954 0.00301848
+ 2.828e+11Hz -0.0171533 0.0030357
+ 2.829e+11Hz -0.017111 0.00305255
+ 2.83e+11Hz -0.0170683 0.00306903
+ 2.831e+11Hz -0.0170254 0.00308512
+ 2.832e+11Hz -0.0169822 0.00310083
+ 2.833e+11Hz -0.0169388 0.00311614
+ 2.834e+11Hz -0.016895 0.00313105
+ 2.835e+11Hz -0.016851 0.00314556
+ 2.836e+11Hz -0.0168068 0.00315967
+ 2.837e+11Hz -0.0167623 0.00317336
+ 2.838e+11Hz -0.0167176 0.00318664
+ 2.839e+11Hz -0.0166727 0.0031995
+ 2.84e+11Hz -0.0166275 0.00321193
+ 2.841e+11Hz -0.0165821 0.00322393
+ 2.842e+11Hz -0.0165366 0.0032355
+ 2.843e+11Hz -0.0164908 0.00324664
+ 2.844e+11Hz -0.0164448 0.00325733
+ 2.845e+11Hz -0.0163986 0.00326758
+ 2.846e+11Hz -0.0163523 0.00327739
+ 2.847e+11Hz -0.0163058 0.00328674
+ 2.848e+11Hz -0.0162591 0.00329564
+ 2.849e+11Hz -0.0162123 0.00330409
+ 2.85e+11Hz -0.0161653 0.00331208
+ 2.851e+11Hz -0.0161182 0.00331961
+ 2.852e+11Hz -0.016071 0.00332667
+ 2.853e+11Hz -0.0160236 0.00333327
+ 2.854e+11Hz -0.0159762 0.0033394
+ 2.855e+11Hz -0.0159286 0.00334506
+ 2.856e+11Hz -0.0158809 0.00335025
+ 2.857e+11Hz -0.0158331 0.00335497
+ 2.858e+11Hz -0.0157853 0.00335922
+ 2.859e+11Hz -0.0157373 0.00336299
+ 2.86e+11Hz -0.0156893 0.00336628
+ 2.861e+11Hz -0.0156413 0.0033691
+ 2.862e+11Hz -0.0155932 0.00337144
+ 2.863e+11Hz -0.015545 0.0033733
+ 2.864e+11Hz -0.0154969 0.00337469
+ 2.865e+11Hz -0.0154487 0.00337559
+ 2.866e+11Hz -0.0154004 0.00337602
+ 2.867e+11Hz -0.0153522 0.00337596
+ 2.868e+11Hz -0.015304 0.00337543
+ 2.869e+11Hz -0.0152558 0.00337442
+ 2.87e+11Hz -0.0152075 0.00337293
+ 2.871e+11Hz -0.0151594 0.00337097
+ 2.872e+11Hz -0.0151112 0.00336853
+ 2.873e+11Hz -0.0150631 0.00336562
+ 2.874e+11Hz -0.015015 0.00336223
+ 2.875e+11Hz -0.014967 0.00335837
+ 2.876e+11Hz -0.014919 0.00335404
+ 2.877e+11Hz -0.0148712 0.00334925
+ 2.878e+11Hz -0.0148234 0.00334398
+ 2.879e+11Hz -0.0147756 0.00333825
+ 2.88e+11Hz -0.014728 0.00333206
+ 2.881e+11Hz -0.0146805 0.00332541
+ 2.882e+11Hz -0.0146331 0.0033183
+ 2.883e+11Hz -0.0145858 0.00331074
+ 2.884e+11Hz -0.0145386 0.00330273
+ 2.885e+11Hz -0.0144916 0.00329427
+ 2.886e+11Hz -0.0144447 0.00328536
+ 2.887e+11Hz -0.014398 0.003276
+ 2.888e+11Hz -0.0143514 0.00326621
+ 2.889e+11Hz -0.0143049 0.00325599
+ 2.89e+11Hz -0.0142587 0.00324533
+ 2.891e+11Hz -0.0142126 0.00323425
+ 2.892e+11Hz -0.0141666 0.00322274
+ 2.893e+11Hz -0.0141209 0.00321081
+ 2.894e+11Hz -0.0140754 0.00319846
+ 2.895e+11Hz -0.0140301 0.0031857
+ 2.896e+11Hz -0.0139849 0.00317254
+ 2.897e+11Hz -0.01394 0.00315898
+ 2.898e+11Hz -0.0138954 0.00314501
+ 2.899e+11Hz -0.0138509 0.00313066
+ 2.9e+11Hz -0.0138067 0.00311591
+ 2.901e+11Hz -0.0137627 0.00310079
+ 2.902e+11Hz -0.0137189 0.00308528
+ 2.903e+11Hz -0.0136754 0.0030694
+ 2.904e+11Hz -0.0136322 0.00305316
+ 2.905e+11Hz -0.0135892 0.00303656
+ 2.906e+11Hz -0.0135465 0.00301959
+ 2.907e+11Hz -0.0135041 0.00300228
+ 2.908e+11Hz -0.0134619 0.00298463
+ 2.909e+11Hz -0.01342 0.00296663
+ 2.91e+11Hz -0.0133784 0.0029483
+ 2.911e+11Hz -0.0133371 0.00292965
+ 2.912e+11Hz -0.013296 0.00291067
+ 2.913e+11Hz -0.0132553 0.00289138
+ 2.914e+11Hz -0.0132149 0.00287178
+ 2.915e+11Hz -0.0131748 0.00285188
+ 2.916e+11Hz -0.013135 0.00283168
+ 2.917e+11Hz -0.0130955 0.0028112
+ 2.918e+11Hz -0.0130563 0.00279043
+ 2.919e+11Hz -0.0130175 0.00276938
+ 2.92e+11Hz -0.0129789 0.00274806
+ 2.921e+11Hz -0.0129407 0.00272648
+ 2.922e+11Hz -0.0129029 0.00270464
+ 2.923e+11Hz -0.0128653 0.00268255
+ 2.924e+11Hz -0.0128281 0.00266022
+ 2.925e+11Hz -0.0127913 0.00263765
+ 2.926e+11Hz -0.0127547 0.00261485
+ 2.927e+11Hz -0.0127186 0.00259183
+ 2.928e+11Hz -0.0126827 0.00256859
+ 2.929e+11Hz -0.0126472 0.00254514
+ 2.93e+11Hz -0.0126121 0.00252149
+ 2.931e+11Hz -0.0125773 0.00249764
+ 2.932e+11Hz -0.0125429 0.0024736
+ 2.933e+11Hz -0.0125088 0.00244938
+ 2.934e+11Hz -0.012475 0.00242498
+ 2.935e+11Hz -0.0124417 0.00240041
+ 2.936e+11Hz -0.0124087 0.00237569
+ 2.937e+11Hz -0.012376 0.0023508
+ 2.938e+11Hz -0.0123437 0.00232577
+ 2.939e+11Hz -0.0123117 0.00230059
+ 2.94e+11Hz -0.0122801 0.00227528
+ 2.941e+11Hz -0.0122489 0.00224984
+ 2.942e+11Hz -0.012218 0.00222428
+ 2.943e+11Hz -0.0121875 0.00219861
+ 2.944e+11Hz -0.0121574 0.00217282
+ 2.945e+11Hz -0.0121276 0.00214693
+ 2.946e+11Hz -0.0120981 0.00212095
+ 2.947e+11Hz -0.012069 0.00209488
+ 2.948e+11Hz -0.0120403 0.00206872
+ 2.949e+11Hz -0.0120119 0.00204249
+ 2.95e+11Hz -0.0119839 0.00201619
+ 2.951e+11Hz -0.0119562 0.00198983
+ 2.952e+11Hz -0.0119289 0.0019634
+ 2.953e+11Hz -0.0119019 0.00193693
+ 2.954e+11Hz -0.0118753 0.00191041
+ 2.955e+11Hz -0.011849 0.00188385
+ 2.956e+11Hz -0.0118231 0.00185725
+ 2.957e+11Hz -0.0117975 0.00183063
+ 2.958e+11Hz -0.0117722 0.00180398
+ 2.959e+11Hz -0.0117473 0.00177732
+ 2.96e+11Hz -0.0117228 0.00175065
+ 2.961e+11Hz -0.0116985 0.00172397
+ 2.962e+11Hz -0.0116746 0.0016973
+ 2.963e+11Hz -0.011651 0.00167063
+ 2.964e+11Hz -0.0116278 0.00164396
+ 2.965e+11Hz -0.0116048 0.00161732
+ 2.966e+11Hz -0.0115822 0.00159069
+ 2.967e+11Hz -0.0115599 0.00156409
+ 2.968e+11Hz -0.0115379 0.00153752
+ 2.969e+11Hz -0.0115163 0.00151099
+ 2.97e+11Hz -0.0114949 0.0014845
+ 2.971e+11Hz -0.0114738 0.00145805
+ 2.972e+11Hz -0.0114531 0.00143165
+ 2.973e+11Hz -0.0114326 0.0014053
+ 2.974e+11Hz -0.0114124 0.00137901
+ 2.975e+11Hz -0.0113926 0.00135278
+ 2.976e+11Hz -0.011373 0.00132662
+ 2.977e+11Hz -0.0113537 0.00130052
+ 2.978e+11Hz -0.0113347 0.0012745
+ 2.979e+11Hz -0.0113159 0.00124856
+ 2.98e+11Hz -0.0112974 0.00122269
+ 2.981e+11Hz -0.0112792 0.00119691
+ 2.982e+11Hz -0.0112613 0.00117122
+ 2.983e+11Hz -0.0112436 0.00114562
+ 2.984e+11Hz -0.0112262 0.00112011
+ 2.985e+11Hz -0.011209 0.0010947
+ 2.986e+11Hz -0.0111921 0.00106938
+ 2.987e+11Hz -0.0111754 0.00104417
+ 2.988e+11Hz -0.011159 0.00101906
+ 2.989e+11Hz -0.0111428 0.000994064
+ 2.99e+11Hz -0.0111268 0.000969174
+ 2.991e+11Hz -0.0111111 0.000944394
+ 2.992e+11Hz -0.0110956 0.000919729
+ 2.993e+11Hz -0.0110803 0.000895179
+ 2.994e+11Hz -0.0110652 0.000870747
+ 2.995e+11Hz -0.0110503 0.000846435
+ 2.996e+11Hz -0.0110357 0.000822244
+ 2.997e+11Hz -0.0110212 0.000798175
+ 2.998e+11Hz -0.0110069 0.000774231
+ 2.999e+11Hz -0.0109929 0.000750413
+ 3e+11Hz -0.010979 0.000726721
+ ]

.ENDS
.SUBCKT Sub_SPfile_X6 1 2 3
R1N 1 10 -50
R1P 10 11 100
R2N 2 20 -50
R2P 20 21 100

A11 %vd(10 3) %vd(11, 12) xfer1
.model xfer1 xfer R_I=true table=[
+ 0Hz 0.00819703 0
+ 1e+08Hz 0.00819728 3.05641e-05
+ 2e+08Hz 0.00819804 6.11124e-05
+ 3e+08Hz 0.00819932 9.16293e-05
+ 4e+08Hz 0.0082011 0.000122099
+ 5e+08Hz 0.00820338 0.000152506
+ 6e+08Hz 0.00820617 0.000182835
+ 7e+08Hz 0.00820946 0.00021307
+ 8e+08Hz 0.00821325 0.000243195
+ 9e+08Hz 0.00821754 0.000273195
+ 1e+09Hz 0.00822232 0.000303056
+ 1.1e+09Hz 0.00822759 0.00033276
+ 1.2e+09Hz 0.00823335 0.000362295
+ 1.3e+09Hz 0.00823959 0.000391643
+ 1.4e+09Hz 0.0082463 0.000420792
+ 1.5e+09Hz 0.00825348 0.000449724
+ 1.6e+09Hz 0.00826113 0.000478427
+ 1.7e+09Hz 0.00826924 0.000506886
+ 1.8e+09Hz 0.00827781 0.000535086
+ 1.9e+09Hz 0.00828682 0.000563013
+ 2e+09Hz 0.00829627 0.000590653
+ 2.1e+09Hz 0.00830615 0.000617993
+ 2.2e+09Hz 0.00831646 0.000645019
+ 2.3e+09Hz 0.00832718 0.000671717
+ 2.4e+09Hz 0.00833831 0.000698074
+ 2.5e+09Hz 0.00834984 0.000724078
+ 2.6e+09Hz 0.00836177 0.000749716
+ 2.7e+09Hz 0.00837407 0.000774974
+ 2.8e+09Hz 0.00838675 0.000799842
+ 2.9e+09Hz 0.00839979 0.000824307
+ 3e+09Hz 0.00841318 0.000848358
+ 3.1e+09Hz 0.00842692 0.000871982
+ 3.2e+09Hz 0.00844098 0.000895169
+ 3.3e+09Hz 0.00845537 0.000917909
+ 3.4e+09Hz 0.00847007 0.000940189
+ 3.5e+09Hz 0.00848506 0.000962001
+ 3.6e+09Hz 0.00850034 0.000983333
+ 3.7e+09Hz 0.0085159 0.00100418
+ 3.8e+09Hz 0.00853172 0.00102452
+ 3.9e+09Hz 0.00854779 0.00104436
+ 4e+09Hz 0.0085641 0.00106368
+ 4.1e+09Hz 0.00858063 0.00108248
+ 4.2e+09Hz 0.00859738 0.00110075
+ 4.3e+09Hz 0.00861432 0.00111847
+ 4.4e+09Hz 0.00863146 0.00113565
+ 4.5e+09Hz 0.00864876 0.00115228
+ 4.6e+09Hz 0.00866623 0.00116834
+ 4.7e+09Hz 0.00868384 0.00118383
+ 4.8e+09Hz 0.00870158 0.00119875
+ 4.9e+09Hz 0.00871945 0.00121309
+ 5e+09Hz 0.00873742 0.00122685
+ 5.1e+09Hz 0.00875548 0.00124001
+ 5.2e+09Hz 0.00877361 0.00125258
+ 5.3e+09Hz 0.00879181 0.00126455
+ 5.4e+09Hz 0.00881006 0.00127592
+ 5.5e+09Hz 0.00882833 0.00128667
+ 5.6e+09Hz 0.00884664 0.00129682
+ 5.7e+09Hz 0.00886494 0.00130636
+ 5.8e+09Hz 0.00888324 0.00131528
+ 5.9e+09Hz 0.00890151 0.00132358
+ 6e+09Hz 0.00891974 0.00133126
+ 6.1e+09Hz 0.00893792 0.00133832
+ 6.2e+09Hz 0.00895604 0.00134476
+ 6.3e+09Hz 0.00897407 0.00135057
+ 6.4e+09Hz 0.00899201 0.00135576
+ 6.5e+09Hz 0.00900983 0.00136033
+ 6.6e+09Hz 0.00902754 0.00136427
+ 6.7e+09Hz 0.0090451 0.00136759
+ 6.8e+09Hz 0.00906251 0.00137028
+ 6.9e+09Hz 0.00907975 0.00137236
+ 7e+09Hz 0.00909681 0.00137381
+ 7.1e+09Hz 0.00911367 0.00137465
+ 7.2e+09Hz 0.00913032 0.00137486
+ 7.3e+09Hz 0.00914676 0.00137447
+ 7.4e+09Hz 0.00916295 0.00137346
+ 7.5e+09Hz 0.00917889 0.00137185
+ 7.6e+09Hz 0.00919457 0.00136963
+ 7.7e+09Hz 0.00920997 0.00136681
+ 7.8e+09Hz 0.00922507 0.0013634
+ 7.9e+09Hz 0.00923988 0.00135939
+ 8e+09Hz 0.00925436 0.0013548
+ 8.1e+09Hz 0.00926852 0.00134962
+ 8.2e+09Hz 0.00928233 0.00134386
+ 8.3e+09Hz 0.00929579 0.00133753
+ 8.4e+09Hz 0.00930887 0.00133064
+ 8.5e+09Hz 0.00932158 0.00132318
+ 8.6e+09Hz 0.0093339 0.00131517
+ 8.7e+09Hz 0.00934581 0.00130661
+ 8.8e+09Hz 0.0093573 0.00129751
+ 8.9e+09Hz 0.00936837 0.00128787
+ 9e+09Hz 0.009379 0.00127771
+ 9.1e+09Hz 0.00938918 0.00126703
+ 9.2e+09Hz 0.0093989 0.00125583
+ 9.3e+09Hz 0.00940815 0.00124413
+ 9.4e+09Hz 0.00941692 0.00123193
+ 9.5e+09Hz 0.00942519 0.00121925
+ 9.6e+09Hz 0.00943297 0.00120608
+ 9.7e+09Hz 0.00944023 0.00119244
+ 9.8e+09Hz 0.00944697 0.00117834
+ 9.9e+09Hz 0.00945318 0.00116378
+ 1e+10Hz 0.00945885 0.00114878
+ 1.01e+10Hz 0.00946397 0.00113334
+ 1.02e+10Hz 0.00946854 0.00111748
+ 1.03e+10Hz 0.00947254 0.0011012
+ 1.04e+10Hz 0.00947597 0.00108451
+ 1.05e+10Hz 0.00947881 0.00106743
+ 1.06e+10Hz 0.00948107 0.00104995
+ 1.07e+10Hz 0.00948273 0.0010321
+ 1.08e+10Hz 0.00948379 0.00101389
+ 1.09e+10Hz 0.00948424 0.000995314
+ 1.1e+10Hz 0.00948407 0.000976393
+ 1.11e+10Hz 0.00948327 0.000957136
+ 1.12e+10Hz 0.00948185 0.000937553
+ 1.13e+10Hz 0.00947979 0.000917656
+ 1.14e+10Hz 0.00947709 0.000897454
+ 1.15e+10Hz 0.00947375 0.000876959
+ 1.16e+10Hz 0.00946975 0.00085618
+ 1.17e+10Hz 0.0094651 0.00083513
+ 1.18e+10Hz 0.00945979 0.00081382
+ 1.19e+10Hz 0.00945381 0.000792259
+ 1.2e+10Hz 0.00944716 0.000770459
+ 1.21e+10Hz 0.00943984 0.000748432
+ 1.22e+10Hz 0.00943184 0.000726188
+ 1.23e+10Hz 0.00942317 0.000703738
+ 1.24e+10Hz 0.00941381 0.000681093
+ 1.25e+10Hz 0.00940376 0.000658265
+ 1.26e+10Hz 0.00939302 0.000635264
+ 1.27e+10Hz 0.0093816 0.000612102
+ 1.28e+10Hz 0.00936948 0.000588789
+ 1.29e+10Hz 0.00935666 0.000565337
+ 1.3e+10Hz 0.00934315 0.000541757
+ 1.31e+10Hz 0.00932894 0.00051806
+ 1.32e+10Hz 0.00931403 0.000494256
+ 1.33e+10Hz 0.00929842 0.000470357
+ 1.34e+10Hz 0.0092821 0.000446374
+ 1.35e+10Hz 0.00926509 0.000422317
+ 1.36e+10Hz 0.00924737 0.000398197
+ 1.37e+10Hz 0.00922895 0.000374025
+ 1.38e+10Hz 0.00920983 0.000349812
+ 1.39e+10Hz 0.00919001 0.000325568
+ 1.4e+10Hz 0.00916949 0.000301304
+ 1.41e+10Hz 0.00914826 0.000277029
+ 1.42e+10Hz 0.00912634 0.000252756
+ 1.43e+10Hz 0.00910371 0.000228493
+ 1.44e+10Hz 0.00908039 0.000204251
+ 1.45e+10Hz 0.00905638 0.00018004
+ 1.46e+10Hz 0.00903167 0.000155871
+ 1.47e+10Hz 0.00900627 0.000131753
+ 1.48e+10Hz 0.00898017 0.000107695
+ 1.49e+10Hz 0.00895339 8.37089e-05
+ 1.5e+10Hz 0.00892593 5.98025e-05
+ 1.51e+10Hz 0.00889778 3.59859e-05
+ 1.52e+10Hz 0.00886895 1.22685e-05
+ 1.53e+10Hz 0.00883945 -1.13405e-05
+ 1.54e+10Hz 0.00880927 -3.4832e-05
+ 1.55e+10Hz 0.00877842 -5.81968e-05
+ 1.56e+10Hz 0.00874691 -8.14261e-05
+ 1.57e+10Hz 0.00871473 -0.000104511
+ 1.58e+10Hz 0.00868189 -0.000127443
+ 1.59e+10Hz 0.00864839 -0.000150214
+ 1.6e+10Hz 0.00861424 -0.000172815
+ 1.61e+10Hz 0.00857944 -0.000195238
+ 1.62e+10Hz 0.008544 -0.000217475
+ 1.63e+10Hz 0.00850792 -0.000239517
+ 1.64e+10Hz 0.0084712 -0.000261358
+ 1.65e+10Hz 0.00843386 -0.000282989
+ 1.66e+10Hz 0.00839588 -0.000304403
+ 1.67e+10Hz 0.00835729 -0.000325593
+ 1.68e+10Hz 0.00831808 -0.000346551
+ 1.69e+10Hz 0.00827826 -0.000367269
+ 1.7e+10Hz 0.00823783 -0.000387743
+ 1.71e+10Hz 0.0081968 -0.000407963
+ 1.72e+10Hz 0.00815517 -0.000427924
+ 1.73e+10Hz 0.00811296 -0.00044762
+ 1.74e+10Hz 0.00807016 -0.000467044
+ 1.75e+10Hz 0.00802677 -0.000486189
+ 1.76e+10Hz 0.00798282 -0.00050505
+ 1.77e+10Hz 0.00793829 -0.00052362
+ 1.78e+10Hz 0.00789321 -0.000541895
+ 1.79e+10Hz 0.00784756 -0.000559869
+ 1.8e+10Hz 0.00780136 -0.000577535
+ 1.81e+10Hz 0.00775462 -0.00059489
+ 1.82e+10Hz 0.00770734 -0.000611927
+ 1.83e+10Hz 0.00765952 -0.000628641
+ 1.84e+10Hz 0.00761118 -0.000645029
+ 1.85e+10Hz 0.00756231 -0.000661085
+ 1.86e+10Hz 0.00751293 -0.000676805
+ 1.87e+10Hz 0.00746304 -0.000692184
+ 1.88e+10Hz 0.00741264 -0.000707218
+ 1.89e+10Hz 0.00736175 -0.000721903
+ 1.9e+10Hz 0.00731036 -0.000736236
+ 1.91e+10Hz 0.00725849 -0.000750212
+ 1.92e+10Hz 0.00720614 -0.000763828
+ 1.93e+10Hz 0.00715331 -0.00077708
+ 1.94e+10Hz 0.00710002 -0.000789965
+ 1.95e+10Hz 0.00704627 -0.00080248
+ 1.96e+10Hz 0.00699206 -0.000814622
+ 1.97e+10Hz 0.0069374 -0.000826387
+ 1.98e+10Hz 0.0068823 -0.000837774
+ 1.99e+10Hz 0.00682676 -0.000848779
+ 2e+10Hz 0.00677079 -0.0008594
+ 2.01e+10Hz 0.00671439 -0.000869634
+ 2.02e+10Hz 0.00665758 -0.00087948
+ 2.03e+10Hz 0.00660035 -0.000888935
+ 2.04e+10Hz 0.00654272 -0.000897997
+ 2.05e+10Hz 0.00648469 -0.000906665
+ 2.06e+10Hz 0.00642626 -0.000914936
+ 2.07e+10Hz 0.00636744 -0.000922809
+ 2.08e+10Hz 0.00630824 -0.000930284
+ 2.09e+10Hz 0.00624866 -0.000937357
+ 2.1e+10Hz 0.00618871 -0.000944028
+ 2.11e+10Hz 0.00612839 -0.000950296
+ 2.12e+10Hz 0.00606771 -0.00095616
+ 2.13e+10Hz 0.00600668 -0.000961618
+ 2.14e+10Hz 0.00594529 -0.000966671
+ 2.15e+10Hz 0.00588356 -0.000971318
+ 2.16e+10Hz 0.0058215 -0.000975556
+ 2.17e+10Hz 0.0057591 -0.000979388
+ 2.18e+10Hz 0.00569637 -0.000982811
+ 2.19e+10Hz 0.00563332 -0.000985826
+ 2.2e+10Hz 0.00556995 -0.000988433
+ 2.21e+10Hz 0.00550627 -0.00099063
+ 2.22e+10Hz 0.00544229 -0.00099242
+ 2.23e+10Hz 0.005378 -0.0009938
+ 2.24e+10Hz 0.00531341 -0.000994772
+ 2.25e+10Hz 0.00524853 -0.000995336
+ 2.26e+10Hz 0.00518336 -0.000995492
+ 2.27e+10Hz 0.00511791 -0.00099524
+ 2.28e+10Hz 0.00505219 -0.000994581
+ 2.29e+10Hz 0.00498618 -0.000993516
+ 2.3e+10Hz 0.00491991 -0.000992045
+ 2.31e+10Hz 0.00485337 -0.000990169
+ 2.32e+10Hz 0.00478658 -0.000987888
+ 2.33e+10Hz 0.00471952 -0.000985204
+ 2.34e+10Hz 0.00465222 -0.000982117
+ 2.35e+10Hz 0.00458466 -0.000978628
+ 2.36e+10Hz 0.00451686 -0.000974738
+ 2.37e+10Hz 0.00444882 -0.000970448
+ 2.38e+10Hz 0.00438055 -0.000965759
+ 2.39e+10Hz 0.00431204 -0.000960673
+ 2.4e+10Hz 0.0042433 -0.00095519
+ 2.41e+10Hz 0.00417434 -0.000949312
+ 2.42e+10Hz 0.00410516 -0.00094304
+ 2.43e+10Hz 0.00403576 -0.000936376
+ 2.44e+10Hz 0.00396614 -0.00092932
+ 2.45e+10Hz 0.00389631 -0.000921874
+ 2.46e+10Hz 0.00382627 -0.000914039
+ 2.47e+10Hz 0.00375603 -0.000905817
+ 2.48e+10Hz 0.00368559 -0.00089721
+ 2.49e+10Hz 0.00361494 -0.000888218
+ 2.5e+10Hz 0.0035441 -0.000878843
+ 2.51e+10Hz 0.00347307 -0.000869088
+ 2.52e+10Hz 0.00340185 -0.000858952
+ 2.53e+10Hz 0.00333043 -0.000848439
+ 2.54e+10Hz 0.00325883 -0.000837548
+ 2.55e+10Hz 0.00318705 -0.000826283
+ 2.56e+10Hz 0.00311509 -0.000814645
+ 2.57e+10Hz 0.00304295 -0.000802635
+ 2.58e+10Hz 0.00297063 -0.000790254
+ 2.59e+10Hz 0.00289814 -0.000777505
+ 2.6e+10Hz 0.00282547 -0.000764389
+ 2.61e+10Hz 0.00275264 -0.000750907
+ 2.62e+10Hz 0.00267964 -0.000737062
+ 2.63e+10Hz 0.00260647 -0.000722855
+ 2.64e+10Hz 0.00253314 -0.000708286
+ 2.65e+10Hz 0.00245964 -0.000693359
+ 2.66e+10Hz 0.00238598 -0.000678075
+ 2.67e+10Hz 0.00231217 -0.000662434
+ 2.68e+10Hz 0.0022382 -0.000646439
+ 2.69e+10Hz 0.00216407 -0.000630091
+ 2.7e+10Hz 0.00208978 -0.000613392
+ 2.71e+10Hz 0.00201534 -0.000596344
+ 2.72e+10Hz 0.00194075 -0.000578946
+ 2.73e+10Hz 0.00186601 -0.000561202
+ 2.74e+10Hz 0.00179112 -0.000543113
+ 2.75e+10Hz 0.00171607 -0.00052468
+ 2.76e+10Hz 0.00164088 -0.000505904
+ 2.77e+10Hz 0.00156555 -0.000486786
+ 2.78e+10Hz 0.00149006 -0.000467329
+ 2.79e+10Hz 0.00141443 -0.000447533
+ 2.8e+10Hz 0.00133866 -0.0004274
+ 2.81e+10Hz 0.00126274 -0.000406931
+ 2.82e+10Hz 0.00118668 -0.000386126
+ 2.83e+10Hz 0.00111048 -0.000364989
+ 2.84e+10Hz 0.00103414 -0.000343518
+ 2.85e+10Hz 0.00095765 -0.000321716
+ 2.86e+10Hz 0.000881023 -0.000299584
+ 2.87e+10Hz 0.000804256 -0.000277122
+ 2.88e+10Hz 0.000727349 -0.000254332
+ 2.89e+10Hz 0.000650302 -0.000231215
+ 2.9e+10Hz 0.000573115 -0.000207771
+ 2.91e+10Hz 0.00049579 -0.000184002
+ 2.92e+10Hz 0.000418326 -0.000159908
+ 2.93e+10Hz 0.000340723 -0.00013549
+ 2.94e+10Hz 0.000262982 -0.000110749
+ 2.95e+10Hz 0.000185103 -8.56851e-05
+ 2.96e+10Hz 0.000107086 -6.02998e-05
+ 2.97e+10Hz 2.89309e-05 -3.45934e-05
+ 2.98e+10Hz -4.93622e-05 -8.56649e-06
+ 2.99e+10Hz -0.000127793 1.77804e-05
+ 3e+10Hz -0.000206362 4.44468e-05
+ 3.01e+10Hz -0.000285069 7.14322e-05
+ 3.02e+10Hz -0.000363913 9.87362e-05
+ 3.03e+10Hz -0.000442896 0.000126359
+ 3.04e+10Hz -0.000522016 0.000154299
+ 3.05e+10Hz -0.000601275 0.000182556
+ 3.06e+10Hz -0.000680671 0.000211131
+ 3.07e+10Hz -0.000760206 0.000240024
+ 3.08e+10Hz -0.00083988 0.000269233
+ 3.09e+10Hz -0.000919691 0.00029876
+ 3.1e+10Hz -0.000999642 0.000328603
+ 3.11e+10Hz -0.00107973 0.000358763
+ 3.12e+10Hz -0.00115996 0.00038924
+ 3.13e+10Hz -0.00124033 0.000420035
+ 3.14e+10Hz -0.00132084 0.000451146
+ 3.15e+10Hz -0.00140148 0.000482574
+ 3.16e+10Hz -0.00148227 0.000514321
+ 3.17e+10Hz -0.00156319 0.000546384
+ 3.18e+10Hz -0.00164426 0.000578766
+ 3.19e+10Hz -0.00172547 0.000611467
+ 3.2e+10Hz -0.00180681 0.000644486
+ 3.21e+10Hz -0.0018883 0.000677825
+ 3.22e+10Hz -0.00196993 0.000711483
+ 3.23e+10Hz -0.0020517 0.000745461
+ 3.24e+10Hz -0.00213361 0.00077976
+ 3.25e+10Hz -0.00221566 0.000814381
+ 3.26e+10Hz -0.00229785 0.000849324
+ 3.27e+10Hz -0.00238019 0.000884589
+ 3.28e+10Hz -0.00246266 0.000920178
+ 3.29e+10Hz -0.00254528 0.00095609
+ 3.3e+10Hz -0.00262804 0.000992328
+ 3.31e+10Hz -0.00271094 0.00102889
+ 3.32e+10Hz -0.00279399 0.00106578
+ 3.33e+10Hz -0.00287717 0.001103
+ 3.34e+10Hz -0.0029605 0.00114055
+ 3.35e+10Hz -0.00304397 0.00117842
+ 3.36e+10Hz -0.00312758 0.00121663
+ 3.37e+10Hz -0.00321133 0.00125517
+ 3.38e+10Hz -0.00329523 0.00129404
+ 3.39e+10Hz -0.00337926 0.00133324
+ 3.4e+10Hz -0.00346344 0.00137278
+ 3.41e+10Hz -0.00354776 0.00141265
+ 3.42e+10Hz -0.00363222 0.00145286
+ 3.43e+10Hz -0.00371682 0.00149341
+ 3.44e+10Hz -0.00380156 0.0015343
+ 3.45e+10Hz -0.00388645 0.00157553
+ 3.46e+10Hz -0.00397147 0.00161711
+ 3.47e+10Hz -0.00405664 0.00165902
+ 3.48e+10Hz -0.00414194 0.00170128
+ 3.49e+10Hz -0.00422738 0.00174389
+ 3.5e+10Hz -0.00431296 0.00178684
+ 3.51e+10Hz -0.00439869 0.00183015
+ 3.52e+10Hz -0.00448454 0.0018738
+ 3.53e+10Hz -0.00457054 0.00191781
+ 3.54e+10Hz -0.00465667 0.00196216
+ 3.55e+10Hz -0.00474294 0.00200688
+ 3.56e+10Hz -0.00482935 0.00205195
+ 3.57e+10Hz -0.00491589 0.00209737
+ 3.58e+10Hz -0.00500257 0.00214316
+ 3.59e+10Hz -0.00508938 0.00218931
+ 3.6e+10Hz -0.00517632 0.00223582
+ 3.61e+10Hz -0.0052634 0.00228269
+ 3.62e+10Hz -0.00535061 0.00232993
+ 3.63e+10Hz -0.00543795 0.00237754
+ 3.64e+10Hz -0.00552542 0.00242551
+ 3.65e+10Hz -0.00561302 0.00247386
+ 3.66e+10Hz -0.00570074 0.00252257
+ 3.67e+10Hz -0.0057886 0.00257166
+ 3.68e+10Hz -0.00587658 0.00262113
+ 3.69e+10Hz -0.00596469 0.00267097
+ 3.7e+10Hz -0.00605292 0.00272119
+ 3.71e+10Hz -0.00614128 0.00277179
+ 3.72e+10Hz -0.00622975 0.00282277
+ 3.73e+10Hz -0.00631835 0.00287414
+ 3.74e+10Hz -0.00640707 0.00292589
+ 3.75e+10Hz -0.00649591 0.00297802
+ 3.76e+10Hz -0.00658486 0.00303054
+ 3.77e+10Hz -0.00667393 0.00308346
+ 3.78e+10Hz -0.00676312 0.00313676
+ 3.79e+10Hz -0.00685242 0.00319046
+ 3.8e+10Hz -0.00694183 0.00324455
+ 3.81e+10Hz -0.00703135 0.00329904
+ 3.82e+10Hz -0.00712098 0.00335393
+ 3.83e+10Hz -0.00721072 0.00340921
+ 3.84e+10Hz -0.00730056 0.0034649
+ 3.85e+10Hz -0.00739051 0.00352098
+ 3.86e+10Hz -0.00748056 0.00357748
+ 3.87e+10Hz -0.00757072 0.00363437
+ 3.88e+10Hz -0.00766097 0.00369168
+ 3.89e+10Hz -0.00775132 0.00374939
+ 3.9e+10Hz -0.00784177 0.00380751
+ 3.91e+10Hz -0.00793231 0.00386604
+ 3.92e+10Hz -0.00802295 0.00392499
+ 3.93e+10Hz -0.00811367 0.00398435
+ 3.94e+10Hz -0.00820449 0.00404412
+ 3.95e+10Hz -0.00829539 0.00410431
+ 3.96e+10Hz -0.00838638 0.00416492
+ 3.97e+10Hz -0.00847745 0.00422596
+ 3.98e+10Hz -0.0085686 0.00428741
+ 3.99e+10Hz -0.00865983 0.00434928
+ 4e+10Hz -0.00875114 0.00441158
+ 4.01e+10Hz -0.00884253 0.0044743
+ 4.02e+10Hz -0.00893399 0.00453745
+ 4.03e+10Hz -0.00902552 0.00460103
+ 4.04e+10Hz -0.00911712 0.00466503
+ 4.05e+10Hz -0.00920878 0.00472947
+ 4.06e+10Hz -0.00930052 0.00479434
+ 4.07e+10Hz -0.00939231 0.00485964
+ 4.08e+10Hz -0.00948417 0.00492537
+ 4.09e+10Hz -0.00957608 0.00499154
+ 4.1e+10Hz -0.00966805 0.00505814
+ 4.11e+10Hz -0.00976007 0.00512518
+ 4.12e+10Hz -0.00985215 0.00519266
+ 4.13e+10Hz -0.00994428 0.00526057
+ 4.14e+10Hz -0.0100365 0.00532893
+ 4.15e+10Hz -0.0101287 0.00539772
+ 4.16e+10Hz -0.0102209 0.00546696
+ 4.17e+10Hz -0.0103132 0.00553664
+ 4.18e+10Hz -0.0104056 0.00560676
+ 4.19e+10Hz -0.0104979 0.00567733
+ 4.2e+10Hz -0.0105904 0.00574834
+ 4.21e+10Hz -0.0106828 0.0058198
+ 4.22e+10Hz -0.0107753 0.00589171
+ 4.23e+10Hz -0.0108677 0.00596406
+ 4.24e+10Hz -0.0109603 0.00603686
+ 4.25e+10Hz -0.0110528 0.0061101
+ 4.26e+10Hz -0.0111454 0.0061838
+ 4.27e+10Hz -0.0112379 0.00625795
+ 4.28e+10Hz -0.0113305 0.00633254
+ 4.29e+10Hz -0.0114231 0.00640759
+ 4.3e+10Hz -0.0115157 0.00648309
+ 4.31e+10Hz -0.0116083 0.00655904
+ 4.32e+10Hz -0.0117009 0.00663544
+ 4.33e+10Hz -0.0117935 0.0067123
+ 4.34e+10Hz -0.0118862 0.0067896
+ 4.35e+10Hz -0.0119788 0.00686737
+ 4.36e+10Hz -0.0120714 0.00694558
+ 4.37e+10Hz -0.012164 0.00702425
+ 4.38e+10Hz -0.0122566 0.00710337
+ 4.39e+10Hz -0.0123491 0.00718295
+ 4.4e+10Hz -0.0124417 0.00726298
+ 4.41e+10Hz -0.0125342 0.00734347
+ 4.42e+10Hz -0.0126267 0.00742441
+ 4.43e+10Hz -0.0127192 0.00750581
+ 4.44e+10Hz -0.0128117 0.00758767
+ 4.45e+10Hz -0.0129041 0.00766997
+ 4.46e+10Hz -0.0129965 0.00775274
+ 4.47e+10Hz -0.0130889 0.00783596
+ 4.48e+10Hz -0.0131813 0.00791963
+ 4.49e+10Hz -0.0132735 0.00800376
+ 4.5e+10Hz -0.0133658 0.00808835
+ 4.51e+10Hz -0.013458 0.00817339
+ 4.52e+10Hz -0.0135502 0.00825888
+ 4.53e+10Hz -0.0136423 0.00834483
+ 4.54e+10Hz -0.0137344 0.00843124
+ 4.55e+10Hz -0.0138264 0.0085181
+ 4.56e+10Hz -0.0139183 0.00860541
+ 4.57e+10Hz -0.0140102 0.00869318
+ 4.58e+10Hz -0.0141021 0.0087814
+ 4.59e+10Hz -0.0141938 0.00887007
+ 4.6e+10Hz -0.0142856 0.0089592
+ 4.61e+10Hz -0.0143772 0.00904878
+ 4.62e+10Hz -0.0144688 0.00913881
+ 4.63e+10Hz -0.0145603 0.0092293
+ 4.64e+10Hz -0.0146517 0.00932024
+ 4.65e+10Hz -0.0147431 0.00941162
+ 4.66e+10Hz -0.0148343 0.00950346
+ 4.67e+10Hz -0.0149255 0.00959575
+ 4.68e+10Hz -0.0150166 0.00968849
+ 4.69e+10Hz -0.0151076 0.00978168
+ 4.7e+10Hz -0.0151986 0.00987531
+ 4.71e+10Hz -0.0152894 0.0099694
+ 4.72e+10Hz -0.0153801 0.0100639
+ 4.73e+10Hz -0.0154708 0.0101589
+ 4.74e+10Hz -0.0155613 0.0102543
+ 4.75e+10Hz -0.0156518 0.0103502
+ 4.76e+10Hz -0.0157422 0.0104465
+ 4.77e+10Hz -0.0158324 0.0105433
+ 4.78e+10Hz -0.0159226 0.0106405
+ 4.79e+10Hz -0.0160126 0.0107381
+ 4.8e+10Hz -0.0161025 0.0108362
+ 4.81e+10Hz -0.0161923 0.0109347
+ 4.82e+10Hz -0.016282 0.0110337
+ 4.83e+10Hz -0.0163716 0.0111331
+ 4.84e+10Hz -0.0164611 0.011233
+ 4.85e+10Hz -0.0165504 0.0113333
+ 4.86e+10Hz -0.0166397 0.011434
+ 4.87e+10Hz -0.0167288 0.0115351
+ 4.88e+10Hz -0.0168177 0.0116367
+ 4.89e+10Hz -0.0169066 0.0117388
+ 4.9e+10Hz -0.0169953 0.0118412
+ 4.91e+10Hz -0.0170839 0.0119442
+ 4.92e+10Hz -0.0171723 0.0120475
+ 4.93e+10Hz -0.0172607 0.0121513
+ 4.94e+10Hz -0.0173489 0.0122554
+ 4.95e+10Hz -0.0174369 0.0123601
+ 4.96e+10Hz -0.0175248 0.0124651
+ 4.97e+10Hz -0.0176126 0.0125706
+ 4.98e+10Hz -0.0177002 0.0126765
+ 4.99e+10Hz -0.0177877 0.0127829
+ 5e+10Hz -0.017875 0.0128896
+ 5.01e+10Hz -0.0179622 0.0129968
+ 5.02e+10Hz -0.0180492 0.0131044
+ 5.03e+10Hz -0.0181361 0.0132125
+ 5.04e+10Hz -0.0182228 0.0133209
+ 5.05e+10Hz -0.0183093 0.0134298
+ 5.06e+10Hz -0.0183958 0.0135391
+ 5.07e+10Hz -0.018482 0.0136488
+ 5.08e+10Hz -0.0185681 0.013759
+ 5.09e+10Hz -0.018654 0.0138695
+ 5.1e+10Hz -0.0187398 0.0139805
+ 5.11e+10Hz -0.0188254 0.0140919
+ 5.12e+10Hz -0.0189108 0.0142037
+ 5.13e+10Hz -0.0189961 0.0143159
+ 5.14e+10Hz -0.0190812 0.0144285
+ 5.15e+10Hz -0.0191661 0.0145416
+ 5.16e+10Hz -0.0192509 0.014655
+ 5.17e+10Hz -0.0193355 0.0147689
+ 5.18e+10Hz -0.0194199 0.0148831
+ 5.19e+10Hz -0.0195041 0.0149978
+ 5.2e+10Hz -0.0195881 0.0151129
+ 5.21e+10Hz -0.019672 0.0152284
+ 5.22e+10Hz -0.0197557 0.0153443
+ 5.23e+10Hz -0.0198392 0.0154606
+ 5.24e+10Hz -0.0199226 0.0155773
+ 5.25e+10Hz -0.0200057 0.0156944
+ 5.26e+10Hz -0.0200887 0.0158119
+ 5.27e+10Hz -0.0201715 0.0159298
+ 5.28e+10Hz -0.020254 0.0160481
+ 5.29e+10Hz -0.0203364 0.0161668
+ 5.3e+10Hz -0.0204187 0.016286
+ 5.31e+10Hz -0.0205007 0.0164055
+ 5.32e+10Hz -0.0205825 0.0165254
+ 5.33e+10Hz -0.0206641 0.0166457
+ 5.34e+10Hz -0.0207456 0.0167664
+ 5.35e+10Hz -0.0208268 0.0168874
+ 5.36e+10Hz -0.0209079 0.0170089
+ 5.37e+10Hz -0.0209887 0.0171308
+ 5.38e+10Hz -0.0210694 0.0172531
+ 5.39e+10Hz -0.0211498 0.0173757
+ 5.4e+10Hz -0.0212301 0.0174988
+ 5.41e+10Hz -0.0213101 0.0176222
+ 5.42e+10Hz -0.02139 0.0177461
+ 5.43e+10Hz -0.0214696 0.0178703
+ 5.44e+10Hz -0.021549 0.0179949
+ 5.45e+10Hz -0.0216283 0.0181199
+ 5.46e+10Hz -0.0217073 0.0182453
+ 5.47e+10Hz -0.0217861 0.018371
+ 5.48e+10Hz -0.0218647 0.0184972
+ 5.49e+10Hz -0.0219431 0.0186237
+ 5.5e+10Hz -0.0220212 0.0187506
+ 5.51e+10Hz -0.0220992 0.0188779
+ 5.52e+10Hz -0.022177 0.0190056
+ 5.53e+10Hz -0.0222545 0.0191337
+ 5.54e+10Hz -0.0223318 0.0192621
+ 5.55e+10Hz -0.0224089 0.019391
+ 5.56e+10Hz -0.0224858 0.0195202
+ 5.57e+10Hz -0.0225624 0.0196498
+ 5.58e+10Hz -0.0226389 0.0197797
+ 5.59e+10Hz -0.0227151 0.0199101
+ 5.6e+10Hz -0.0227911 0.0200408
+ 5.61e+10Hz -0.0228669 0.0201719
+ 5.62e+10Hz -0.0229424 0.0203034
+ 5.63e+10Hz -0.0230178 0.0204352
+ 5.64e+10Hz -0.0230928 0.0205674
+ 5.65e+10Hz -0.0231677 0.0207
+ 5.66e+10Hz -0.0232423 0.020833
+ 5.67e+10Hz -0.0233168 0.0209664
+ 5.68e+10Hz -0.0233909 0.0211001
+ 5.69e+10Hz -0.0234649 0.0212342
+ 5.7e+10Hz -0.0235386 0.0213686
+ 5.71e+10Hz -0.0236121 0.0215035
+ 5.72e+10Hz -0.0236853 0.0216387
+ 5.73e+10Hz -0.0237584 0.0217743
+ 5.74e+10Hz -0.0238311 0.0219102
+ 5.75e+10Hz -0.0239037 0.0220465
+ 5.76e+10Hz -0.0239759 0.0221832
+ 5.77e+10Hz -0.024048 0.0223203
+ 5.78e+10Hz -0.0241198 0.0224577
+ 5.79e+10Hz -0.0241914 0.0225955
+ 5.8e+10Hz -0.0242627 0.0227337
+ 5.81e+10Hz -0.0243338 0.0228722
+ 5.82e+10Hz -0.0244046 0.0230111
+ 5.83e+10Hz -0.0244753 0.0231504
+ 5.84e+10Hz -0.0245456 0.02329
+ 5.85e+10Hz -0.0246157 0.02343
+ 5.86e+10Hz -0.0246855 0.0235704
+ 5.87e+10Hz -0.0247551 0.0237111
+ 5.88e+10Hz -0.0248245 0.0238522
+ 5.89e+10Hz -0.0248936 0.0239937
+ 5.9e+10Hz -0.0249624 0.0241355
+ 5.91e+10Hz -0.025031 0.0242777
+ 5.92e+10Hz -0.0250993 0.0244203
+ 5.93e+10Hz -0.0251674 0.0245632
+ 5.94e+10Hz -0.0252352 0.0247065
+ 5.95e+10Hz -0.0253027 0.0248501
+ 5.96e+10Hz -0.02537 0.0249941
+ 5.97e+10Hz -0.025437 0.0251385
+ 5.98e+10Hz -0.0255037 0.0252832
+ 5.99e+10Hz -0.0255702 0.0254283
+ 6e+10Hz -0.0256365 0.0255738
+ 6.01e+10Hz -0.0257024 0.0257196
+ 6.02e+10Hz -0.0257681 0.0258658
+ 6.03e+10Hz -0.0258335 0.0260123
+ 6.04e+10Hz -0.0258986 0.0261592
+ 6.05e+10Hz -0.0259635 0.0263064
+ 6.06e+10Hz -0.0260281 0.0264541
+ 6.07e+10Hz -0.0260924 0.026602
+ 6.08e+10Hz -0.0261564 0.0267504
+ 6.09e+10Hz -0.0262202 0.0268991
+ 6.1e+10Hz -0.0262837 0.0270481
+ 6.11e+10Hz -0.0263469 0.0271975
+ 6.12e+10Hz -0.0264098 0.0273473
+ 6.13e+10Hz -0.0264724 0.0274974
+ 6.14e+10Hz -0.0265347 0.0276479
+ 6.15e+10Hz -0.0265968 0.0277987
+ 6.16e+10Hz -0.0266586 0.0279499
+ 6.17e+10Hz -0.02672 0.0281014
+ 6.18e+10Hz -0.0267812 0.0282533
+ 6.19e+10Hz -0.0268421 0.0284056
+ 6.2e+10Hz -0.0269027 0.0285582
+ 6.21e+10Hz -0.026963 0.0287111
+ 6.22e+10Hz -0.027023 0.0288644
+ 6.23e+10Hz -0.0270827 0.0290181
+ 6.24e+10Hz -0.0271421 0.0291721
+ 6.25e+10Hz -0.0272012 0.0293265
+ 6.26e+10Hz -0.0272601 0.0294812
+ 6.27e+10Hz -0.0273185 0.0296363
+ 6.28e+10Hz -0.0273767 0.0297917
+ 6.29e+10Hz -0.0274346 0.0299475
+ 6.3e+10Hz -0.0274922 0.0301036
+ 6.31e+10Hz -0.0275494 0.0302601
+ 6.32e+10Hz -0.0276064 0.030417
+ 6.33e+10Hz -0.027663 0.0305741
+ 6.34e+10Hz -0.0277193 0.0307316
+ 6.35e+10Hz -0.0277753 0.0308895
+ 6.36e+10Hz -0.027831 0.0310477
+ 6.37e+10Hz -0.0278864 0.0312063
+ 6.38e+10Hz -0.0279414 0.0313652
+ 6.39e+10Hz -0.0279961 0.0315245
+ 6.4e+10Hz -0.0280505 0.0316841
+ 6.41e+10Hz -0.0281045 0.031844
+ 6.42e+10Hz -0.0281583 0.0320043
+ 6.43e+10Hz -0.0282117 0.0321649
+ 6.44e+10Hz -0.0282647 0.0323259
+ 6.45e+10Hz -0.0283174 0.0324872
+ 6.46e+10Hz -0.0283698 0.0326489
+ 6.47e+10Hz -0.0284219 0.0328109
+ 6.48e+10Hz -0.0284736 0.0329732
+ 6.49e+10Hz -0.028525 0.0331359
+ 6.5e+10Hz -0.028576 0.0332989
+ 6.51e+10Hz -0.0286267 0.0334622
+ 6.52e+10Hz -0.028677 0.0336259
+ 6.53e+10Hz -0.028727 0.03379
+ 6.54e+10Hz -0.0287767 0.0339543
+ 6.55e+10Hz -0.0288259 0.034119
+ 6.56e+10Hz -0.0288749 0.0342841
+ 6.57e+10Hz -0.0289234 0.0344494
+ 6.58e+10Hz -0.0289717 0.0346151
+ 6.59e+10Hz -0.0290195 0.0347811
+ 6.6e+10Hz -0.029067 0.0349475
+ 6.61e+10Hz -0.0291142 0.0351142
+ 6.62e+10Hz -0.029161 0.0352812
+ 6.63e+10Hz -0.0292074 0.0354485
+ 6.64e+10Hz -0.0292534 0.0356162
+ 6.65e+10Hz -0.0292991 0.0357842
+ 6.66e+10Hz -0.0293444 0.0359525
+ 6.67e+10Hz -0.0293893 0.0361212
+ 6.68e+10Hz -0.0294339 0.0362902
+ 6.69e+10Hz -0.0294781 0.0364594
+ 6.7e+10Hz -0.0295219 0.0366291
+ 6.71e+10Hz -0.0295653 0.036799
+ 6.72e+10Hz -0.0296083 0.0369692
+ 6.73e+10Hz -0.029651 0.0371398
+ 6.74e+10Hz -0.0296933 0.0373107
+ 6.75e+10Hz -0.0297352 0.0374819
+ 6.76e+10Hz -0.0297767 0.0376534
+ 6.77e+10Hz -0.0298178 0.0378253
+ 6.78e+10Hz -0.0298585 0.0379974
+ 6.79e+10Hz -0.0298988 0.0381699
+ 6.8e+10Hz -0.0299387 0.0383426
+ 6.81e+10Hz -0.0299783 0.0385157
+ 6.82e+10Hz -0.0300174 0.0386891
+ 6.83e+10Hz -0.0300561 0.0388628
+ 6.84e+10Hz -0.0300944 0.0390368
+ 6.85e+10Hz -0.0301324 0.0392111
+ 6.86e+10Hz -0.0301699 0.0393857
+ 6.87e+10Hz -0.030207 0.0395606
+ 6.88e+10Hz -0.0302437 0.0397358
+ 6.89e+10Hz -0.03028 0.0399113
+ 6.9e+10Hz -0.0303159 0.0400871
+ 6.91e+10Hz -0.0303513 0.0402632
+ 6.92e+10Hz -0.0303864 0.0404396
+ 6.93e+10Hz -0.030421 0.0406163
+ 6.94e+10Hz -0.0304552 0.0407933
+ 6.95e+10Hz -0.030489 0.0409705
+ 6.96e+10Hz -0.0305224 0.0411481
+ 6.97e+10Hz -0.0305554 0.0413259
+ 6.98e+10Hz -0.0305879 0.0415041
+ 6.99e+10Hz -0.03062 0.0416825
+ 7e+10Hz -0.0306516 0.0418612
+ 7.01e+10Hz -0.0306829 0.0420402
+ 7.02e+10Hz -0.0307137 0.0422194
+ 7.03e+10Hz -0.0307441 0.042399
+ 7.04e+10Hz -0.030774 0.0425788
+ 7.05e+10Hz -0.0308035 0.0427589
+ 7.06e+10Hz -0.0308326 0.0429393
+ 7.07e+10Hz -0.0308612 0.0431199
+ 7.08e+10Hz -0.0308894 0.0433009
+ 7.09e+10Hz -0.0309171 0.043482
+ 7.1e+10Hz -0.0309444 0.0436635
+ 7.11e+10Hz -0.0309713 0.0438452
+ 7.12e+10Hz -0.0309977 0.0440272
+ 7.13e+10Hz -0.0310236 0.0442095
+ 7.14e+10Hz -0.0310491 0.044392
+ 7.15e+10Hz -0.0310742 0.0445748
+ 7.16e+10Hz -0.0310988 0.0447578
+ 7.17e+10Hz -0.031123 0.0449411
+ 7.18e+10Hz -0.0311467 0.0451246
+ 7.19e+10Hz -0.0311699 0.0453084
+ 7.2e+10Hz -0.0311927 0.0454925
+ 7.21e+10Hz -0.031215 0.0456768
+ 7.22e+10Hz -0.0312369 0.0458613
+ 7.23e+10Hz -0.0312583 0.0460461
+ 7.24e+10Hz -0.0312792 0.0462311
+ 7.25e+10Hz -0.0312997 0.0464164
+ 7.26e+10Hz -0.0313197 0.046602
+ 7.27e+10Hz -0.0313393 0.0467877
+ 7.28e+10Hz -0.0313583 0.0469737
+ 7.29e+10Hz -0.031377 0.04716
+ 7.3e+10Hz -0.0313951 0.0473464
+ 7.31e+10Hz -0.0314128 0.0475332
+ 7.32e+10Hz -0.03143 0.0477201
+ 7.33e+10Hz -0.0314467 0.0479073
+ 7.34e+10Hz -0.0314629 0.0480947
+ 7.35e+10Hz -0.0314787 0.0482823
+ 7.36e+10Hz -0.031494 0.0484701
+ 7.37e+10Hz -0.0315088 0.0486582
+ 7.38e+10Hz -0.0315232 0.0488465
+ 7.39e+10Hz -0.031537 0.049035
+ 7.4e+10Hz -0.0315504 0.0492237
+ 7.41e+10Hz -0.0315633 0.0494127
+ 7.42e+10Hz -0.0315757 0.0496018
+ 7.43e+10Hz -0.0315876 0.0497912
+ 7.44e+10Hz -0.0315991 0.0499808
+ 7.45e+10Hz -0.03161 0.0501706
+ 7.46e+10Hz -0.0316205 0.0503605
+ 7.47e+10Hz -0.0316305 0.0505507
+ 7.48e+10Hz -0.03164 0.0507411
+ 7.49e+10Hz -0.031649 0.0509317
+ 7.5e+10Hz -0.0316575 0.0511225
+ 7.51e+10Hz -0.0316655 0.0513135
+ 7.52e+10Hz -0.031673 0.0515047
+ 7.53e+10Hz -0.0316801 0.0516961
+ 7.54e+10Hz -0.0316866 0.0518877
+ 7.55e+10Hz -0.0316927 0.0520794
+ 7.56e+10Hz -0.0316982 0.0522714
+ 7.57e+10Hz -0.0317033 0.0524635
+ 7.58e+10Hz -0.0317078 0.0526559
+ 7.59e+10Hz -0.0317119 0.0528484
+ 7.6e+10Hz -0.0317154 0.053041
+ 7.61e+10Hz -0.0317185 0.0532339
+ 7.62e+10Hz -0.031721 0.053427
+ 7.63e+10Hz -0.0317231 0.0536202
+ 7.64e+10Hz -0.0317246 0.0538136
+ 7.65e+10Hz -0.0317257 0.0540071
+ 7.66e+10Hz -0.0317262 0.0542009
+ 7.67e+10Hz -0.0317263 0.0543948
+ 7.68e+10Hz -0.0317258 0.0545889
+ 7.69e+10Hz -0.0317248 0.0547831
+ 7.7e+10Hz -0.0317234 0.0549775
+ 7.71e+10Hz -0.0317214 0.0551721
+ 7.72e+10Hz -0.0317189 0.0553668
+ 7.73e+10Hz -0.0317159 0.0555617
+ 7.74e+10Hz -0.0317124 0.0557567
+ 7.75e+10Hz -0.0317084 0.0559519
+ 7.76e+10Hz -0.0317039 0.0561473
+ 7.77e+10Hz -0.0316988 0.0563427
+ 7.78e+10Hz -0.0316933 0.0565384
+ 7.79e+10Hz -0.0316872 0.0567342
+ 7.8e+10Hz -0.0316806 0.0569301
+ 7.81e+10Hz -0.0316736 0.0571262
+ 7.82e+10Hz -0.031666 0.0573224
+ 7.83e+10Hz -0.0316579 0.0575188
+ 7.84e+10Hz -0.0316492 0.0577153
+ 7.85e+10Hz -0.0316401 0.057912
+ 7.86e+10Hz -0.0316304 0.0581087
+ 7.87e+10Hz -0.0316203 0.0583057
+ 7.88e+10Hz -0.0316096 0.0585027
+ 7.89e+10Hz -0.0315983 0.0586999
+ 7.9e+10Hz -0.0315866 0.0588972
+ 7.91e+10Hz -0.0315744 0.0590946
+ 7.92e+10Hz -0.0315616 0.0592922
+ 7.93e+10Hz -0.0315483 0.0594899
+ 7.94e+10Hz -0.0315345 0.0596877
+ 7.95e+10Hz -0.0315202 0.0598856
+ 7.96e+10Hz -0.0315054 0.0600837
+ 7.97e+10Hz -0.03149 0.0602818
+ 7.98e+10Hz -0.0314741 0.0604801
+ 7.99e+10Hz -0.0314577 0.0606785
+ 8e+10Hz -0.0314408 0.0608771
+ 8.01e+10Hz -0.0314233 0.0610757
+ 8.02e+10Hz -0.0314054 0.0612744
+ 8.03e+10Hz -0.0313869 0.0614733
+ 8.04e+10Hz -0.0313678 0.0616722
+ 8.05e+10Hz -0.0313483 0.0618713
+ 8.06e+10Hz -0.0313282 0.0620704
+ 8.07e+10Hz -0.0313076 0.0622697
+ 8.08e+10Hz -0.0312865 0.0624691
+ 8.09e+10Hz -0.0312648 0.0626685
+ 8.1e+10Hz -0.0312427 0.0628681
+ 8.11e+10Hz -0.0312199 0.0630678
+ 8.12e+10Hz -0.0311967 0.0632675
+ 8.13e+10Hz -0.031173 0.0634674
+ 8.14e+10Hz -0.0311487 0.0636673
+ 8.15e+10Hz -0.0311238 0.0638673
+ 8.16e+10Hz -0.0310985 0.0640675
+ 8.17e+10Hz -0.0310726 0.0642677
+ 8.18e+10Hz -0.0310462 0.064468
+ 8.19e+10Hz -0.0310193 0.0646683
+ 8.2e+10Hz -0.0309918 0.0648688
+ 8.21e+10Hz -0.0309638 0.0650693
+ 8.22e+10Hz -0.0309352 0.06527
+ 8.23e+10Hz -0.0309062 0.0654707
+ 8.24e+10Hz -0.0308766 0.0656715
+ 8.25e+10Hz -0.0308464 0.0658723
+ 8.26e+10Hz -0.0308157 0.0660732
+ 8.27e+10Hz -0.0307846 0.0662742
+ 8.28e+10Hz -0.0307528 0.0664753
+ 8.29e+10Hz -0.0307205 0.0666765
+ 8.3e+10Hz -0.0306877 0.0668777
+ 8.31e+10Hz -0.0306544 0.0670789
+ 8.32e+10Hz -0.0306205 0.0672803
+ 8.33e+10Hz -0.0305861 0.0674817
+ 8.34e+10Hz -0.0305511 0.0676832
+ 8.35e+10Hz -0.0305156 0.0678847
+ 8.36e+10Hz -0.0304796 0.0680863
+ 8.37e+10Hz -0.030443 0.068288
+ 8.38e+10Hz -0.0304059 0.0684897
+ 8.39e+10Hz -0.0303682 0.0686914
+ 8.4e+10Hz -0.03033 0.0688933
+ 8.41e+10Hz -0.0302913 0.0690951
+ 8.42e+10Hz -0.030252 0.0692971
+ 8.43e+10Hz -0.0302122 0.069499
+ 8.44e+10Hz -0.0301718 0.0697011
+ 8.45e+10Hz -0.0301309 0.0699031
+ 8.46e+10Hz -0.0300894 0.0701052
+ 8.47e+10Hz -0.0300474 0.0703074
+ 8.48e+10Hz -0.0300049 0.0705096
+ 8.49e+10Hz -0.0299618 0.0707119
+ 8.5e+10Hz -0.0299182 0.0709141
+ 8.51e+10Hz -0.029874 0.0711165
+ 8.52e+10Hz -0.0298293 0.0713188
+ 8.53e+10Hz -0.029784 0.0715212
+ 8.54e+10Hz -0.0297382 0.0717236
+ 8.55e+10Hz -0.0296918 0.0719261
+ 8.56e+10Hz -0.0296449 0.0721286
+ 8.57e+10Hz -0.0295974 0.0723311
+ 8.58e+10Hz -0.0295494 0.0725337
+ 8.59e+10Hz -0.0295008 0.0727363
+ 8.6e+10Hz -0.0294517 0.0729389
+ 8.61e+10Hz -0.029402 0.0731415
+ 8.62e+10Hz -0.0293518 0.0733442
+ 8.63e+10Hz -0.029301 0.0735468
+ 8.64e+10Hz -0.0292496 0.0737495
+ 8.65e+10Hz -0.0291978 0.0739522
+ 8.66e+10Hz -0.0291453 0.074155
+ 8.67e+10Hz -0.0290923 0.0743577
+ 8.68e+10Hz -0.0290387 0.0745605
+ 8.69e+10Hz -0.0289846 0.0747633
+ 8.7e+10Hz -0.0289299 0.074966
+ 8.71e+10Hz -0.0288747 0.0751688
+ 8.72e+10Hz -0.0288189 0.0753716
+ 8.73e+10Hz -0.0287626 0.0755744
+ 8.74e+10Hz -0.0287057 0.0757772
+ 8.75e+10Hz -0.0286482 0.07598
+ 8.76e+10Hz -0.0285902 0.0761828
+ 8.77e+10Hz -0.0285316 0.0763857
+ 8.78e+10Hz -0.0284724 0.0765885
+ 8.79e+10Hz -0.0284127 0.0767913
+ 8.8e+10Hz -0.0283524 0.0769941
+ 8.81e+10Hz -0.0282916 0.0771969
+ 8.82e+10Hz -0.0282302 0.0773997
+ 8.83e+10Hz -0.0281682 0.0776024
+ 8.84e+10Hz -0.0281056 0.0778052
+ 8.85e+10Hz -0.0280425 0.078008
+ 8.86e+10Hz -0.0279788 0.0782107
+ 8.87e+10Hz -0.0279146 0.0784134
+ 8.88e+10Hz -0.0278498 0.0786161
+ 8.89e+10Hz -0.0277844 0.0788188
+ 8.9e+10Hz -0.0277184 0.0790215
+ 8.91e+10Hz -0.0276519 0.0792241
+ 8.92e+10Hz -0.0275848 0.0794267
+ 8.93e+10Hz -0.0275172 0.0796293
+ 8.94e+10Hz -0.0274489 0.0798318
+ 8.95e+10Hz -0.0273801 0.0800344
+ 8.96e+10Hz -0.0273107 0.0802369
+ 8.97e+10Hz -0.0272408 0.0804393
+ 8.98e+10Hz -0.0271702 0.0806418
+ 8.99e+10Hz -0.0270991 0.0808442
+ 9e+10Hz -0.0270274 0.0810465
+ 9.01e+10Hz -0.0269551 0.0812488
+ 9.02e+10Hz -0.0268823 0.0814511
+ 9.03e+10Hz -0.0268089 0.0816533
+ 9.04e+10Hz -0.0267349 0.0818555
+ 9.05e+10Hz -0.0266603 0.0820576
+ 9.06e+10Hz -0.0265851 0.0822597
+ 9.07e+10Hz -0.0265094 0.0824617
+ 9.08e+10Hz -0.0264331 0.0826637
+ 9.09e+10Hz -0.0263562 0.0828656
+ 9.1e+10Hz -0.0262787 0.0830674
+ 9.11e+10Hz -0.0262006 0.0832692
+ 9.12e+10Hz -0.026122 0.083471
+ 9.13e+10Hz -0.0260427 0.0836727
+ 9.14e+10Hz -0.0259629 0.0838743
+ 9.15e+10Hz -0.0258825 0.0840758
+ 9.16e+10Hz -0.0258015 0.0842773
+ 9.17e+10Hz -0.0257199 0.0844787
+ 9.18e+10Hz -0.0256378 0.08468
+ 9.19e+10Hz -0.025555 0.0848813
+ 9.2e+10Hz -0.0254717 0.0850824
+ 9.21e+10Hz -0.0253878 0.0852835
+ 9.22e+10Hz -0.0253032 0.0854845
+ 9.23e+10Hz -0.0252181 0.0856855
+ 9.24e+10Hz -0.0251325 0.0858863
+ 9.25e+10Hz -0.0250462 0.0860871
+ 9.26e+10Hz -0.0249593 0.0862877
+ 9.27e+10Hz -0.0248718 0.0864883
+ 9.28e+10Hz -0.0247838 0.0866888
+ 9.29e+10Hz -0.0246951 0.0868892
+ 9.3e+10Hz -0.0246059 0.0870894
+ 9.31e+10Hz -0.0245161 0.0872896
+ 9.32e+10Hz -0.0244257 0.0874897
+ 9.33e+10Hz -0.0243346 0.0876897
+ 9.34e+10Hz -0.024243 0.0878896
+ 9.35e+10Hz -0.0241508 0.0880893
+ 9.36e+10Hz -0.024058 0.088289
+ 9.37e+10Hz -0.0239646 0.0884885
+ 9.38e+10Hz -0.0238707 0.088688
+ 9.39e+10Hz -0.0237761 0.0888873
+ 9.4e+10Hz -0.0236809 0.0890864
+ 9.41e+10Hz -0.0235851 0.0892855
+ 9.42e+10Hz -0.0234888 0.0894844
+ 9.43e+10Hz -0.0233918 0.0896833
+ 9.44e+10Hz -0.0232942 0.089882
+ 9.45e+10Hz -0.0231961 0.0900805
+ 9.46e+10Hz -0.0230973 0.0902789
+ 9.47e+10Hz -0.022998 0.0904772
+ 9.48e+10Hz -0.022898 0.0906754
+ 9.49e+10Hz -0.0227975 0.0908734
+ 9.5e+10Hz -0.0226964 0.0910712
+ 9.51e+10Hz -0.0225946 0.091269
+ 9.52e+10Hz -0.0224923 0.0914665
+ 9.53e+10Hz -0.0223893 0.0916639
+ 9.54e+10Hz -0.0222858 0.0918612
+ 9.55e+10Hz -0.0221817 0.0920583
+ 9.56e+10Hz -0.022077 0.0922553
+ 9.57e+10Hz -0.0219716 0.0924521
+ 9.58e+10Hz -0.0218657 0.0926488
+ 9.59e+10Hz -0.0217592 0.0928452
+ 9.6e+10Hz -0.0216521 0.0930416
+ 9.61e+10Hz -0.0215444 0.0932377
+ 9.62e+10Hz -0.0214361 0.0934337
+ 9.63e+10Hz -0.0213271 0.0936295
+ 9.64e+10Hz -0.0212176 0.0938251
+ 9.65e+10Hz -0.0211075 0.0940206
+ 9.66e+10Hz -0.0209968 0.0942159
+ 9.67e+10Hz -0.0208855 0.0944109
+ 9.68e+10Hz -0.0207736 0.0946059
+ 9.69e+10Hz -0.0206611 0.0948006
+ 9.7e+10Hz -0.020548 0.0949951
+ 9.71e+10Hz -0.0204343 0.0951894
+ 9.72e+10Hz -0.02032 0.0953836
+ 9.73e+10Hz -0.0202052 0.0955776
+ 9.74e+10Hz -0.0200897 0.0957713
+ 9.75e+10Hz -0.0199736 0.0959649
+ 9.76e+10Hz -0.019857 0.0961582
+ 9.77e+10Hz -0.0197397 0.0963514
+ 9.78e+10Hz -0.0196218 0.0965443
+ 9.79e+10Hz -0.0195034 0.0967371
+ 9.8e+10Hz -0.0193843 0.0969296
+ 9.81e+10Hz -0.0192647 0.0971219
+ 9.82e+10Hz -0.0191444 0.097314
+ 9.83e+10Hz -0.0190236 0.0975059
+ 9.84e+10Hz -0.0189022 0.0976975
+ 9.85e+10Hz -0.0187801 0.0978889
+ 9.86e+10Hz -0.0186575 0.0980801
+ 9.87e+10Hz -0.0185343 0.0982711
+ 9.88e+10Hz -0.0184106 0.0984618
+ 9.89e+10Hz -0.0182862 0.0986523
+ 9.9e+10Hz -0.0181612 0.0988426
+ 9.91e+10Hz -0.0180356 0.0990327
+ 9.92e+10Hz -0.0179095 0.0992225
+ 9.93e+10Hz -0.0177827 0.099412
+ 9.94e+10Hz -0.0176554 0.0996013
+ 9.95e+10Hz -0.0175275 0.0997904
+ 9.96e+10Hz -0.017399 0.0999792
+ 9.97e+10Hz -0.0172699 0.100168
+ 9.98e+10Hz -0.0171402 0.100356
+ 9.99e+10Hz -0.0170099 0.100544
+ 1e+11Hz -0.0168791 0.100732
+ 1.001e+11Hz -0.0167476 0.100919
+ 1.002e+11Hz -0.0166156 0.101107
+ 1.003e+11Hz -0.016483 0.101294
+ 1.004e+11Hz -0.0163498 0.101481
+ 1.005e+11Hz -0.0162161 0.101667
+ 1.006e+11Hz -0.0160817 0.101853
+ 1.007e+11Hz -0.0159468 0.102039
+ 1.008e+11Hz -0.0158113 0.102225
+ 1.009e+11Hz -0.0156752 0.10241
+ 1.01e+11Hz -0.0155385 0.102595
+ 1.011e+11Hz -0.0154013 0.10278
+ 1.012e+11Hz -0.0152635 0.102965
+ 1.013e+11Hz -0.0151251 0.103149
+ 1.014e+11Hz -0.0149861 0.103333
+ 1.015e+11Hz -0.0148466 0.103517
+ 1.016e+11Hz -0.0147064 0.1037
+ 1.017e+11Hz -0.0145658 0.103883
+ 1.018e+11Hz -0.0144245 0.104066
+ 1.019e+11Hz -0.0142827 0.104248
+ 1.02e+11Hz -0.0141403 0.10443
+ 1.021e+11Hz -0.0139973 0.104612
+ 1.022e+11Hz -0.0138537 0.104794
+ 1.023e+11Hz -0.0137096 0.104975
+ 1.024e+11Hz -0.0135649 0.105156
+ 1.025e+11Hz -0.0134197 0.105337
+ 1.026e+11Hz -0.0132739 0.105517
+ 1.027e+11Hz -0.0131275 0.105697
+ 1.028e+11Hz -0.0129806 0.105877
+ 1.029e+11Hz -0.0128331 0.106056
+ 1.03e+11Hz -0.012685 0.106235
+ 1.031e+11Hz -0.0125364 0.106414
+ 1.032e+11Hz -0.0123872 0.106593
+ 1.033e+11Hz -0.0122375 0.106771
+ 1.034e+11Hz -0.0120872 0.106949
+ 1.035e+11Hz -0.0119363 0.107126
+ 1.036e+11Hz -0.0117849 0.107303
+ 1.037e+11Hz -0.0116329 0.10748
+ 1.038e+11Hz -0.0114804 0.107656
+ 1.039e+11Hz -0.0113273 0.107832
+ 1.04e+11Hz -0.0111737 0.108008
+ 1.041e+11Hz -0.0110195 0.108184
+ 1.042e+11Hz -0.0108648 0.108359
+ 1.043e+11Hz -0.0107095 0.108534
+ 1.044e+11Hz -0.0105536 0.108708
+ 1.045e+11Hz -0.0103973 0.108882
+ 1.046e+11Hz -0.0102403 0.109056
+ 1.047e+11Hz -0.0100829 0.109229
+ 1.048e+11Hz -0.00992485 0.109402
+ 1.049e+11Hz -0.00976628 0.109575
+ 1.05e+11Hz -0.00960718 0.109747
+ 1.051e+11Hz -0.00944753 0.109919
+ 1.052e+11Hz -0.00928734 0.11009
+ 1.053e+11Hz -0.0091266 0.110262
+ 1.054e+11Hz -0.00896533 0.110433
+ 1.055e+11Hz -0.00880352 0.110603
+ 1.056e+11Hz -0.00864118 0.110773
+ 1.057e+11Hz -0.00847829 0.110943
+ 1.058e+11Hz -0.00831487 0.111112
+ 1.059e+11Hz -0.00815092 0.111281
+ 1.06e+11Hz -0.00798643 0.11145
+ 1.061e+11Hz -0.00782141 0.111618
+ 1.062e+11Hz -0.00765585 0.111786
+ 1.063e+11Hz -0.00748977 0.111953
+ 1.064e+11Hz -0.00732316 0.11212
+ 1.065e+11Hz -0.00715601 0.112287
+ 1.066e+11Hz -0.00698834 0.112454
+ 1.067e+11Hz -0.00682014 0.112619
+ 1.068e+11Hz -0.00665141 0.112785
+ 1.069e+11Hz -0.00648216 0.11295
+ 1.07e+11Hz -0.00631239 0.113115
+ 1.071e+11Hz -0.00614209 0.11328
+ 1.072e+11Hz -0.00597126 0.113444
+ 1.073e+11Hz -0.00579992 0.113607
+ 1.074e+11Hz -0.00562806 0.11377
+ 1.075e+11Hz -0.00545567 0.113933
+ 1.076e+11Hz -0.00528277 0.114096
+ 1.077e+11Hz -0.00510934 0.114257
+ 1.078e+11Hz -0.0049354 0.114419
+ 1.079e+11Hz -0.00476094 0.11458
+ 1.08e+11Hz -0.00458597 0.114741
+ 1.081e+11Hz -0.00441048 0.114902
+ 1.082e+11Hz -0.00423448 0.115061
+ 1.083e+11Hz -0.00405797 0.115221
+ 1.084e+11Hz -0.00388094 0.11538
+ 1.085e+11Hz -0.0037034 0.115539
+ 1.086e+11Hz -0.00352535 0.115697
+ 1.087e+11Hz -0.0033468 0.115855
+ 1.088e+11Hz -0.00316773 0.116013
+ 1.089e+11Hz -0.00298816 0.11617
+ 1.09e+11Hz -0.00280807 0.116326
+ 1.091e+11Hz -0.00262748 0.116483
+ 1.092e+11Hz -0.00244639 0.116639
+ 1.093e+11Hz -0.00226479 0.116794
+ 1.094e+11Hz -0.00208269 0.116949
+ 1.095e+11Hz -0.00190008 0.117103
+ 1.096e+11Hz -0.00171697 0.117258
+ 1.097e+11Hz -0.00153336 0.117411
+ 1.098e+11Hz -0.00134925 0.117564
+ 1.099e+11Hz -0.00116464 0.117717
+ 1.1e+11Hz -0.000979534 0.11787
+ 1.101e+11Hz -0.000793926 0.118022
+ 1.102e+11Hz -0.00060782 0.118173
+ 1.103e+11Hz -0.000421218 0.118324
+ 1.104e+11Hz -0.00023412 0.118475
+ 1.105e+11Hz -4.6527e-05 0.118625
+ 1.106e+11Hz 0.000141561 0.118774
+ 1.107e+11Hz 0.000330142 0.118924
+ 1.108e+11Hz 0.000519217 0.119072
+ 1.109e+11Hz 0.000708783 0.119221
+ 1.11e+11Hz 0.000898841 0.119369
+ 1.111e+11Hz 0.00108939 0.119516
+ 1.112e+11Hz 0.00128043 0.119663
+ 1.113e+11Hz 0.00147196 0.11981
+ 1.114e+11Hz 0.00166397 0.119956
+ 1.115e+11Hz 0.00185648 0.120101
+ 1.116e+11Hz 0.00204947 0.120247
+ 1.117e+11Hz 0.00224295 0.120391
+ 1.118e+11Hz 0.00243691 0.120536
+ 1.119e+11Hz 0.00263136 0.120679
+ 1.12e+11Hz 0.00282629 0.120822
+ 1.121e+11Hz 0.0030217 0.120965
+ 1.122e+11Hz 0.0032176 0.121108
+ 1.123e+11Hz 0.00341398 0.121249
+ 1.124e+11Hz 0.00361084 0.121391
+ 1.125e+11Hz 0.00380818 0.121532
+ 1.126e+11Hz 0.004006 0.121672
+ 1.127e+11Hz 0.0042043 0.121812
+ 1.128e+11Hz 0.00440307 0.121952
+ 1.129e+11Hz 0.00460233 0.122091
+ 1.13e+11Hz 0.00480206 0.122229
+ 1.131e+11Hz 0.00500226 0.122367
+ 1.132e+11Hz 0.00520295 0.122505
+ 1.133e+11Hz 0.0054041 0.122642
+ 1.134e+11Hz 0.00560573 0.122778
+ 1.135e+11Hz 0.00580783 0.122914
+ 1.136e+11Hz 0.00601041 0.12305
+ 1.137e+11Hz 0.00621345 0.123185
+ 1.138e+11Hz 0.00641697 0.12332
+ 1.139e+11Hz 0.00662096 0.123454
+ 1.14e+11Hz 0.00682541 0.123587
+ 1.141e+11Hz 0.00703034 0.12372
+ 1.142e+11Hz 0.00723573 0.123853
+ 1.143e+11Hz 0.00744159 0.123985
+ 1.144e+11Hz 0.00764791 0.124116
+ 1.145e+11Hz 0.0078547 0.124247
+ 1.146e+11Hz 0.00806195 0.124378
+ 1.147e+11Hz 0.00826967 0.124508
+ 1.148e+11Hz 0.00847785 0.124637
+ 1.149e+11Hz 0.00868649 0.124766
+ 1.15e+11Hz 0.00889559 0.124895
+ 1.151e+11Hz 0.00910515 0.125023
+ 1.152e+11Hz 0.00931517 0.12515
+ 1.153e+11Hz 0.00952565 0.125277
+ 1.154e+11Hz 0.00973659 0.125403
+ 1.155e+11Hz 0.00994798 0.125529
+ 1.156e+11Hz 0.0101598 0.125654
+ 1.157e+11Hz 0.0103721 0.125779
+ 1.158e+11Hz 0.0105849 0.125903
+ 1.159e+11Hz 0.0107981 0.126027
+ 1.16e+11Hz 0.0110118 0.12615
+ 1.161e+11Hz 0.0112259 0.126272
+ 1.162e+11Hz 0.0114404 0.126394
+ 1.163e+11Hz 0.0116555 0.126516
+ 1.164e+11Hz 0.0118709 0.126637
+ 1.165e+11Hz 0.0120868 0.126757
+ 1.166e+11Hz 0.0123032 0.126877
+ 1.167e+11Hz 0.01252 0.126996
+ 1.168e+11Hz 0.0127372 0.127115
+ 1.169e+11Hz 0.0129549 0.127233
+ 1.17e+11Hz 0.013173 0.127351
+ 1.171e+11Hz 0.0133916 0.127468
+ 1.172e+11Hz 0.0136106 0.127584
+ 1.173e+11Hz 0.0138301 0.1277
+ 1.174e+11Hz 0.01405 0.127815
+ 1.175e+11Hz 0.0142703 0.12793
+ 1.176e+11Hz 0.014491 0.128044
+ 1.177e+11Hz 0.0147122 0.128158
+ 1.178e+11Hz 0.0149339 0.128271
+ 1.179e+11Hz 0.0151559 0.128383
+ 1.18e+11Hz 0.0153784 0.128495
+ 1.181e+11Hz 0.0156013 0.128606
+ 1.182e+11Hz 0.0158246 0.128717
+ 1.183e+11Hz 0.0160484 0.128827
+ 1.184e+11Hz 0.0162726 0.128936
+ 1.185e+11Hz 0.0164972 0.129045
+ 1.186e+11Hz 0.0167223 0.129154
+ 1.187e+11Hz 0.0169478 0.129261
+ 1.188e+11Hz 0.0171736 0.129368
+ 1.189e+11Hz 0.0173999 0.129475
+ 1.19e+11Hz 0.0176267 0.129581
+ 1.191e+11Hz 0.0178538 0.129686
+ 1.192e+11Hz 0.0180814 0.129791
+ 1.193e+11Hz 0.0183093 0.129895
+ 1.194e+11Hz 0.0185377 0.129998
+ 1.195e+11Hz 0.0187665 0.130101
+ 1.196e+11Hz 0.0189957 0.130203
+ 1.197e+11Hz 0.0192253 0.130305
+ 1.198e+11Hz 0.0194553 0.130406
+ 1.199e+11Hz 0.0196857 0.130506
+ 1.2e+11Hz 0.0199165 0.130606
+ 1.201e+11Hz 0.0201478 0.130705
+ 1.202e+11Hz 0.0203794 0.130804
+ 1.203e+11Hz 0.0206114 0.130902
+ 1.204e+11Hz 0.0208438 0.130999
+ 1.205e+11Hz 0.0210766 0.131095
+ 1.206e+11Hz 0.0213098 0.131191
+ 1.207e+11Hz 0.0215434 0.131287
+ 1.208e+11Hz 0.0217774 0.131381
+ 1.209e+11Hz 0.0220118 0.131475
+ 1.21e+11Hz 0.0222465 0.131569
+ 1.211e+11Hz 0.0224816 0.131661
+ 1.212e+11Hz 0.0227172 0.131753
+ 1.213e+11Hz 0.0229531 0.131845
+ 1.214e+11Hz 0.0231894 0.131936
+ 1.215e+11Hz 0.023426 0.132026
+ 1.216e+11Hz 0.0236631 0.132115
+ 1.217e+11Hz 0.0239005 0.132204
+ 1.218e+11Hz 0.0241382 0.132292
+ 1.219e+11Hz 0.0243764 0.13238
+ 1.22e+11Hz 0.0246149 0.132466
+ 1.221e+11Hz 0.0248538 0.132552
+ 1.222e+11Hz 0.025093 0.132638
+ 1.223e+11Hz 0.0253326 0.132723
+ 1.224e+11Hz 0.0255726 0.132807
+ 1.225e+11Hz 0.0258129 0.13289
+ 1.226e+11Hz 0.0260536 0.132973
+ 1.227e+11Hz 0.0262946 0.133055
+ 1.228e+11Hz 0.026536 0.133136
+ 1.229e+11Hz 0.0267777 0.133217
+ 1.23e+11Hz 0.0270198 0.133297
+ 1.231e+11Hz 0.0272622 0.133377
+ 1.232e+11Hz 0.027505 0.133455
+ 1.233e+11Hz 0.0277481 0.133533
+ 1.234e+11Hz 0.0279916 0.13361
+ 1.235e+11Hz 0.0282354 0.133687
+ 1.236e+11Hz 0.0284795 0.133763
+ 1.237e+11Hz 0.0287239 0.133838
+ 1.238e+11Hz 0.0289687 0.133912
+ 1.239e+11Hz 0.0292138 0.133986
+ 1.24e+11Hz 0.0294592 0.134059
+ 1.241e+11Hz 0.029705 0.134132
+ 1.242e+11Hz 0.0299511 0.134203
+ 1.243e+11Hz 0.0301975 0.134274
+ 1.244e+11Hz 0.0304442 0.134345
+ 1.245e+11Hz 0.0306912 0.134414
+ 1.246e+11Hz 0.0309386 0.134483
+ 1.247e+11Hz 0.0311862 0.134551
+ 1.248e+11Hz 0.0314342 0.134618
+ 1.249e+11Hz 0.0316824 0.134685
+ 1.25e+11Hz 0.031931 0.134751
+ 1.251e+11Hz 0.0321799 0.134816
+ 1.252e+11Hz 0.032429 0.134881
+ 1.253e+11Hz 0.0326785 0.134944
+ 1.254e+11Hz 0.0329282 0.135007
+ 1.255e+11Hz 0.0331783 0.13507
+ 1.256e+11Hz 0.0334286 0.135131
+ 1.257e+11Hz 0.0336792 0.135192
+ 1.258e+11Hz 0.0339301 0.135252
+ 1.259e+11Hz 0.0341813 0.135312
+ 1.26e+11Hz 0.0344327 0.13537
+ 1.261e+11Hz 0.0346845 0.135428
+ 1.262e+11Hz 0.0349365 0.135486
+ 1.263e+11Hz 0.0351888 0.135542
+ 1.264e+11Hz 0.0354413 0.135598
+ 1.265e+11Hz 0.0356941 0.135653
+ 1.266e+11Hz 0.0359472 0.135707
+ 1.267e+11Hz 0.0362005 0.13576
+ 1.268e+11Hz 0.0364541 0.135813
+ 1.269e+11Hz 0.036708 0.135865
+ 1.27e+11Hz 0.0369621 0.135916
+ 1.271e+11Hz 0.0372165 0.135967
+ 1.272e+11Hz 0.0374711 0.136017
+ 1.273e+11Hz 0.0377259 0.136066
+ 1.274e+11Hz 0.037981 0.136114
+ 1.275e+11Hz 0.0382364 0.136161
+ 1.276e+11Hz 0.038492 0.136208
+ 1.277e+11Hz 0.0387478 0.136254
+ 1.278e+11Hz 0.0390038 0.136299
+ 1.279e+11Hz 0.0392601 0.136344
+ 1.28e+11Hz 0.0395167 0.136387
+ 1.281e+11Hz 0.0397734 0.136431
+ 1.282e+11Hz 0.0400304 0.136473
+ 1.283e+11Hz 0.0402876 0.136514
+ 1.284e+11Hz 0.040545 0.136555
+ 1.285e+11Hz 0.0408026 0.136595
+ 1.286e+11Hz 0.0410605 0.136634
+ 1.287e+11Hz 0.0413185 0.136672
+ 1.288e+11Hz 0.0415768 0.13671
+ 1.289e+11Hz 0.0418353 0.136747
+ 1.29e+11Hz 0.042094 0.136783
+ 1.291e+11Hz 0.0423529 0.136818
+ 1.292e+11Hz 0.042612 0.136853
+ 1.293e+11Hz 0.0428712 0.136887
+ 1.294e+11Hz 0.0431307 0.13692
+ 1.295e+11Hz 0.0433904 0.136952
+ 1.296e+11Hz 0.0436503 0.136984
+ 1.297e+11Hz 0.0439104 0.137014
+ 1.298e+11Hz 0.0441706 0.137044
+ 1.299e+11Hz 0.044431 0.137073
+ 1.3e+11Hz 0.0446917 0.137102
+ 1.301e+11Hz 0.0449525 0.13713
+ 1.302e+11Hz 0.0452135 0.137156
+ 1.303e+11Hz 0.0454746 0.137183
+ 1.304e+11Hz 0.0457359 0.137208
+ 1.305e+11Hz 0.0459974 0.137233
+ 1.306e+11Hz 0.0462591 0.137256
+ 1.307e+11Hz 0.0465209 0.137279
+ 1.308e+11Hz 0.0467829 0.137301
+ 1.309e+11Hz 0.0470451 0.137323
+ 1.31e+11Hz 0.0473074 0.137344
+ 1.311e+11Hz 0.0475699 0.137363
+ 1.312e+11Hz 0.0478326 0.137383
+ 1.313e+11Hz 0.0480954 0.137401
+ 1.314e+11Hz 0.0483583 0.137419
+ 1.315e+11Hz 0.0486214 0.137435
+ 1.316e+11Hz 0.0488846 0.137451
+ 1.317e+11Hz 0.049148 0.137467
+ 1.318e+11Hz 0.0494116 0.137481
+ 1.319e+11Hz 0.0496752 0.137495
+ 1.32e+11Hz 0.0499391 0.137508
+ 1.321e+11Hz 0.050203 0.13752
+ 1.322e+11Hz 0.0504671 0.137531
+ 1.323e+11Hz 0.0507313 0.137542
+ 1.324e+11Hz 0.0509957 0.137551
+ 1.325e+11Hz 0.0512602 0.13756
+ 1.326e+11Hz 0.0515248 0.137568
+ 1.327e+11Hz 0.0517895 0.137576
+ 1.328e+11Hz 0.0520544 0.137582
+ 1.329e+11Hz 0.0523194 0.137588
+ 1.33e+11Hz 0.0525845 0.137593
+ 1.331e+11Hz 0.0528497 0.137597
+ 1.332e+11Hz 0.0531151 0.137601
+ 1.333e+11Hz 0.0533805 0.137604
+ 1.334e+11Hz 0.0536461 0.137605
+ 1.335e+11Hz 0.0539118 0.137607
+ 1.336e+11Hz 0.0541776 0.137607
+ 1.337e+11Hz 0.0544435 0.137606
+ 1.338e+11Hz 0.0547095 0.137605
+ 1.339e+11Hz 0.0549756 0.137603
+ 1.34e+11Hz 0.0552418 0.1376
+ 1.341e+11Hz 0.0555081 0.137597
+ 1.342e+11Hz 0.0557745 0.137592
+ 1.343e+11Hz 0.0560411 0.137587
+ 1.344e+11Hz 0.0563077 0.137581
+ 1.345e+11Hz 0.0565744 0.137574
+ 1.346e+11Hz 0.0568412 0.137567
+ 1.347e+11Hz 0.0571081 0.137558
+ 1.348e+11Hz 0.057375 0.137549
+ 1.349e+11Hz 0.0576421 0.137539
+ 1.35e+11Hz 0.0579092 0.137528
+ 1.351e+11Hz 0.0581764 0.137517
+ 1.352e+11Hz 0.0584438 0.137504
+ 1.353e+11Hz 0.0587111 0.137491
+ 1.354e+11Hz 0.0589786 0.137477
+ 1.355e+11Hz 0.0592462 0.137462
+ 1.356e+11Hz 0.0595138 0.137447
+ 1.357e+11Hz 0.0597815 0.13743
+ 1.358e+11Hz 0.0600493 0.137413
+ 1.359e+11Hz 0.0603171 0.137395
+ 1.36e+11Hz 0.060585 0.137377
+ 1.361e+11Hz 0.060853 0.137357
+ 1.362e+11Hz 0.061121 0.137337
+ 1.363e+11Hz 0.0613892 0.137315
+ 1.364e+11Hz 0.0616573 0.137293
+ 1.365e+11Hz 0.0619256 0.137271
+ 1.366e+11Hz 0.0621939 0.137247
+ 1.367e+11Hz 0.0624622 0.137223
+ 1.368e+11Hz 0.0627306 0.137198
+ 1.369e+11Hz 0.0629991 0.137172
+ 1.37e+11Hz 0.0632676 0.137145
+ 1.371e+11Hz 0.0635362 0.137117
+ 1.372e+11Hz 0.0638048 0.137089
+ 1.373e+11Hz 0.0640735 0.137059
+ 1.374e+11Hz 0.0643422 0.137029
+ 1.375e+11Hz 0.064611 0.136998
+ 1.376e+11Hz 0.0648798 0.136967
+ 1.377e+11Hz 0.0651487 0.136934
+ 1.378e+11Hz 0.0654175 0.136901
+ 1.379e+11Hz 0.0656865 0.136867
+ 1.38e+11Hz 0.0659555 0.136832
+ 1.381e+11Hz 0.0662245 0.136796
+ 1.382e+11Hz 0.0664935 0.13676
+ 1.383e+11Hz 0.0667626 0.136722
+ 1.384e+11Hz 0.0670317 0.136684
+ 1.385e+11Hz 0.0673009 0.136645
+ 1.386e+11Hz 0.06757 0.136605
+ 1.387e+11Hz 0.0678392 0.136565
+ 1.388e+11Hz 0.0681085 0.136523
+ 1.389e+11Hz 0.0683777 0.136481
+ 1.39e+11Hz 0.068647 0.136438
+ 1.391e+11Hz 0.0689163 0.136394
+ 1.392e+11Hz 0.0691856 0.136349
+ 1.393e+11Hz 0.0694549 0.136303
+ 1.394e+11Hz 0.0697243 0.136257
+ 1.395e+11Hz 0.0699937 0.13621
+ 1.396e+11Hz 0.070263 0.136161
+ 1.397e+11Hz 0.0705324 0.136113
+ 1.398e+11Hz 0.0708018 0.136063
+ 1.399e+11Hz 0.0710712 0.136012
+ 1.4e+11Hz 0.0713406 0.135961
+ 1.401e+11Hz 0.07161 0.135908
+ 1.402e+11Hz 0.0718794 0.135855
+ 1.403e+11Hz 0.0721489 0.135801
+ 1.404e+11Hz 0.0724183 0.135747
+ 1.405e+11Hz 0.0726877 0.135691
+ 1.406e+11Hz 0.0729571 0.135634
+ 1.407e+11Hz 0.0732264 0.135577
+ 1.408e+11Hz 0.0734958 0.135519
+ 1.409e+11Hz 0.0737652 0.13546
+ 1.41e+11Hz 0.0740346 0.1354
+ 1.411e+11Hz 0.0743039 0.135339
+ 1.412e+11Hz 0.0745732 0.135278
+ 1.413e+11Hz 0.0748425 0.135215
+ 1.414e+11Hz 0.0751118 0.135152
+ 1.415e+11Hz 0.0753811 0.135088
+ 1.416e+11Hz 0.0756503 0.135023
+ 1.417e+11Hz 0.0759195 0.134957
+ 1.418e+11Hz 0.0761887 0.13489
+ 1.419e+11Hz 0.0764578 0.134823
+ 1.42e+11Hz 0.0767269 0.134754
+ 1.421e+11Hz 0.076996 0.134685
+ 1.422e+11Hz 0.077265 0.134615
+ 1.423e+11Hz 0.077534 0.134544
+ 1.424e+11Hz 0.077803 0.134472
+ 1.425e+11Hz 0.0780718 0.134399
+ 1.426e+11Hz 0.0783407 0.134325
+ 1.427e+11Hz 0.0786095 0.134251
+ 1.428e+11Hz 0.0788782 0.134175
+ 1.429e+11Hz 0.0791469 0.134099
+ 1.43e+11Hz 0.0794156 0.134022
+ 1.431e+11Hz 0.0796841 0.133944
+ 1.432e+11Hz 0.0799526 0.133865
+ 1.433e+11Hz 0.0802211 0.133785
+ 1.434e+11Hz 0.0804895 0.133705
+ 1.435e+11Hz 0.0807578 0.133623
+ 1.436e+11Hz 0.081026 0.133541
+ 1.437e+11Hz 0.0812941 0.133457
+ 1.438e+11Hz 0.0815622 0.133373
+ 1.439e+11Hz 0.0818302 0.133288
+ 1.44e+11Hz 0.0820981 0.133202
+ 1.441e+11Hz 0.0823659 0.133115
+ 1.442e+11Hz 0.0826336 0.133027
+ 1.443e+11Hz 0.0829012 0.132939
+ 1.444e+11Hz 0.0831688 0.132849
+ 1.445e+11Hz 0.0834362 0.132759
+ 1.446e+11Hz 0.0837035 0.132668
+ 1.447e+11Hz 0.0839708 0.132575
+ 1.448e+11Hz 0.0842379 0.132482
+ 1.449e+11Hz 0.0845049 0.132388
+ 1.45e+11Hz 0.0847718 0.132293
+ 1.451e+11Hz 0.0850386 0.132197
+ 1.452e+11Hz 0.0853052 0.132101
+ 1.453e+11Hz 0.0855717 0.132003
+ 1.454e+11Hz 0.0858381 0.131905
+ 1.455e+11Hz 0.0861044 0.131805
+ 1.456e+11Hz 0.0863705 0.131705
+ 1.457e+11Hz 0.0866365 0.131604
+ 1.458e+11Hz 0.0869024 0.131501
+ 1.459e+11Hz 0.0871681 0.131398
+ 1.46e+11Hz 0.0874337 0.131294
+ 1.461e+11Hz 0.0876991 0.131189
+ 1.462e+11Hz 0.0879644 0.131083
+ 1.463e+11Hz 0.0882295 0.130977
+ 1.464e+11Hz 0.0884944 0.130869
+ 1.465e+11Hz 0.0887592 0.130761
+ 1.466e+11Hz 0.0890238 0.130651
+ 1.467e+11Hz 0.0892883 0.130541
+ 1.468e+11Hz 0.0895525 0.13043
+ 1.469e+11Hz 0.0898166 0.130317
+ 1.47e+11Hz 0.0900805 0.130204
+ 1.471e+11Hz 0.0903443 0.13009
+ 1.472e+11Hz 0.0906078 0.129975
+ 1.473e+11Hz 0.0908711 0.129859
+ 1.474e+11Hz 0.0911343 0.129742
+ 1.475e+11Hz 0.0913972 0.129625
+ 1.476e+11Hz 0.09166 0.129506
+ 1.477e+11Hz 0.0919225 0.129386
+ 1.478e+11Hz 0.0921848 0.129266
+ 1.479e+11Hz 0.0924469 0.129144
+ 1.48e+11Hz 0.0927088 0.129022
+ 1.481e+11Hz 0.0929705 0.128899
+ 1.482e+11Hz 0.0932319 0.128775
+ 1.483e+11Hz 0.0934931 0.128649
+ 1.484e+11Hz 0.0937541 0.128523
+ 1.485e+11Hz 0.0940148 0.128396
+ 1.486e+11Hz 0.0942753 0.128269
+ 1.487e+11Hz 0.0945356 0.12814
+ 1.488e+11Hz 0.0947956 0.12801
+ 1.489e+11Hz 0.0950553 0.127879
+ 1.49e+11Hz 0.0953148 0.127748
+ 1.491e+11Hz 0.095574 0.127615
+ 1.492e+11Hz 0.095833 0.127482
+ 1.493e+11Hz 0.0960917 0.127348
+ 1.494e+11Hz 0.0963501 0.127212
+ 1.495e+11Hz 0.0966083 0.127076
+ 1.496e+11Hz 0.0968661 0.126939
+ 1.497e+11Hz 0.0971237 0.126801
+ 1.498e+11Hz 0.097381 0.126662
+ 1.499e+11Hz 0.097638 0.126522
+ 1.5e+11Hz 0.0978947 0.126381
+ ]

A12 %vd(20 3) %vd(12, 3) xfer2
.model xfer2 xfer R_I=true table=[
+ 0Hz 0.991964 0
+ 1e+08Hz 0.991963 -0.00133515
+ 2e+08Hz 0.991959 -0.00267028
+ 3e+08Hz 0.991952 -0.00400535
+ 4e+08Hz 0.991943 -0.00534036
+ 5e+08Hz 0.991931 -0.00667526
+ 6e+08Hz 0.991916 -0.00801005
+ 7e+08Hz 0.991899 -0.00934468
+ 8e+08Hz 0.991878 -0.0106792
+ 9e+08Hz 0.991856 -0.0120134
+ 1e+09Hz 0.99183 -0.0133475
+ 1.1e+09Hz 0.991802 -0.0146813
+ 1.2e+09Hz 0.991771 -0.0160148
+ 1.3e+09Hz 0.991738 -0.0173481
+ 1.4e+09Hz 0.991702 -0.018681
+ 1.5e+09Hz 0.991663 -0.0200136
+ 1.6e+09Hz 0.991622 -0.0213459
+ 1.7e+09Hz 0.991578 -0.0226777
+ 1.8e+09Hz 0.991531 -0.0240092
+ 1.9e+09Hz 0.991482 -0.0253402
+ 2e+09Hz 0.991431 -0.0266708
+ 2.1e+09Hz 0.991376 -0.0280009
+ 2.2e+09Hz 0.991319 -0.0293305
+ 2.3e+09Hz 0.99126 -0.0306596
+ 2.4e+09Hz 0.991198 -0.0319882
+ 2.5e+09Hz 0.991133 -0.0333162
+ 2.6e+09Hz 0.991066 -0.0346437
+ 2.7e+09Hz 0.990997 -0.0359705
+ 2.8e+09Hz 0.990925 -0.0372968
+ 2.9e+09Hz 0.99085 -0.0386224
+ 3e+09Hz 0.990773 -0.0399474
+ 3.1e+09Hz 0.990694 -0.0412717
+ 3.2e+09Hz 0.990612 -0.0425953
+ 3.3e+09Hz 0.990528 -0.0439182
+ 3.4e+09Hz 0.990441 -0.0452404
+ 3.5e+09Hz 0.990352 -0.0465618
+ 3.6e+09Hz 0.990261 -0.0478825
+ 3.7e+09Hz 0.990167 -0.0492024
+ 3.8e+09Hz 0.990071 -0.0505216
+ 3.9e+09Hz 0.989972 -0.0518399
+ 4e+09Hz 0.989871 -0.0531575
+ 4.1e+09Hz 0.989768 -0.0544742
+ 4.2e+09Hz 0.989663 -0.0557901
+ 4.3e+09Hz 0.989555 -0.0571051
+ 4.4e+09Hz 0.989446 -0.0584192
+ 4.5e+09Hz 0.989334 -0.0597325
+ 4.6e+09Hz 0.989219 -0.0610449
+ 4.7e+09Hz 0.989103 -0.0623564
+ 4.8e+09Hz 0.988984 -0.063667
+ 4.9e+09Hz 0.988864 -0.0649766
+ 5e+09Hz 0.988741 -0.0662854
+ 5.1e+09Hz 0.988616 -0.0675932
+ 5.2e+09Hz 0.988489 -0.0689001
+ 5.3e+09Hz 0.98836 -0.070206
+ 5.4e+09Hz 0.988229 -0.0715109
+ 5.5e+09Hz 0.988096 -0.0728149
+ 5.6e+09Hz 0.987961 -0.0741179
+ 5.7e+09Hz 0.987823 -0.0754199
+ 5.8e+09Hz 0.987684 -0.076721
+ 5.9e+09Hz 0.987543 -0.078021
+ 6e+09Hz 0.9874 -0.0793201
+ 6.1e+09Hz 0.987255 -0.0806182
+ 6.2e+09Hz 0.987109 -0.0819152
+ 6.3e+09Hz 0.98696 -0.0832113
+ 6.4e+09Hz 0.98681 -0.0845064
+ 6.5e+09Hz 0.986657 -0.0858004
+ 6.6e+09Hz 0.986503 -0.0870935
+ 6.7e+09Hz 0.986348 -0.0883855
+ 6.8e+09Hz 0.98619 -0.0896765
+ 6.9e+09Hz 0.986031 -0.0909665
+ 7e+09Hz 0.985869 -0.0922555
+ 7.1e+09Hz 0.985707 -0.0935435
+ 7.2e+09Hz 0.985542 -0.0948305
+ 7.3e+09Hz 0.985376 -0.0961165
+ 7.4e+09Hz 0.985208 -0.0974015
+ 7.5e+09Hz 0.985038 -0.0986855
+ 7.6e+09Hz 0.984867 -0.0999684
+ 7.7e+09Hz 0.984695 -0.10125
+ 7.8e+09Hz 0.98452 -0.102531
+ 7.9e+09Hz 0.984344 -0.103811
+ 8e+09Hz 0.984167 -0.105091
+ 8.1e+09Hz 0.983988 -0.106369
+ 8.2e+09Hz 0.983807 -0.107646
+ 8.3e+09Hz 0.983625 -0.108922
+ 8.4e+09Hz 0.983442 -0.110197
+ 8.5e+09Hz 0.983257 -0.111471
+ 8.6e+09Hz 0.98307 -0.112744
+ 8.7e+09Hz 0.982882 -0.114017
+ 8.8e+09Hz 0.982693 -0.115288
+ 8.9e+09Hz 0.982502 -0.116558
+ 9e+09Hz 0.98231 -0.117828
+ 9.1e+09Hz 0.982116 -0.119096
+ 9.2e+09Hz 0.981922 -0.120364
+ 9.3e+09Hz 0.981725 -0.121631
+ 9.4e+09Hz 0.981527 -0.122897
+ 9.5e+09Hz 0.981329 -0.124162
+ 9.6e+09Hz 0.981128 -0.125426
+ 9.7e+09Hz 0.980927 -0.12669
+ 9.8e+09Hz 0.980724 -0.127952
+ 9.9e+09Hz 0.980519 -0.129214
+ 1e+10Hz 0.980314 -0.130474
+ 1.01e+10Hz 0.980107 -0.131735
+ 1.02e+10Hz 0.979899 -0.132994
+ 1.03e+10Hz 0.979689 -0.134252
+ 1.04e+10Hz 0.979479 -0.13551
+ 1.05e+10Hz 0.979267 -0.136767
+ 1.06e+10Hz 0.979054 -0.138023
+ 1.07e+10Hz 0.97884 -0.139278
+ 1.08e+10Hz 0.978624 -0.140532
+ 1.09e+10Hz 0.978407 -0.141786
+ 1.1e+10Hz 0.97819 -0.143039
+ 1.11e+10Hz 0.97797 -0.144292
+ 1.12e+10Hz 0.97775 -0.145543
+ 1.13e+10Hz 0.977529 -0.146794
+ 1.14e+10Hz 0.977306 -0.148045
+ 1.15e+10Hz 0.977082 -0.149294
+ 1.16e+10Hz 0.976857 -0.150543
+ 1.17e+10Hz 0.976631 -0.151792
+ 1.18e+10Hz 0.976404 -0.153039
+ 1.19e+10Hz 0.976175 -0.154287
+ 1.2e+10Hz 0.975945 -0.155533
+ 1.21e+10Hz 0.975715 -0.156779
+ 1.22e+10Hz 0.975483 -0.158024
+ 1.23e+10Hz 0.975249 -0.159269
+ 1.24e+10Hz 0.975015 -0.160513
+ 1.25e+10Hz 0.97478 -0.161757
+ 1.26e+10Hz 0.974543 -0.163
+ 1.27e+10Hz 0.974306 -0.164242
+ 1.28e+10Hz 0.974067 -0.165485
+ 1.29e+10Hz 0.973827 -0.166726
+ 1.3e+10Hz 0.973586 -0.167967
+ 1.31e+10Hz 0.973343 -0.169208
+ 1.32e+10Hz 0.9731 -0.170448
+ 1.33e+10Hz 0.972855 -0.171687
+ 1.34e+10Hz 0.97261 -0.172926
+ 1.35e+10Hz 0.972363 -0.174165
+ 1.36e+10Hz 0.972115 -0.175403
+ 1.37e+10Hz 0.971866 -0.176641
+ 1.38e+10Hz 0.971615 -0.177878
+ 1.39e+10Hz 0.971364 -0.179115
+ 1.4e+10Hz 0.971111 -0.180352
+ 1.41e+10Hz 0.970857 -0.181588
+ 1.42e+10Hz 0.970603 -0.182823
+ 1.43e+10Hz 0.970346 -0.184059
+ 1.44e+10Hz 0.970089 -0.185294
+ 1.45e+10Hz 0.969831 -0.186529
+ 1.46e+10Hz 0.969571 -0.187763
+ 1.47e+10Hz 0.96931 -0.188997
+ 1.48e+10Hz 0.969048 -0.19023
+ 1.49e+10Hz 0.968785 -0.191464
+ 1.5e+10Hz 0.96852 -0.192696
+ 1.51e+10Hz 0.968255 -0.193929
+ 1.52e+10Hz 0.967988 -0.195161
+ 1.53e+10Hz 0.96772 -0.196393
+ 1.54e+10Hz 0.967451 -0.197625
+ 1.55e+10Hz 0.96718 -0.198857
+ 1.56e+10Hz 0.966908 -0.200088
+ 1.57e+10Hz 0.966635 -0.201319
+ 1.58e+10Hz 0.966361 -0.202549
+ 1.59e+10Hz 0.966086 -0.20378
+ 1.6e+10Hz 0.965809 -0.20501
+ 1.61e+10Hz 0.965531 -0.206239
+ 1.62e+10Hz 0.965252 -0.207469
+ 1.63e+10Hz 0.964971 -0.208698
+ 1.64e+10Hz 0.964689 -0.209927
+ 1.65e+10Hz 0.964406 -0.211156
+ 1.66e+10Hz 0.964122 -0.212385
+ 1.67e+10Hz 0.963836 -0.213613
+ 1.68e+10Hz 0.963549 -0.214841
+ 1.69e+10Hz 0.963261 -0.216069
+ 1.7e+10Hz 0.962971 -0.217296
+ 1.71e+10Hz 0.96268 -0.218524
+ 1.72e+10Hz 0.962388 -0.219751
+ 1.73e+10Hz 0.962094 -0.220978
+ 1.74e+10Hz 0.961799 -0.222204
+ 1.75e+10Hz 0.961503 -0.223431
+ 1.76e+10Hz 0.961205 -0.224657
+ 1.77e+10Hz 0.960906 -0.225883
+ 1.78e+10Hz 0.960606 -0.227109
+ 1.79e+10Hz 0.960304 -0.228335
+ 1.8e+10Hz 0.960001 -0.22956
+ 1.81e+10Hz 0.959696 -0.230785
+ 1.82e+10Hz 0.95939 -0.23201
+ 1.83e+10Hz 0.959082 -0.233235
+ 1.84e+10Hz 0.958773 -0.234459
+ 1.85e+10Hz 0.958463 -0.235684
+ 1.86e+10Hz 0.958151 -0.236908
+ 1.87e+10Hz 0.957838 -0.238131
+ 1.88e+10Hz 0.957524 -0.239355
+ 1.89e+10Hz 0.957207 -0.240579
+ 1.9e+10Hz 0.95689 -0.241802
+ 1.91e+10Hz 0.956571 -0.243025
+ 1.92e+10Hz 0.95625 -0.244247
+ 1.93e+10Hz 0.955928 -0.24547
+ 1.94e+10Hz 0.955605 -0.246692
+ 1.95e+10Hz 0.95528 -0.247914
+ 1.96e+10Hz 0.954953 -0.249136
+ 1.97e+10Hz 0.954625 -0.250357
+ 1.98e+10Hz 0.954296 -0.251579
+ 1.99e+10Hz 0.953965 -0.2528
+ 2e+10Hz 0.953632 -0.25402
+ 2.01e+10Hz 0.953298 -0.255241
+ 2.02e+10Hz 0.952963 -0.256461
+ 2.03e+10Hz 0.952626 -0.257681
+ 2.04e+10Hz 0.952287 -0.258901
+ 2.05e+10Hz 0.951947 -0.26012
+ 2.06e+10Hz 0.951605 -0.26134
+ 2.07e+10Hz 0.951262 -0.262558
+ 2.08e+10Hz 0.950917 -0.263777
+ 2.09e+10Hz 0.95057 -0.264995
+ 2.1e+10Hz 0.950222 -0.266213
+ 2.11e+10Hz 0.949873 -0.267431
+ 2.12e+10Hz 0.949522 -0.268649
+ 2.13e+10Hz 0.949169 -0.269866
+ 2.14e+10Hz 0.948814 -0.271082
+ 2.15e+10Hz 0.948458 -0.272299
+ 2.16e+10Hz 0.948101 -0.273515
+ 2.17e+10Hz 0.947742 -0.274731
+ 2.18e+10Hz 0.947381 -0.275946
+ 2.19e+10Hz 0.947019 -0.277161
+ 2.2e+10Hz 0.946655 -0.278376
+ 2.21e+10Hz 0.946289 -0.279591
+ 2.22e+10Hz 0.945922 -0.280805
+ 2.23e+10Hz 0.945553 -0.282018
+ 2.24e+10Hz 0.945183 -0.283232
+ 2.25e+10Hz 0.944811 -0.284445
+ 2.26e+10Hz 0.944437 -0.285657
+ 2.27e+10Hz 0.944062 -0.286869
+ 2.28e+10Hz 0.943685 -0.288081
+ 2.29e+10Hz 0.943306 -0.289293
+ 2.3e+10Hz 0.942926 -0.290504
+ 2.31e+10Hz 0.942544 -0.291714
+ 2.32e+10Hz 0.942161 -0.292924
+ 2.33e+10Hz 0.941776 -0.294134
+ 2.34e+10Hz 0.941389 -0.295343
+ 2.35e+10Hz 0.941001 -0.296552
+ 2.36e+10Hz 0.940611 -0.29776
+ 2.37e+10Hz 0.940219 -0.298969
+ 2.38e+10Hz 0.939826 -0.300176
+ 2.39e+10Hz 0.939431 -0.301383
+ 2.4e+10Hz 0.939035 -0.30259
+ 2.41e+10Hz 0.938637 -0.303796
+ 2.42e+10Hz 0.938237 -0.305001
+ 2.43e+10Hz 0.937835 -0.306206
+ 2.44e+10Hz 0.937432 -0.307411
+ 2.45e+10Hz 0.937028 -0.308615
+ 2.46e+10Hz 0.936621 -0.309819
+ 2.47e+10Hz 0.936213 -0.311022
+ 2.48e+10Hz 0.935804 -0.312225
+ 2.49e+10Hz 0.935393 -0.313427
+ 2.5e+10Hz 0.93498 -0.314629
+ 2.51e+10Hz 0.934565 -0.31583
+ 2.52e+10Hz 0.934149 -0.31703
+ 2.53e+10Hz 0.933731 -0.31823
+ 2.54e+10Hz 0.933312 -0.31943
+ 2.55e+10Hz 0.932891 -0.320629
+ 2.56e+10Hz 0.932468 -0.321827
+ 2.57e+10Hz 0.932044 -0.323025
+ 2.58e+10Hz 0.931618 -0.324222
+ 2.59e+10Hz 0.931191 -0.325419
+ 2.6e+10Hz 0.930762 -0.326615
+ 2.61e+10Hz 0.930331 -0.32781
+ 2.62e+10Hz 0.929899 -0.329005
+ 2.63e+10Hz 0.929465 -0.330199
+ 2.64e+10Hz 0.929029 -0.331393
+ 2.65e+10Hz 0.928592 -0.332586
+ 2.66e+10Hz 0.928153 -0.333779
+ 2.67e+10Hz 0.927713 -0.334971
+ 2.68e+10Hz 0.927271 -0.336162
+ 2.69e+10Hz 0.926828 -0.337353
+ 2.7e+10Hz 0.926383 -0.338543
+ 2.71e+10Hz 0.925936 -0.339732
+ 2.72e+10Hz 0.925488 -0.340921
+ 2.73e+10Hz 0.925038 -0.342109
+ 2.74e+10Hz 0.924586 -0.343297
+ 2.75e+10Hz 0.924133 -0.344484
+ 2.76e+10Hz 0.923679 -0.34567
+ 2.77e+10Hz 0.923222 -0.346856
+ 2.78e+10Hz 0.922765 -0.348041
+ 2.79e+10Hz 0.922306 -0.349225
+ 2.8e+10Hz 0.921845 -0.350409
+ 2.81e+10Hz 0.921382 -0.351592
+ 2.82e+10Hz 0.920918 -0.352774
+ 2.83e+10Hz 0.920453 -0.353955
+ 2.84e+10Hz 0.919986 -0.355137
+ 2.85e+10Hz 0.919517 -0.356317
+ 2.86e+10Hz 0.919047 -0.357496
+ 2.87e+10Hz 0.918575 -0.358675
+ 2.88e+10Hz 0.918102 -0.359854
+ 2.89e+10Hz 0.917627 -0.361031
+ 2.9e+10Hz 0.917151 -0.362208
+ 2.91e+10Hz 0.916673 -0.363384
+ 2.92e+10Hz 0.916194 -0.36456
+ 2.93e+10Hz 0.915713 -0.365735
+ 2.94e+10Hz 0.915231 -0.366909
+ 2.95e+10Hz 0.914747 -0.368082
+ 2.96e+10Hz 0.914261 -0.369255
+ 2.97e+10Hz 0.913775 -0.370427
+ 2.98e+10Hz 0.913286 -0.371598
+ 2.99e+10Hz 0.912796 -0.372769
+ 3e+10Hz 0.912305 -0.373939
+ 3.01e+10Hz 0.911812 -0.375108
+ 3.02e+10Hz 0.911318 -0.376277
+ 3.03e+10Hz 0.910822 -0.377444
+ 3.04e+10Hz 0.910325 -0.378611
+ 3.05e+10Hz 0.909826 -0.379778
+ 3.06e+10Hz 0.909326 -0.380943
+ 3.07e+10Hz 0.908824 -0.382108
+ 3.08e+10Hz 0.90832 -0.383273
+ 3.09e+10Hz 0.907816 -0.384436
+ 3.1e+10Hz 0.90731 -0.385599
+ 3.11e+10Hz 0.906802 -0.386761
+ 3.12e+10Hz 0.906293 -0.387922
+ 3.13e+10Hz 0.905783 -0.389083
+ 3.14e+10Hz 0.90527 -0.390243
+ 3.15e+10Hz 0.904757 -0.391402
+ 3.16e+10Hz 0.904242 -0.39256
+ 3.17e+10Hz 0.903726 -0.393718
+ 3.18e+10Hz 0.903208 -0.394875
+ 3.19e+10Hz 0.902689 -0.396031
+ 3.2e+10Hz 0.902168 -0.397187
+ 3.21e+10Hz 0.901646 -0.398342
+ 3.22e+10Hz 0.901123 -0.399496
+ 3.23e+10Hz 0.900598 -0.400649
+ 3.24e+10Hz 0.900072 -0.401802
+ 3.25e+10Hz 0.899544 -0.402954
+ 3.26e+10Hz 0.899015 -0.404105
+ 3.27e+10Hz 0.898484 -0.405255
+ 3.28e+10Hz 0.897952 -0.406405
+ 3.29e+10Hz 0.897418 -0.407554
+ 3.3e+10Hz 0.896883 -0.408702
+ 3.31e+10Hz 0.896347 -0.40985
+ 3.32e+10Hz 0.89581 -0.410997
+ 3.33e+10Hz 0.89527 -0.412143
+ 3.34e+10Hz 0.89473 -0.413288
+ 3.35e+10Hz 0.894188 -0.414433
+ 3.36e+10Hz 0.893645 -0.415577
+ 3.37e+10Hz 0.8931 -0.41672
+ 3.38e+10Hz 0.892554 -0.417863
+ 3.39e+10Hz 0.892006 -0.419004
+ 3.4e+10Hz 0.891457 -0.420145
+ 3.41e+10Hz 0.890907 -0.421286
+ 3.42e+10Hz 0.890355 -0.422425
+ 3.43e+10Hz 0.889802 -0.423564
+ 3.44e+10Hz 0.889248 -0.424702
+ 3.45e+10Hz 0.888692 -0.42584
+ 3.46e+10Hz 0.888134 -0.426976
+ 3.47e+10Hz 0.887576 -0.428112
+ 3.48e+10Hz 0.887016 -0.429248
+ 3.49e+10Hz 0.886454 -0.430382
+ 3.5e+10Hz 0.885891 -0.431516
+ 3.51e+10Hz 0.885327 -0.432649
+ 3.52e+10Hz 0.884761 -0.433781
+ 3.53e+10Hz 0.884194 -0.434913
+ 3.54e+10Hz 0.883626 -0.436044
+ 3.55e+10Hz 0.883056 -0.437174
+ 3.56e+10Hz 0.882485 -0.438303
+ 3.57e+10Hz 0.881912 -0.439432
+ 3.58e+10Hz 0.881339 -0.44056
+ 3.59e+10Hz 0.880763 -0.441687
+ 3.6e+10Hz 0.880186 -0.442814
+ 3.61e+10Hz 0.879608 -0.44394
+ 3.62e+10Hz 0.879029 -0.445065
+ 3.63e+10Hz 0.878448 -0.446189
+ 3.64e+10Hz 0.877866 -0.447313
+ 3.65e+10Hz 0.877282 -0.448436
+ 3.66e+10Hz 0.876697 -0.449558
+ 3.67e+10Hz 0.876111 -0.45068
+ 3.68e+10Hz 0.875523 -0.4518
+ 3.69e+10Hz 0.874934 -0.45292
+ 3.7e+10Hz 0.874343 -0.45404
+ 3.71e+10Hz 0.873751 -0.455158
+ 3.72e+10Hz 0.873158 -0.456276
+ 3.73e+10Hz 0.872563 -0.457393
+ 3.74e+10Hz 0.871967 -0.45851
+ 3.75e+10Hz 0.871369 -0.459625
+ 3.76e+10Hz 0.870771 -0.46074
+ 3.77e+10Hz 0.87017 -0.461854
+ 3.78e+10Hz 0.869569 -0.462968
+ 3.79e+10Hz 0.868966 -0.464081
+ 3.8e+10Hz 0.868361 -0.465193
+ 3.81e+10Hz 0.867755 -0.466304
+ 3.82e+10Hz 0.867148 -0.467415
+ 3.83e+10Hz 0.86654 -0.468524
+ 3.84e+10Hz 0.86593 -0.469633
+ 3.85e+10Hz 0.865318 -0.470742
+ 3.86e+10Hz 0.864705 -0.471849
+ 3.87e+10Hz 0.864091 -0.472956
+ 3.88e+10Hz 0.863476 -0.474062
+ 3.89e+10Hz 0.862859 -0.475168
+ 3.9e+10Hz 0.86224 -0.476273
+ 3.91e+10Hz 0.861621 -0.477376
+ 3.92e+10Hz 0.861 -0.47848
+ 3.93e+10Hz 0.860377 -0.479582
+ 3.94e+10Hz 0.859753 -0.480684
+ 3.95e+10Hz 0.859128 -0.481785
+ 3.96e+10Hz 0.858501 -0.482885
+ 3.97e+10Hz 0.857873 -0.483984
+ 3.98e+10Hz 0.857243 -0.485083
+ 3.99e+10Hz 0.856612 -0.486181
+ 4e+10Hz 0.85598 -0.487278
+ 4.01e+10Hz 0.855346 -0.488375
+ 4.02e+10Hz 0.854711 -0.48947
+ 4.03e+10Hz 0.854075 -0.490565
+ 4.04e+10Hz 0.853437 -0.491659
+ 4.05e+10Hz 0.852797 -0.492753
+ 4.06e+10Hz 0.852157 -0.493845
+ 4.07e+10Hz 0.851514 -0.494937
+ 4.08e+10Hz 0.850871 -0.496028
+ 4.09e+10Hz 0.850226 -0.497119
+ 4.1e+10Hz 0.84958 -0.498208
+ 4.11e+10Hz 0.848932 -0.499297
+ 4.12e+10Hz 0.848283 -0.500385
+ 4.13e+10Hz 0.847632 -0.501472
+ 4.14e+10Hz 0.84698 -0.502558
+ 4.15e+10Hz 0.846326 -0.503644
+ 4.16e+10Hz 0.845672 -0.504729
+ 4.17e+10Hz 0.845015 -0.505813
+ 4.18e+10Hz 0.844358 -0.506896
+ 4.19e+10Hz 0.843699 -0.507978
+ 4.2e+10Hz 0.843038 -0.50906
+ 4.21e+10Hz 0.842376 -0.510141
+ 4.22e+10Hz 0.841713 -0.511221
+ 4.23e+10Hz 0.841048 -0.5123
+ 4.24e+10Hz 0.840382 -0.513378
+ 4.25e+10Hz 0.839715 -0.514456
+ 4.26e+10Hz 0.839045 -0.515533
+ 4.27e+10Hz 0.838375 -0.516609
+ 4.28e+10Hz 0.837703 -0.517684
+ 4.29e+10Hz 0.83703 -0.518758
+ 4.3e+10Hz 0.836356 -0.519832
+ 4.31e+10Hz 0.835679 -0.520904
+ 4.32e+10Hz 0.835002 -0.521976
+ 4.33e+10Hz 0.834323 -0.523047
+ 4.34e+10Hz 0.833643 -0.524118
+ 4.35e+10Hz 0.832961 -0.525187
+ 4.36e+10Hz 0.832278 -0.526255
+ 4.37e+10Hz 0.831593 -0.527323
+ 4.38e+10Hz 0.830908 -0.52839
+ 4.39e+10Hz 0.83022 -0.529456
+ 4.4e+10Hz 0.829531 -0.530521
+ 4.41e+10Hz 0.828841 -0.531585
+ 4.42e+10Hz 0.82815 -0.532648
+ 4.43e+10Hz 0.827457 -0.533711
+ 4.44e+10Hz 0.826762 -0.534772
+ 4.45e+10Hz 0.826066 -0.535833
+ 4.46e+10Hz 0.825369 -0.536893
+ 4.47e+10Hz 0.82467 -0.537952
+ 4.48e+10Hz 0.82397 -0.53901
+ 4.49e+10Hz 0.823269 -0.540067
+ 4.5e+10Hz 0.822566 -0.541124
+ 4.51e+10Hz 0.821862 -0.542179
+ 4.52e+10Hz 0.821156 -0.543234
+ 4.53e+10Hz 0.820449 -0.544287
+ 4.54e+10Hz 0.81974 -0.54534
+ 4.55e+10Hz 0.81903 -0.546392
+ 4.56e+10Hz 0.818319 -0.547443
+ 4.57e+10Hz 0.817607 -0.548493
+ 4.58e+10Hz 0.816892 -0.549542
+ 4.59e+10Hz 0.816177 -0.55059
+ 4.6e+10Hz 0.81546 -0.551638
+ 4.61e+10Hz 0.814742 -0.552684
+ 4.62e+10Hz 0.814022 -0.55373
+ 4.63e+10Hz 0.813301 -0.554774
+ 4.64e+10Hz 0.812578 -0.555818
+ 4.65e+10Hz 0.811854 -0.55686
+ 4.66e+10Hz 0.811129 -0.557902
+ 4.67e+10Hz 0.810403 -0.558943
+ 4.68e+10Hz 0.809674 -0.559983
+ 4.69e+10Hz 0.808945 -0.561022
+ 4.7e+10Hz 0.808214 -0.56206
+ 4.71e+10Hz 0.807482 -0.563096
+ 4.72e+10Hz 0.806748 -0.564133
+ 4.73e+10Hz 0.806013 -0.565168
+ 4.74e+10Hz 0.805277 -0.566202
+ 4.75e+10Hz 0.804539 -0.567235
+ 4.76e+10Hz 0.8038 -0.568267
+ 4.77e+10Hz 0.80306 -0.569298
+ 4.78e+10Hz 0.802318 -0.570329
+ 4.79e+10Hz 0.801575 -0.571358
+ 4.8e+10Hz 0.80083 -0.572386
+ 4.81e+10Hz 0.800084 -0.573413
+ 4.82e+10Hz 0.799337 -0.57444
+ 4.83e+10Hz 0.798588 -0.575465
+ 4.84e+10Hz 0.797838 -0.576489
+ 4.85e+10Hz 0.797087 -0.577513
+ 4.86e+10Hz 0.796334 -0.578535
+ 4.87e+10Hz 0.79558 -0.579556
+ 4.88e+10Hz 0.794824 -0.580577
+ 4.89e+10Hz 0.794068 -0.581596
+ 4.9e+10Hz 0.793309 -0.582614
+ 4.91e+10Hz 0.79255 -0.583632
+ 4.92e+10Hz 0.791789 -0.584648
+ 4.93e+10Hz 0.791027 -0.585663
+ 4.94e+10Hz 0.790263 -0.586677
+ 4.95e+10Hz 0.789498 -0.587691
+ 4.96e+10Hz 0.788732 -0.588703
+ 4.97e+10Hz 0.787965 -0.589714
+ 4.98e+10Hz 0.787196 -0.590724
+ 4.99e+10Hz 0.786426 -0.591734
+ 5e+10Hz 0.785654 -0.592742
+ 5.01e+10Hz 0.784881 -0.593749
+ 5.02e+10Hz 0.784107 -0.594755
+ 5.03e+10Hz 0.783331 -0.59576
+ 5.04e+10Hz 0.782555 -0.596764
+ 5.05e+10Hz 0.781777 -0.597767
+ 5.06e+10Hz 0.780997 -0.598769
+ 5.07e+10Hz 0.780216 -0.59977
+ 5.08e+10Hz 0.779434 -0.600769
+ 5.09e+10Hz 0.778651 -0.601768
+ 5.1e+10Hz 0.777866 -0.602766
+ 5.11e+10Hz 0.77708 -0.603763
+ 5.12e+10Hz 0.776293 -0.604758
+ 5.13e+10Hz 0.775505 -0.605753
+ 5.14e+10Hz 0.774715 -0.606746
+ 5.15e+10Hz 0.773924 -0.607739
+ 5.16e+10Hz 0.773131 -0.60873
+ 5.17e+10Hz 0.772338 -0.60972
+ 5.18e+10Hz 0.771543 -0.61071
+ 5.19e+10Hz 0.770746 -0.611698
+ 5.2e+10Hz 0.769949 -0.612685
+ 5.21e+10Hz 0.76915 -0.613671
+ 5.22e+10Hz 0.76835 -0.614656
+ 5.23e+10Hz 0.767548 -0.61564
+ 5.24e+10Hz 0.766746 -0.616622
+ 5.25e+10Hz 0.765942 -0.617604
+ 5.26e+10Hz 0.765137 -0.618585
+ 5.27e+10Hz 0.76433 -0.619564
+ 5.28e+10Hz 0.763523 -0.620543
+ 5.29e+10Hz 0.762714 -0.62152
+ 5.3e+10Hz 0.761903 -0.622497
+ 5.31e+10Hz 0.761092 -0.623472
+ 5.32e+10Hz 0.760279 -0.624446
+ 5.33e+10Hz 0.759465 -0.625419
+ 5.34e+10Hz 0.75865 -0.626391
+ 5.35e+10Hz 0.757834 -0.627362
+ 5.36e+10Hz 0.757016 -0.628332
+ 5.37e+10Hz 0.756197 -0.6293
+ 5.38e+10Hz 0.755377 -0.630268
+ 5.39e+10Hz 0.754556 -0.631235
+ 5.4e+10Hz 0.753733 -0.6322
+ 5.41e+10Hz 0.752909 -0.633164
+ 5.42e+10Hz 0.752084 -0.634127
+ 5.43e+10Hz 0.751258 -0.63509
+ 5.44e+10Hz 0.75043 -0.636051
+ 5.45e+10Hz 0.749601 -0.637011
+ 5.46e+10Hz 0.748771 -0.637969
+ 5.47e+10Hz 0.74794 -0.638927
+ 5.48e+10Hz 0.747108 -0.639884
+ 5.49e+10Hz 0.746274 -0.640839
+ 5.5e+10Hz 0.745439 -0.641794
+ 5.51e+10Hz 0.744603 -0.642747
+ 5.52e+10Hz 0.743766 -0.643699
+ 5.53e+10Hz 0.742927 -0.64465
+ 5.54e+10Hz 0.742088 -0.6456
+ 5.55e+10Hz 0.741247 -0.646549
+ 5.56e+10Hz 0.740405 -0.647497
+ 5.57e+10Hz 0.739562 -0.648444
+ 5.58e+10Hz 0.738717 -0.649389
+ 5.59e+10Hz 0.737872 -0.650334
+ 5.6e+10Hz 0.737025 -0.651277
+ 5.61e+10Hz 0.736177 -0.652219
+ 5.62e+10Hz 0.735327 -0.65316
+ 5.63e+10Hz 0.734477 -0.6541
+ 5.64e+10Hz 0.733625 -0.655039
+ 5.65e+10Hz 0.732772 -0.655977
+ 5.66e+10Hz 0.731918 -0.656913
+ 5.67e+10Hz 0.731063 -0.657849
+ 5.68e+10Hz 0.730207 -0.658783
+ 5.69e+10Hz 0.729349 -0.659717
+ 5.7e+10Hz 0.728491 -0.660649
+ 5.71e+10Hz 0.727631 -0.66158
+ 5.72e+10Hz 0.72677 -0.66251
+ 5.73e+10Hz 0.725907 -0.663438
+ 5.74e+10Hz 0.725044 -0.664366
+ 5.75e+10Hz 0.724179 -0.665293
+ 5.76e+10Hz 0.723314 -0.666218
+ 5.77e+10Hz 0.722447 -0.667142
+ 5.78e+10Hz 0.721579 -0.668065
+ 5.79e+10Hz 0.720709 -0.668988
+ 5.8e+10Hz 0.719839 -0.669909
+ 5.81e+10Hz 0.718967 -0.670828
+ 5.82e+10Hz 0.718095 -0.671747
+ 5.83e+10Hz 0.717221 -0.672664
+ 5.84e+10Hz 0.716346 -0.673581
+ 5.85e+10Hz 0.715469 -0.674496
+ 5.86e+10Hz 0.714592 -0.67541
+ 5.87e+10Hz 0.713714 -0.676323
+ 5.88e+10Hz 0.712834 -0.677235
+ 5.89e+10Hz 0.711953 -0.678146
+ 5.9e+10Hz 0.711071 -0.679056
+ 5.91e+10Hz 0.710188 -0.679964
+ 5.92e+10Hz 0.709303 -0.680871
+ 5.93e+10Hz 0.708418 -0.681778
+ 5.94e+10Hz 0.707531 -0.682683
+ 5.95e+10Hz 0.706644 -0.683586
+ 5.96e+10Hz 0.705755 -0.684489
+ 5.97e+10Hz 0.704865 -0.685391
+ 5.98e+10Hz 0.703974 -0.686291
+ 5.99e+10Hz 0.703081 -0.687191
+ 6e+10Hz 0.702188 -0.688089
+ 6.01e+10Hz 0.701293 -0.688986
+ 6.02e+10Hz 0.700397 -0.689882
+ 6.03e+10Hz 0.6995 -0.690777
+ 6.04e+10Hz 0.698602 -0.69167
+ 6.05e+10Hz 0.697703 -0.692563
+ 6.06e+10Hz 0.696803 -0.693454
+ 6.07e+10Hz 0.695901 -0.694344
+ 6.08e+10Hz 0.694998 -0.695233
+ 6.09e+10Hz 0.694095 -0.696121
+ 6.1e+10Hz 0.69319 -0.697008
+ 6.11e+10Hz 0.692284 -0.697894
+ 6.12e+10Hz 0.691377 -0.698778
+ 6.13e+10Hz 0.690468 -0.699661
+ 6.14e+10Hz 0.689559 -0.700543
+ 6.15e+10Hz 0.688648 -0.701424
+ 6.16e+10Hz 0.687737 -0.702304
+ 6.17e+10Hz 0.686824 -0.703183
+ 6.18e+10Hz 0.68591 -0.70406
+ 6.19e+10Hz 0.684995 -0.704936
+ 6.2e+10Hz 0.684079 -0.705811
+ 6.21e+10Hz 0.683161 -0.706685
+ 6.22e+10Hz 0.682243 -0.707558
+ 6.23e+10Hz 0.681323 -0.70843
+ 6.24e+10Hz 0.680402 -0.7093
+ 6.25e+10Hz 0.679481 -0.710169
+ 6.26e+10Hz 0.678558 -0.711037
+ 6.27e+10Hz 0.677633 -0.711904
+ 6.28e+10Hz 0.676708 -0.71277
+ 6.29e+10Hz 0.675782 -0.713634
+ 6.3e+10Hz 0.674854 -0.714498
+ 6.31e+10Hz 0.673926 -0.71536
+ 6.32e+10Hz 0.672996 -0.716221
+ 6.33e+10Hz 0.672065 -0.717081
+ 6.34e+10Hz 0.671133 -0.717939
+ 6.35e+10Hz 0.6702 -0.718797
+ 6.36e+10Hz 0.669266 -0.719653
+ 6.37e+10Hz 0.668331 -0.720508
+ 6.38e+10Hz 0.667394 -0.721362
+ 6.39e+10Hz 0.666457 -0.722214
+ 6.4e+10Hz 0.665518 -0.723066
+ 6.41e+10Hz 0.664578 -0.723916
+ 6.42e+10Hz 0.663637 -0.724765
+ 6.43e+10Hz 0.662695 -0.725613
+ 6.44e+10Hz 0.661752 -0.72646
+ 6.45e+10Hz 0.660808 -0.727305
+ 6.46e+10Hz 0.659863 -0.728149
+ 6.47e+10Hz 0.658916 -0.728992
+ 6.48e+10Hz 0.657969 -0.729834
+ 6.49e+10Hz 0.65702 -0.730674
+ 6.5e+10Hz 0.65607 -0.731514
+ 6.51e+10Hz 0.655119 -0.732352
+ 6.52e+10Hz 0.654168 -0.733189
+ 6.53e+10Hz 0.653215 -0.734024
+ 6.54e+10Hz 0.65226 -0.734859
+ 6.55e+10Hz 0.651305 -0.735692
+ 6.56e+10Hz 0.650349 -0.736524
+ 6.57e+10Hz 0.649391 -0.737355
+ 6.58e+10Hz 0.648433 -0.738184
+ 6.59e+10Hz 0.647473 -0.739013
+ 6.6e+10Hz 0.646512 -0.73984
+ 6.61e+10Hz 0.64555 -0.740665
+ 6.62e+10Hz 0.644587 -0.74149
+ 6.63e+10Hz 0.643623 -0.742313
+ 6.64e+10Hz 0.642658 -0.743135
+ 6.65e+10Hz 0.641692 -0.743956
+ 6.66e+10Hz 0.640725 -0.744776
+ 6.67e+10Hz 0.639756 -0.745594
+ 6.68e+10Hz 0.638787 -0.746411
+ 6.69e+10Hz 0.637816 -0.747227
+ 6.7e+10Hz 0.636845 -0.748041
+ 6.71e+10Hz 0.635872 -0.748854
+ 6.72e+10Hz 0.634898 -0.749667
+ 6.73e+10Hz 0.633923 -0.750477
+ 6.74e+10Hz 0.632947 -0.751287
+ 6.75e+10Hz 0.63197 -0.752095
+ 6.76e+10Hz 0.630992 -0.752902
+ 6.77e+10Hz 0.630013 -0.753707
+ 6.78e+10Hz 0.629033 -0.754512
+ 6.79e+10Hz 0.628051 -0.755315
+ 6.8e+10Hz 0.627069 -0.756117
+ 6.81e+10Hz 0.626086 -0.756917
+ 6.82e+10Hz 0.625101 -0.757716
+ 6.83e+10Hz 0.624116 -0.758514
+ 6.84e+10Hz 0.623129 -0.759311
+ 6.85e+10Hz 0.622141 -0.760106
+ 6.86e+10Hz 0.621153 -0.7609
+ 6.87e+10Hz 0.620163 -0.761693
+ 6.88e+10Hz 0.619172 -0.762484
+ 6.89e+10Hz 0.61818 -0.763275
+ 6.9e+10Hz 0.617187 -0.764063
+ 6.91e+10Hz 0.616193 -0.764851
+ 6.92e+10Hz 0.615198 -0.765637
+ 6.93e+10Hz 0.614202 -0.766422
+ 6.94e+10Hz 0.613205 -0.767206
+ 6.95e+10Hz 0.612207 -0.767988
+ 6.96e+10Hz 0.611208 -0.768769
+ 6.97e+10Hz 0.610207 -0.769548
+ 6.98e+10Hz 0.609206 -0.770327
+ 6.99e+10Hz 0.608204 -0.771104
+ 7e+10Hz 0.6072 -0.77188
+ 7.01e+10Hz 0.606196 -0.772654
+ 7.02e+10Hz 0.605191 -0.773427
+ 7.03e+10Hz 0.604184 -0.774199
+ 7.04e+10Hz 0.603177 -0.774969
+ 7.05e+10Hz 0.602168 -0.775738
+ 7.06e+10Hz 0.601159 -0.776505
+ 7.07e+10Hz 0.600148 -0.777272
+ 7.08e+10Hz 0.599137 -0.778037
+ 7.09e+10Hz 0.598124 -0.7788
+ 7.1e+10Hz 0.597111 -0.779563
+ 7.11e+10Hz 0.596096 -0.780324
+ 7.12e+10Hz 0.595081 -0.781083
+ 7.13e+10Hz 0.594064 -0.781841
+ 7.14e+10Hz 0.593047 -0.782598
+ 7.15e+10Hz 0.592028 -0.783354
+ 7.16e+10Hz 0.591009 -0.784108
+ 7.17e+10Hz 0.589988 -0.784861
+ 7.18e+10Hz 0.588967 -0.785612
+ 7.19e+10Hz 0.587944 -0.786362
+ 7.2e+10Hz 0.586921 -0.787111
+ 7.21e+10Hz 0.585897 -0.787859
+ 7.22e+10Hz 0.584871 -0.788605
+ 7.23e+10Hz 0.583845 -0.789349
+ 7.24e+10Hz 0.582817 -0.790092
+ 7.25e+10Hz 0.581789 -0.790834
+ 7.26e+10Hz 0.58076 -0.791575
+ 7.27e+10Hz 0.57973 -0.792314
+ 7.28e+10Hz 0.578698 -0.793052
+ 7.29e+10Hz 0.577666 -0.793788
+ 7.3e+10Hz 0.576633 -0.794523
+ 7.31e+10Hz 0.575599 -0.795257
+ 7.32e+10Hz 0.574564 -0.795989
+ 7.33e+10Hz 0.573528 -0.79672
+ 7.34e+10Hz 0.572491 -0.797449
+ 7.35e+10Hz 0.571453 -0.798177
+ 7.36e+10Hz 0.570414 -0.798904
+ 7.37e+10Hz 0.569374 -0.799629
+ 7.38e+10Hz 0.568334 -0.800353
+ 7.39e+10Hz 0.567292 -0.801076
+ 7.4e+10Hz 0.566249 -0.801797
+ 7.41e+10Hz 0.565206 -0.802516
+ 7.42e+10Hz 0.564161 -0.803235
+ 7.43e+10Hz 0.563116 -0.803952
+ 7.44e+10Hz 0.56207 -0.804667
+ 7.45e+10Hz 0.561023 -0.805381
+ 7.46e+10Hz 0.559975 -0.806094
+ 7.47e+10Hz 0.558925 -0.806805
+ 7.48e+10Hz 0.557876 -0.807515
+ 7.49e+10Hz 0.556825 -0.808224
+ 7.5e+10Hz 0.555773 -0.808931
+ 7.51e+10Hz 0.55472 -0.809637
+ 7.52e+10Hz 0.553667 -0.810341
+ 7.53e+10Hz 0.552612 -0.811044
+ 7.54e+10Hz 0.551557 -0.811745
+ 7.55e+10Hz 0.550501 -0.812445
+ 7.56e+10Hz 0.549444 -0.813144
+ 7.57e+10Hz 0.548386 -0.813841
+ 7.58e+10Hz 0.547327 -0.814537
+ 7.59e+10Hz 0.546267 -0.815232
+ 7.6e+10Hz 0.545206 -0.815925
+ 7.61e+10Hz 0.544145 -0.816616
+ 7.62e+10Hz 0.543082 -0.817306
+ 7.63e+10Hz 0.542019 -0.817995
+ 7.64e+10Hz 0.540955 -0.818682
+ 7.65e+10Hz 0.53989 -0.819369
+ 7.66e+10Hz 0.538824 -0.820053
+ 7.67e+10Hz 0.537757 -0.820736
+ 7.68e+10Hz 0.536689 -0.821418
+ 7.69e+10Hz 0.535621 -0.822098
+ 7.7e+10Hz 0.534552 -0.822777
+ 7.71e+10Hz 0.533481 -0.823454
+ 7.72e+10Hz 0.53241 -0.82413
+ 7.73e+10Hz 0.531339 -0.824805
+ 7.74e+10Hz 0.530266 -0.825478
+ 7.75e+10Hz 0.529192 -0.82615
+ 7.76e+10Hz 0.528118 -0.82682
+ 7.77e+10Hz 0.527042 -0.827489
+ 7.78e+10Hz 0.525966 -0.828156
+ 7.79e+10Hz 0.52489 -0.828823
+ 7.8e+10Hz 0.523812 -0.829487
+ 7.81e+10Hz 0.522733 -0.83015
+ 7.82e+10Hz 0.521654 -0.830812
+ 7.83e+10Hz 0.520573 -0.831472
+ 7.84e+10Hz 0.519492 -0.832131
+ 7.85e+10Hz 0.51841 -0.832789
+ 7.86e+10Hz 0.517328 -0.833445
+ 7.87e+10Hz 0.516244 -0.834099
+ 7.88e+10Hz 0.51516 -0.834753
+ 7.89e+10Hz 0.514075 -0.835404
+ 7.9e+10Hz 0.512989 -0.836055
+ 7.91e+10Hz 0.511902 -0.836704
+ 7.92e+10Hz 0.510814 -0.837351
+ 7.93e+10Hz 0.509726 -0.837997
+ 7.94e+10Hz 0.508637 -0.838642
+ 7.95e+10Hz 0.507547 -0.839285
+ 7.96e+10Hz 0.506456 -0.839927
+ 7.97e+10Hz 0.505364 -0.840567
+ 7.98e+10Hz 0.504272 -0.841206
+ 7.99e+10Hz 0.503179 -0.841844
+ 8e+10Hz 0.502085 -0.84248
+ 8.01e+10Hz 0.50099 -0.843114
+ 8.02e+10Hz 0.499894 -0.843747
+ 8.03e+10Hz 0.498798 -0.844379
+ 8.04e+10Hz 0.497701 -0.845009
+ 8.05e+10Hz 0.496603 -0.845638
+ 8.06e+10Hz 0.495504 -0.846266
+ 8.07e+10Hz 0.494405 -0.846892
+ 8.08e+10Hz 0.493304 -0.847517
+ 8.09e+10Hz 0.492204 -0.84814
+ 8.1e+10Hz 0.491102 -0.848761
+ 8.11e+10Hz 0.489999 -0.849382
+ 8.12e+10Hz 0.488896 -0.85
+ 8.13e+10Hz 0.487792 -0.850618
+ 8.14e+10Hz 0.486687 -0.851234
+ 8.15e+10Hz 0.485581 -0.851848
+ 8.16e+10Hz 0.484475 -0.852461
+ 8.17e+10Hz 0.483368 -0.853073
+ 8.18e+10Hz 0.48226 -0.853683
+ 8.19e+10Hz 0.481151 -0.854292
+ 8.2e+10Hz 0.480041 -0.854899
+ 8.21e+10Hz 0.478931 -0.855505
+ 8.22e+10Hz 0.47782 -0.85611
+ 8.23e+10Hz 0.476708 -0.856713
+ 8.24e+10Hz 0.475596 -0.857314
+ 8.25e+10Hz 0.474483 -0.857915
+ 8.26e+10Hz 0.473369 -0.858513
+ 8.27e+10Hz 0.472254 -0.85911
+ 8.28e+10Hz 0.471138 -0.859706
+ 8.29e+10Hz 0.470022 -0.860301
+ 8.3e+10Hz 0.468905 -0.860893
+ 8.31e+10Hz 0.467788 -0.861485
+ 8.32e+10Hz 0.466669 -0.862075
+ 8.33e+10Hz 0.46555 -0.862664
+ 8.34e+10Hz 0.46443 -0.863251
+ 8.35e+10Hz 0.463309 -0.863837
+ 8.36e+10Hz 0.462188 -0.864421
+ 8.37e+10Hz 0.461066 -0.865004
+ 8.38e+10Hz 0.459943 -0.865585
+ 8.39e+10Hz 0.458819 -0.866165
+ 8.4e+10Hz 0.457695 -0.866743
+ 8.41e+10Hz 0.45657 -0.86732
+ 8.42e+10Hz 0.455444 -0.867896
+ 8.43e+10Hz 0.454317 -0.86847
+ 8.44e+10Hz 0.45319 -0.869043
+ 8.45e+10Hz 0.452062 -0.869614
+ 8.46e+10Hz 0.450933 -0.870184
+ 8.47e+10Hz 0.449804 -0.870752
+ 8.48e+10Hz 0.448674 -0.871319
+ 8.49e+10Hz 0.447543 -0.871884
+ 8.5e+10Hz 0.446411 -0.872448
+ 8.51e+10Hz 0.445279 -0.873011
+ 8.52e+10Hz 0.444146 -0.873572
+ 8.53e+10Hz 0.443012 -0.874131
+ 8.54e+10Hz 0.441877 -0.874689
+ 8.55e+10Hz 0.440742 -0.875246
+ 8.56e+10Hz 0.439606 -0.875801
+ 8.57e+10Hz 0.43847 -0.876355
+ 8.58e+10Hz 0.437332 -0.876907
+ 8.59e+10Hz 0.436194 -0.877458
+ 8.6e+10Hz 0.435056 -0.878007
+ 8.61e+10Hz 0.433916 -0.878555
+ 8.62e+10Hz 0.432776 -0.879101
+ 8.63e+10Hz 0.431635 -0.879646
+ 8.64e+10Hz 0.430493 -0.88019
+ 8.65e+10Hz 0.429351 -0.880732
+ 8.66e+10Hz 0.428208 -0.881272
+ 8.67e+10Hz 0.427065 -0.881811
+ 8.68e+10Hz 0.42592 -0.882349
+ 8.69e+10Hz 0.424775 -0.882885
+ 8.7e+10Hz 0.423629 -0.883419
+ 8.71e+10Hz 0.422483 -0.883952
+ 8.72e+10Hz 0.421336 -0.884484
+ 8.73e+10Hz 0.420188 -0.885014
+ 8.74e+10Hz 0.41904 -0.885543
+ 8.75e+10Hz 0.41789 -0.88607
+ 8.76e+10Hz 0.41674 -0.886596
+ 8.77e+10Hz 0.41559 -0.88712
+ 8.78e+10Hz 0.414439 -0.887643
+ 8.79e+10Hz 0.413287 -0.888164
+ 8.8e+10Hz 0.412134 -0.888684
+ 8.81e+10Hz 0.410981 -0.889202
+ 8.82e+10Hz 0.409827 -0.889719
+ 8.83e+10Hz 0.408672 -0.890234
+ 8.84e+10Hz 0.407517 -0.890748
+ 8.85e+10Hz 0.406361 -0.89126
+ 8.86e+10Hz 0.405204 -0.891771
+ 8.87e+10Hz 0.404047 -0.89228
+ 8.88e+10Hz 0.402889 -0.892788
+ 8.89e+10Hz 0.40173 -0.893294
+ 8.9e+10Hz 0.400571 -0.893799
+ 8.91e+10Hz 0.399411 -0.894302
+ 8.92e+10Hz 0.39825 -0.894804
+ 8.93e+10Hz 0.397089 -0.895304
+ 8.94e+10Hz 0.395927 -0.895803
+ 8.95e+10Hz 0.394764 -0.8963
+ 8.96e+10Hz 0.393601 -0.896795
+ 8.97e+10Hz 0.392437 -0.89729
+ 8.98e+10Hz 0.391272 -0.897782
+ 8.99e+10Hz 0.390107 -0.898273
+ 9e+10Hz 0.388941 -0.898763
+ 9.01e+10Hz 0.387774 -0.899251
+ 9.02e+10Hz 0.386607 -0.899738
+ 9.03e+10Hz 0.385439 -0.900223
+ 9.04e+10Hz 0.384271 -0.900706
+ 9.05e+10Hz 0.383102 -0.901188
+ 9.06e+10Hz 0.381932 -0.901669
+ 9.07e+10Hz 0.380762 -0.902148
+ 9.08e+10Hz 0.379591 -0.902625
+ 9.09e+10Hz 0.378419 -0.903101
+ 9.1e+10Hz 0.377247 -0.903575
+ 9.11e+10Hz 0.376074 -0.904048
+ 9.12e+10Hz 0.3749 -0.904519
+ 9.13e+10Hz 0.373726 -0.904989
+ 9.14e+10Hz 0.372551 -0.905457
+ 9.15e+10Hz 0.371376 -0.905924
+ 9.16e+10Hz 0.3702 -0.906389
+ 9.17e+10Hz 0.369023 -0.906852
+ 9.18e+10Hz 0.367846 -0.907315
+ 9.19e+10Hz 0.366668 -0.907775
+ 9.2e+10Hz 0.36549 -0.908234
+ 9.21e+10Hz 0.364311 -0.908691
+ 9.22e+10Hz 0.363131 -0.909147
+ 9.23e+10Hz 0.361951 -0.909601
+ 9.24e+10Hz 0.36077 -0.910054
+ 9.25e+10Hz 0.359588 -0.910505
+ 9.26e+10Hz 0.358407 -0.910955
+ 9.27e+10Hz 0.357224 -0.911403
+ 9.28e+10Hz 0.356041 -0.911849
+ 9.29e+10Hz 0.354857 -0.912294
+ 9.3e+10Hz 0.353673 -0.912737
+ 9.31e+10Hz 0.352488 -0.913179
+ 9.32e+10Hz 0.351302 -0.913619
+ 9.33e+10Hz 0.350116 -0.914058
+ 9.34e+10Hz 0.348929 -0.914495
+ 9.35e+10Hz 0.347742 -0.91493
+ 9.36e+10Hz 0.346554 -0.915364
+ 9.37e+10Hz 0.345366 -0.915796
+ 9.38e+10Hz 0.344177 -0.916227
+ 9.39e+10Hz 0.342987 -0.916656
+ 9.4e+10Hz 0.341797 -0.917084
+ 9.41e+10Hz 0.340607 -0.91751
+ 9.42e+10Hz 0.339415 -0.917934
+ 9.43e+10Hz 0.338224 -0.918357
+ 9.44e+10Hz 0.337032 -0.918779
+ 9.45e+10Hz 0.335839 -0.919198
+ 9.46e+10Hz 0.334645 -0.919616
+ 9.47e+10Hz 0.333452 -0.920033
+ 9.48e+10Hz 0.332257 -0.920448
+ 9.49e+10Hz 0.331062 -0.920861
+ 9.5e+10Hz 0.329867 -0.921273
+ 9.51e+10Hz 0.328671 -0.921683
+ 9.52e+10Hz 0.327474 -0.922092
+ 9.53e+10Hz 0.326277 -0.922499
+ 9.54e+10Hz 0.32508 -0.922904
+ 9.55e+10Hz 0.323882 -0.923308
+ 9.56e+10Hz 0.322683 -0.92371
+ 9.57e+10Hz 0.321484 -0.924111
+ 9.58e+10Hz 0.320285 -0.92451
+ 9.59e+10Hz 0.319084 -0.924907
+ 9.6e+10Hz 0.317884 -0.925303
+ 9.61e+10Hz 0.316683 -0.925697
+ 9.62e+10Hz 0.315481 -0.92609
+ 9.63e+10Hz 0.314279 -0.926481
+ 9.64e+10Hz 0.313077 -0.92687
+ 9.65e+10Hz 0.311874 -0.927258
+ 9.66e+10Hz 0.31067 -0.927644
+ 9.67e+10Hz 0.309466 -0.928029
+ 9.68e+10Hz 0.308262 -0.928412
+ 9.69e+10Hz 0.307057 -0.928793
+ 9.7e+10Hz 0.305851 -0.929173
+ 9.71e+10Hz 0.304645 -0.929551
+ 9.72e+10Hz 0.303439 -0.929928
+ 9.73e+10Hz 0.302232 -0.930303
+ 9.74e+10Hz 0.301025 -0.930677
+ 9.75e+10Hz 0.299817 -0.931048
+ 9.76e+10Hz 0.298609 -0.931419
+ 9.77e+10Hz 0.297401 -0.931787
+ 9.78e+10Hz 0.296192 -0.932154
+ 9.79e+10Hz 0.294982 -0.93252
+ 9.8e+10Hz 0.293772 -0.932883
+ 9.81e+10Hz 0.292562 -0.933246
+ 9.82e+10Hz 0.291351 -0.933606
+ 9.83e+10Hz 0.29014 -0.933965
+ 9.84e+10Hz 0.288928 -0.934322
+ 9.85e+10Hz 0.287716 -0.934678
+ 9.86e+10Hz 0.286504 -0.935033
+ 9.87e+10Hz 0.285291 -0.935385
+ 9.88e+10Hz 0.284077 -0.935736
+ 9.89e+10Hz 0.282863 -0.936085
+ 9.9e+10Hz 0.281649 -0.936433
+ 9.91e+10Hz 0.280435 -0.936779
+ 9.92e+10Hz 0.27922 -0.937124
+ 9.93e+10Hz 0.278004 -0.937467
+ 9.94e+10Hz 0.276789 -0.937808
+ 9.95e+10Hz 0.275572 -0.938148
+ 9.96e+10Hz 0.274356 -0.938486
+ 9.97e+10Hz 0.273139 -0.938822
+ 9.98e+10Hz 0.271922 -0.939157
+ 9.99e+10Hz 0.270704 -0.939491
+ 1e+11Hz 0.269486 -0.939822
+ 1.001e+11Hz 0.268267 -0.940152
+ 1.002e+11Hz 0.267048 -0.940481
+ 1.003e+11Hz 0.265829 -0.940808
+ 1.004e+11Hz 0.264609 -0.941133
+ 1.005e+11Hz 0.263389 -0.941457
+ 1.006e+11Hz 0.262169 -0.941779
+ 1.007e+11Hz 0.260948 -0.942099
+ 1.008e+11Hz 0.259727 -0.942418
+ 1.009e+11Hz 0.258506 -0.942735
+ 1.01e+11Hz 0.257284 -0.943051
+ 1.011e+11Hz 0.256062 -0.943365
+ 1.012e+11Hz 0.254839 -0.943678
+ 1.013e+11Hz 0.253617 -0.943989
+ 1.014e+11Hz 0.252393 -0.944298
+ 1.015e+11Hz 0.25117 -0.944606
+ 1.016e+11Hz 0.249946 -0.944912
+ 1.017e+11Hz 0.248722 -0.945216
+ 1.018e+11Hz 0.247497 -0.945519
+ 1.019e+11Hz 0.246272 -0.94582
+ 1.02e+11Hz 0.245047 -0.94612
+ 1.021e+11Hz 0.243821 -0.946418
+ 1.022e+11Hz 0.242595 -0.946715
+ 1.023e+11Hz 0.241369 -0.94701
+ 1.024e+11Hz 0.240142 -0.947303
+ 1.025e+11Hz 0.238916 -0.947595
+ 1.026e+11Hz 0.237688 -0.947885
+ 1.027e+11Hz 0.236461 -0.948174
+ 1.028e+11Hz 0.235233 -0.948461
+ 1.029e+11Hz 0.234005 -0.948746
+ 1.03e+11Hz 0.232776 -0.94903
+ 1.031e+11Hz 0.231547 -0.949312
+ 1.032e+11Hz 0.230318 -0.949593
+ 1.033e+11Hz 0.229089 -0.949872
+ 1.034e+11Hz 0.227859 -0.950149
+ 1.035e+11Hz 0.226629 -0.950425
+ 1.036e+11Hz 0.225399 -0.9507
+ 1.037e+11Hz 0.224168 -0.950972
+ 1.038e+11Hz 0.222937 -0.951244
+ 1.039e+11Hz 0.221706 -0.951513
+ 1.04e+11Hz 0.220474 -0.951781
+ 1.041e+11Hz 0.219242 -0.952048
+ 1.042e+11Hz 0.21801 -0.952312
+ 1.043e+11Hz 0.216778 -0.952576
+ 1.044e+11Hz 0.215545 -0.952837
+ 1.045e+11Hz 0.214312 -0.953097
+ 1.046e+11Hz 0.213079 -0.953356
+ 1.047e+11Hz 0.211845 -0.953613
+ 1.048e+11Hz 0.210611 -0.953868
+ 1.049e+11Hz 0.209377 -0.954122
+ 1.05e+11Hz 0.208143 -0.954374
+ 1.051e+11Hz 0.206908 -0.954625
+ 1.052e+11Hz 0.205673 -0.954874
+ 1.053e+11Hz 0.204438 -0.955121
+ 1.054e+11Hz 0.203202 -0.955367
+ 1.055e+11Hz 0.201966 -0.955611
+ 1.056e+11Hz 0.200731 -0.955854
+ 1.057e+11Hz 0.199494 -0.956095
+ 1.058e+11Hz 0.198258 -0.956335
+ 1.059e+11Hz 0.197021 -0.956573
+ 1.06e+11Hz 0.195783 -0.956809
+ 1.061e+11Hz 0.194546 -0.957044
+ 1.062e+11Hz 0.193308 -0.957278
+ 1.063e+11Hz 0.19207 -0.957509
+ 1.064e+11Hz 0.190832 -0.95774
+ 1.065e+11Hz 0.189594 -0.957968
+ 1.066e+11Hz 0.188355 -0.958195
+ 1.067e+11Hz 0.187116 -0.958421
+ 1.068e+11Hz 0.185877 -0.958645
+ 1.069e+11Hz 0.184637 -0.958867
+ 1.07e+11Hz 0.183397 -0.959088
+ 1.071e+11Hz 0.182157 -0.959307
+ 1.072e+11Hz 0.180917 -0.959524
+ 1.073e+11Hz 0.179676 -0.95974
+ 1.074e+11Hz 0.178435 -0.959955
+ 1.075e+11Hz 0.177195 -0.960168
+ 1.076e+11Hz 0.175953 -0.960379
+ 1.077e+11Hz 0.174712 -0.960589
+ 1.078e+11Hz 0.17347 -0.960797
+ 1.079e+11Hz 0.172228 -0.961004
+ 1.08e+11Hz 0.170985 -0.961209
+ 1.081e+11Hz 0.169743 -0.961412
+ 1.082e+11Hz 0.1685 -0.961614
+ 1.083e+11Hz 0.167257 -0.961814
+ 1.084e+11Hz 0.166014 -0.962013
+ 1.085e+11Hz 0.16477 -0.96221
+ 1.086e+11Hz 0.163526 -0.962406
+ 1.087e+11Hz 0.162282 -0.9626
+ 1.088e+11Hz 0.161038 -0.962792
+ 1.089e+11Hz 0.159794 -0.962983
+ 1.09e+11Hz 0.158549 -0.963172
+ 1.091e+11Hz 0.157304 -0.96336
+ 1.092e+11Hz 0.156059 -0.963546
+ 1.093e+11Hz 0.154813 -0.963731
+ 1.094e+11Hz 0.153568 -0.963914
+ 1.095e+11Hz 0.152322 -0.964095
+ 1.096e+11Hz 0.151076 -0.964275
+ 1.097e+11Hz 0.14983 -0.964453
+ 1.098e+11Hz 0.148583 -0.96463
+ 1.099e+11Hz 0.147336 -0.964805
+ 1.1e+11Hz 0.146089 -0.964978
+ 1.101e+11Hz 0.144842 -0.96515
+ 1.102e+11Hz 0.143595 -0.965321
+ 1.103e+11Hz 0.142347 -0.96549
+ 1.104e+11Hz 0.141099 -0.965657
+ 1.105e+11Hz 0.139851 -0.965822
+ 1.106e+11Hz 0.138602 -0.965986
+ 1.107e+11Hz 0.137354 -0.966149
+ 1.108e+11Hz 0.136105 -0.966309
+ 1.109e+11Hz 0.134856 -0.966469
+ 1.11e+11Hz 0.133607 -0.966626
+ 1.111e+11Hz 0.132357 -0.966782
+ 1.112e+11Hz 0.131108 -0.966937
+ 1.113e+11Hz 0.129858 -0.96709
+ 1.114e+11Hz 0.128608 -0.967241
+ 1.115e+11Hz 0.127358 -0.967391
+ 1.116e+11Hz 0.126107 -0.967539
+ 1.117e+11Hz 0.124856 -0.967685
+ 1.118e+11Hz 0.123606 -0.96783
+ 1.119e+11Hz 0.122355 -0.967973
+ 1.12e+11Hz 0.121103 -0.968115
+ 1.121e+11Hz 0.119852 -0.968255
+ 1.122e+11Hz 0.1186 -0.968394
+ 1.123e+11Hz 0.117348 -0.96853
+ 1.124e+11Hz 0.116096 -0.968666
+ 1.125e+11Hz 0.114844 -0.968799
+ 1.126e+11Hz 0.113591 -0.968931
+ 1.127e+11Hz 0.112339 -0.969062
+ 1.128e+11Hz 0.111086 -0.96919
+ 1.129e+11Hz 0.109833 -0.969318
+ 1.13e+11Hz 0.10858 -0.969443
+ 1.131e+11Hz 0.107327 -0.969567
+ 1.132e+11Hz 0.106073 -0.96969
+ 1.133e+11Hz 0.104819 -0.96981
+ 1.134e+11Hz 0.103566 -0.969929
+ 1.135e+11Hz 0.102311 -0.970047
+ 1.136e+11Hz 0.101057 -0.970163
+ 1.137e+11Hz 0.0998028 -0.970277
+ 1.138e+11Hz 0.0985482 -0.97039
+ 1.139e+11Hz 0.0972935 -0.970501
+ 1.14e+11Hz 0.0960386 -0.97061
+ 1.141e+11Hz 0.0947836 -0.970718
+ 1.142e+11Hz 0.0935283 -0.970824
+ 1.143e+11Hz 0.092273 -0.970928
+ 1.144e+11Hz 0.0910175 -0.971031
+ 1.145e+11Hz 0.0897618 -0.971133
+ 1.146e+11Hz 0.088506 -0.971232
+ 1.147e+11Hz 0.08725 -0.97133
+ 1.148e+11Hz 0.0859939 -0.971426
+ 1.149e+11Hz 0.0847377 -0.971521
+ 1.15e+11Hz 0.0834813 -0.971614
+ 1.151e+11Hz 0.0822248 -0.971705
+ 1.152e+11Hz 0.0809682 -0.971795
+ 1.153e+11Hz 0.0797114 -0.971883
+ 1.154e+11Hz 0.0784545 -0.97197
+ 1.155e+11Hz 0.0771975 -0.972055
+ 1.156e+11Hz 0.0759403 -0.972138
+ 1.157e+11Hz 0.074683 -0.972219
+ 1.158e+11Hz 0.0734256 -0.972299
+ 1.159e+11Hz 0.0721681 -0.972378
+ 1.16e+11Hz 0.0709105 -0.972454
+ 1.161e+11Hz 0.0696528 -0.972529
+ 1.162e+11Hz 0.068395 -0.972602
+ 1.163e+11Hz 0.0671371 -0.972674
+ 1.164e+11Hz 0.065879 -0.972744
+ 1.165e+11Hz 0.0646209 -0.972812
+ 1.166e+11Hz 0.0633627 -0.972879
+ 1.167e+11Hz 0.0621044 -0.972944
+ 1.168e+11Hz 0.060846 -0.973007
+ 1.169e+11Hz 0.0595875 -0.973069
+ 1.17e+11Hz 0.058329 -0.973129
+ 1.171e+11Hz 0.0570703 -0.973187
+ 1.172e+11Hz 0.0558116 -0.973244
+ 1.173e+11Hz 0.0545528 -0.973299
+ 1.174e+11Hz 0.053294 -0.973352
+ 1.175e+11Hz 0.0520351 -0.973404
+ 1.176e+11Hz 0.0507761 -0.973454
+ 1.177e+11Hz 0.0495171 -0.973502
+ 1.178e+11Hz 0.048258 -0.973549
+ 1.179e+11Hz 0.0469989 -0.973594
+ 1.18e+11Hz 0.0457397 -0.973637
+ 1.181e+11Hz 0.0444805 -0.973679
+ 1.182e+11Hz 0.0432212 -0.973719
+ 1.183e+11Hz 0.0419619 -0.973757
+ 1.184e+11Hz 0.0407026 -0.973794
+ 1.185e+11Hz 0.0394432 -0.973829
+ 1.186e+11Hz 0.0381838 -0.973862
+ 1.187e+11Hz 0.0369244 -0.973894
+ 1.188e+11Hz 0.035665 -0.973924
+ 1.189e+11Hz 0.0344055 -0.973952
+ 1.19e+11Hz 0.0331461 -0.973979
+ 1.191e+11Hz 0.0318866 -0.974004
+ 1.192e+11Hz 0.0306271 -0.974027
+ 1.193e+11Hz 0.0293676 -0.974049
+ 1.194e+11Hz 0.0281082 -0.974069
+ 1.195e+11Hz 0.0268487 -0.974087
+ 1.196e+11Hz 0.0255892 -0.974104
+ 1.197e+11Hz 0.0243298 -0.974118
+ 1.198e+11Hz 0.0230704 -0.974132
+ 1.199e+11Hz 0.0218109 -0.974143
+ 1.2e+11Hz 0.0205515 -0.974153
+ 1.201e+11Hz 0.0192922 -0.974162
+ 1.202e+11Hz 0.0180329 -0.974168
+ 1.203e+11Hz 0.0167736 -0.974173
+ 1.204e+11Hz 0.0155143 -0.974177
+ 1.205e+11Hz 0.0142551 -0.974178
+ 1.206e+11Hz 0.0129959 -0.974178
+ 1.207e+11Hz 0.0117368 -0.974176
+ 1.208e+11Hz 0.0104777 -0.974173
+ 1.209e+11Hz 0.00921866 -0.974168
+ 1.21e+11Hz 0.00795969 -0.974161
+ 1.211e+11Hz 0.00670079 -0.974153
+ 1.212e+11Hz 0.00544195 -0.974143
+ 1.213e+11Hz 0.00418318 -0.974131
+ 1.214e+11Hz 0.00292449 -0.974118
+ 1.215e+11Hz 0.00166586 -0.974103
+ 1.216e+11Hz 0.00040732 -0.974086
+ 1.217e+11Hz -0.000851141 -0.974068
+ 1.218e+11Hz -0.00210952 -0.974048
+ 1.219e+11Hz -0.0033678 -0.974026
+ 1.22e+11Hz -0.004626 -0.974003
+ 1.221e+11Hz -0.0058841 -0.973978
+ 1.222e+11Hz -0.0071421 -0.973951
+ 1.223e+11Hz -0.0084 -0.973923
+ 1.224e+11Hz -0.00965779 -0.973893
+ 1.225e+11Hz -0.0109155 -0.973862
+ 1.226e+11Hz -0.0121731 -0.973828
+ 1.227e+11Hz -0.0134305 -0.973794
+ 1.228e+11Hz -0.0146879 -0.973757
+ 1.229e+11Hz -0.0159451 -0.973719
+ 1.23e+11Hz -0.0172022 -0.97368
+ 1.231e+11Hz -0.0184592 -0.973638
+ 1.232e+11Hz -0.019716 -0.973595
+ 1.233e+11Hz -0.0209727 -0.97355
+ 1.234e+11Hz -0.0222293 -0.973504
+ 1.235e+11Hz -0.0234857 -0.973456
+ 1.236e+11Hz -0.0247421 -0.973407
+ 1.237e+11Hz -0.0259982 -0.973356
+ 1.238e+11Hz -0.0272542 -0.973303
+ 1.239e+11Hz -0.0285101 -0.973248
+ 1.24e+11Hz -0.0297658 -0.973193
+ 1.241e+11Hz -0.0310214 -0.973135
+ 1.242e+11Hz -0.0322768 -0.973076
+ 1.243e+11Hz -0.0335321 -0.973015
+ 1.244e+11Hz -0.0347872 -0.972952
+ 1.245e+11Hz -0.0360421 -0.972888
+ 1.246e+11Hz -0.0372969 -0.972823
+ 1.247e+11Hz -0.0385515 -0.972755
+ 1.248e+11Hz -0.0398059 -0.972686
+ 1.249e+11Hz -0.0410601 -0.972616
+ 1.25e+11Hz -0.0423142 -0.972544
+ 1.251e+11Hz -0.0435682 -0.97247
+ 1.252e+11Hz -0.0448219 -0.972395
+ 1.253e+11Hz -0.0460755 -0.972318
+ 1.254e+11Hz -0.0473288 -0.972239
+ 1.255e+11Hz -0.048582 -0.972159
+ 1.256e+11Hz -0.049835 -0.972078
+ 1.257e+11Hz -0.0510879 -0.971994
+ 1.258e+11Hz -0.0523405 -0.971909
+ 1.259e+11Hz -0.053593 -0.971823
+ 1.26e+11Hz -0.0548452 -0.971735
+ 1.261e+11Hz -0.0560973 -0.971646
+ 1.262e+11Hz -0.0573492 -0.971554
+ 1.263e+11Hz -0.0586009 -0.971462
+ 1.264e+11Hz -0.0598524 -0.971367
+ 1.265e+11Hz -0.0611037 -0.971272
+ 1.266e+11Hz -0.0623548 -0.971174
+ 1.267e+11Hz -0.0636057 -0.971075
+ 1.268e+11Hz -0.0648564 -0.970975
+ 1.269e+11Hz -0.0661069 -0.970873
+ 1.27e+11Hz -0.0673572 -0.970769
+ 1.271e+11Hz -0.0686072 -0.970664
+ 1.272e+11Hz -0.0698571 -0.970557
+ 1.273e+11Hz -0.0711068 -0.970449
+ 1.274e+11Hz -0.0723563 -0.970339
+ 1.275e+11Hz -0.0736056 -0.970227
+ 1.276e+11Hz -0.0748546 -0.970114
+ 1.277e+11Hz -0.0761035 -0.97
+ 1.278e+11Hz -0.0773522 -0.969884
+ 1.279e+11Hz -0.0786006 -0.969766
+ 1.28e+11Hz -0.0798488 -0.969647
+ 1.281e+11Hz -0.0810969 -0.969526
+ 1.282e+11Hz -0.0823447 -0.969404
+ 1.283e+11Hz -0.0835923 -0.96928
+ 1.284e+11Hz -0.0848397 -0.969155
+ 1.285e+11Hz -0.0860869 -0.969028
+ 1.286e+11Hz -0.0873339 -0.9689
+ 1.287e+11Hz -0.0885806 -0.96877
+ 1.288e+11Hz -0.0898272 -0.968638
+ 1.289e+11Hz -0.0910735 -0.968505
+ 1.29e+11Hz -0.0923197 -0.968371
+ 1.291e+11Hz -0.0935656 -0.968235
+ 1.292e+11Hz -0.0948113 -0.968097
+ 1.293e+11Hz -0.0960568 -0.967958
+ 1.294e+11Hz -0.0973021 -0.967817
+ 1.295e+11Hz -0.0985472 -0.967675
+ 1.296e+11Hz -0.0997921 -0.967532
+ 1.297e+11Hz -0.101037 -0.967387
+ 1.298e+11Hz -0.102281 -0.96724
+ 1.299e+11Hz -0.103526 -0.967092
+ 1.3e+11Hz -0.10477 -0.966942
+ 1.301e+11Hz -0.106013 -0.966791
+ 1.302e+11Hz -0.107257 -0.966638
+ 1.303e+11Hz -0.1085 -0.966484
+ 1.304e+11Hz -0.109744 -0.966328
+ 1.305e+11Hz -0.110987 -0.966171
+ 1.306e+11Hz -0.112229 -0.966012
+ 1.307e+11Hz -0.113472 -0.965852
+ 1.308e+11Hz -0.114714 -0.96569
+ 1.309e+11Hz -0.115957 -0.965527
+ 1.31e+11Hz -0.117198 -0.965362
+ 1.311e+11Hz -0.11844 -0.965196
+ 1.312e+11Hz -0.119682 -0.965028
+ 1.313e+11Hz -0.120923 -0.964858
+ 1.314e+11Hz -0.122164 -0.964688
+ 1.315e+11Hz -0.123405 -0.964515
+ 1.316e+11Hz -0.124646 -0.964341
+ 1.317e+11Hz -0.125887 -0.964166
+ 1.318e+11Hz -0.127127 -0.963989
+ 1.319e+11Hz -0.128367 -0.96381
+ 1.32e+11Hz -0.129607 -0.96363
+ 1.321e+11Hz -0.130847 -0.963449
+ 1.322e+11Hz -0.132086 -0.963266
+ 1.323e+11Hz -0.133326 -0.963082
+ 1.324e+11Hz -0.134565 -0.962895
+ 1.325e+11Hz -0.135804 -0.962708
+ 1.326e+11Hz -0.137043 -0.962519
+ 1.327e+11Hz -0.138281 -0.962328
+ 1.328e+11Hz -0.139519 -0.962136
+ 1.329e+11Hz -0.140758 -0.961943
+ 1.33e+11Hz -0.141996 -0.961747
+ 1.331e+11Hz -0.143233 -0.961551
+ 1.332e+11Hz -0.144471 -0.961353
+ 1.333e+11Hz -0.145708 -0.961153
+ 1.334e+11Hz -0.146946 -0.960951
+ 1.335e+11Hz -0.148182 -0.960749
+ 1.336e+11Hz -0.149419 -0.960544
+ 1.337e+11Hz -0.150656 -0.960339
+ 1.338e+11Hz -0.151892 -0.960131
+ 1.339e+11Hz -0.153128 -0.959922
+ 1.34e+11Hz -0.154364 -0.959712
+ 1.341e+11Hz -0.1556 -0.9595
+ 1.342e+11Hz -0.156836 -0.959286
+ 1.343e+11Hz -0.158071 -0.959071
+ 1.344e+11Hz -0.159306 -0.958855
+ 1.345e+11Hz -0.160541 -0.958636
+ 1.346e+11Hz -0.161776 -0.958417
+ 1.347e+11Hz -0.163011 -0.958195
+ 1.348e+11Hz -0.164245 -0.957973
+ 1.349e+11Hz -0.165479 -0.957748
+ 1.35e+11Hz -0.166713 -0.957522
+ 1.351e+11Hz -0.167947 -0.957295
+ 1.352e+11Hz -0.169181 -0.957066
+ 1.353e+11Hz -0.170414 -0.956835
+ 1.354e+11Hz -0.171647 -0.956603
+ 1.355e+11Hz -0.17288 -0.956369
+ 1.356e+11Hz -0.174113 -0.956134
+ 1.357e+11Hz -0.175346 -0.955897
+ 1.358e+11Hz -0.176578 -0.955658
+ 1.359e+11Hz -0.17781 -0.955418
+ 1.36e+11Hz -0.179042 -0.955176
+ 1.361e+11Hz -0.180274 -0.954933
+ 1.362e+11Hz -0.181505 -0.954688
+ 1.363e+11Hz -0.182737 -0.954442
+ 1.364e+11Hz -0.183968 -0.954194
+ 1.365e+11Hz -0.185198 -0.953944
+ 1.366e+11Hz -0.186429 -0.953693
+ 1.367e+11Hz -0.187659 -0.95344
+ 1.368e+11Hz -0.18889 -0.953186
+ 1.369e+11Hz -0.190119 -0.95293
+ 1.37e+11Hz -0.191349 -0.952672
+ 1.371e+11Hz -0.192579 -0.952413
+ 1.372e+11Hz -0.193808 -0.952152
+ 1.373e+11Hz -0.195037 -0.951889
+ 1.374e+11Hz -0.196266 -0.951625
+ 1.375e+11Hz -0.197494 -0.951359
+ 1.376e+11Hz -0.198722 -0.951092
+ 1.377e+11Hz -0.19995 -0.950823
+ 1.378e+11Hz -0.201178 -0.950552
+ 1.379e+11Hz -0.202405 -0.95028
+ 1.38e+11Hz -0.203633 -0.950006
+ 1.381e+11Hz -0.20486 -0.949731
+ 1.382e+11Hz -0.206086 -0.949453
+ 1.383e+11Hz -0.207313 -0.949175
+ 1.384e+11Hz -0.208539 -0.948894
+ 1.385e+11Hz -0.209765 -0.948612
+ 1.386e+11Hz -0.21099 -0.948328
+ 1.387e+11Hz -0.212216 -0.948043
+ 1.388e+11Hz -0.213441 -0.947756
+ 1.389e+11Hz -0.214665 -0.947467
+ 1.39e+11Hz -0.21589 -0.947176
+ 1.391e+11Hz -0.217114 -0.946884
+ 1.392e+11Hz -0.218338 -0.946591
+ 1.393e+11Hz -0.219561 -0.946295
+ 1.394e+11Hz -0.220784 -0.945998
+ 1.395e+11Hz -0.222007 -0.945699
+ 1.396e+11Hz -0.22323 -0.945399
+ 1.397e+11Hz -0.224452 -0.945097
+ 1.398e+11Hz -0.225674 -0.944793
+ 1.399e+11Hz -0.226895 -0.944488
+ 1.4e+11Hz -0.228116 -0.94418
+ 1.401e+11Hz -0.229337 -0.943872
+ 1.402e+11Hz -0.230558 -0.943561
+ 1.403e+11Hz -0.231778 -0.943249
+ 1.404e+11Hz -0.232998 -0.942935
+ 1.405e+11Hz -0.234217 -0.94262
+ 1.406e+11Hz -0.235436 -0.942302
+ 1.407e+11Hz -0.236655 -0.941983
+ 1.408e+11Hz -0.237873 -0.941663
+ 1.409e+11Hz -0.239091 -0.94134
+ 1.41e+11Hz -0.240309 -0.941016
+ 1.411e+11Hz -0.241526 -0.940691
+ 1.412e+11Hz -0.242742 -0.940363
+ 1.413e+11Hz -0.243958 -0.940034
+ 1.414e+11Hz -0.245174 -0.939703
+ 1.415e+11Hz -0.24639 -0.939371
+ 1.416e+11Hz -0.247605 -0.939037
+ 1.417e+11Hz -0.248819 -0.938701
+ 1.418e+11Hz -0.250034 -0.938363
+ 1.419e+11Hz -0.251247 -0.938024
+ 1.42e+11Hz -0.25246 -0.937683
+ 1.421e+11Hz -0.253673 -0.937341
+ 1.422e+11Hz -0.254885 -0.936996
+ 1.423e+11Hz -0.256097 -0.93665
+ 1.424e+11Hz -0.257309 -0.936303
+ 1.425e+11Hz -0.25852 -0.935953
+ 1.426e+11Hz -0.25973 -0.935602
+ 1.427e+11Hz -0.26094 -0.935249
+ 1.428e+11Hz -0.262149 -0.934895
+ 1.429e+11Hz -0.263358 -0.934539
+ 1.43e+11Hz -0.264567 -0.934181
+ 1.431e+11Hz -0.265775 -0.933821
+ 1.432e+11Hz -0.266982 -0.93346
+ 1.433e+11Hz -0.268189 -0.933097
+ 1.434e+11Hz -0.269395 -0.932733
+ 1.435e+11Hz -0.270601 -0.932366
+ 1.436e+11Hz -0.271806 -0.931998
+ 1.437e+11Hz -0.273011 -0.931629
+ 1.438e+11Hz -0.274215 -0.931258
+ 1.439e+11Hz -0.275418 -0.930885
+ 1.44e+11Hz -0.276621 -0.93051
+ 1.441e+11Hz -0.277824 -0.930134
+ 1.442e+11Hz -0.279026 -0.929756
+ 1.443e+11Hz -0.280227 -0.929377
+ 1.444e+11Hz -0.281428 -0.928995
+ 1.445e+11Hz -0.282628 -0.928613
+ 1.446e+11Hz -0.283827 -0.928228
+ 1.447e+11Hz -0.285026 -0.927842
+ 1.448e+11Hz -0.286224 -0.927454
+ 1.449e+11Hz -0.287422 -0.927065
+ 1.45e+11Hz -0.288619 -0.926674
+ 1.451e+11Hz -0.289815 -0.926281
+ 1.452e+11Hz -0.291011 -0.925887
+ 1.453e+11Hz -0.292206 -0.925491
+ 1.454e+11Hz -0.293401 -0.925094
+ 1.455e+11Hz -0.294594 -0.924695
+ 1.456e+11Hz -0.295788 -0.924294
+ 1.457e+11Hz -0.29698 -0.923892
+ 1.458e+11Hz -0.298172 -0.923488
+ 1.459e+11Hz -0.299363 -0.923082
+ 1.46e+11Hz -0.300554 -0.922675
+ 1.461e+11Hz -0.301744 -0.922267
+ 1.462e+11Hz -0.302933 -0.921856
+ 1.463e+11Hz -0.304121 -0.921445
+ 1.464e+11Hz -0.305309 -0.921031
+ 1.465e+11Hz -0.306496 -0.920616
+ 1.466e+11Hz -0.307683 -0.9202
+ 1.467e+11Hz -0.308868 -0.919782
+ 1.468e+11Hz -0.310054 -0.919362
+ 1.469e+11Hz -0.311238 -0.918941
+ 1.47e+11Hz -0.312422 -0.918519
+ 1.471e+11Hz -0.313605 -0.918095
+ 1.472e+11Hz -0.314787 -0.917669
+ 1.473e+11Hz -0.315968 -0.917242
+ 1.474e+11Hz -0.317149 -0.916813
+ 1.475e+11Hz -0.318329 -0.916383
+ 1.476e+11Hz -0.319509 -0.915952
+ 1.477e+11Hz -0.320688 -0.915519
+ 1.478e+11Hz -0.321865 -0.915084
+ 1.479e+11Hz -0.323043 -0.914648
+ 1.48e+11Hz -0.324219 -0.91421
+ 1.481e+11Hz -0.325395 -0.913771
+ 1.482e+11Hz -0.32657 -0.913331
+ 1.483e+11Hz -0.327744 -0.912889
+ 1.484e+11Hz -0.328918 -0.912446
+ 1.485e+11Hz -0.330091 -0.912001
+ 1.486e+11Hz -0.331263 -0.911555
+ 1.487e+11Hz -0.332435 -0.911107
+ 1.488e+11Hz -0.333605 -0.910658
+ 1.489e+11Hz -0.334775 -0.910207
+ 1.49e+11Hz -0.335944 -0.909755
+ 1.491e+11Hz -0.337113 -0.909302
+ 1.492e+11Hz -0.338281 -0.908848
+ 1.493e+11Hz -0.339448 -0.908391
+ 1.494e+11Hz -0.340614 -0.907934
+ 1.495e+11Hz -0.34178 -0.907475
+ 1.496e+11Hz -0.342945 -0.907015
+ 1.497e+11Hz -0.344109 -0.906553
+ 1.498e+11Hz -0.345272 -0.906091
+ 1.499e+11Hz -0.346435 -0.905626
+ 1.5e+11Hz -0.347597 -0.905161
+ ]

A21 %vd(10 3) %vd(21, 22) xfer3
.model xfer3 xfer R_I=true table=[
+ 0Hz 0.992005 0
+ 1e+08Hz 0.992004 -0.00131293
+ 2e+08Hz 0.992 -0.00262583
+ 3e+08Hz 0.991993 -0.00393869
+ 4e+08Hz 0.991984 -0.00525147
+ 5e+08Hz 0.991972 -0.00656415
+ 6e+08Hz 0.991958 -0.0078767
+ 7e+08Hz 0.991941 -0.00918911
+ 8e+08Hz 0.991921 -0.0105013
+ 9e+08Hz 0.991899 -0.0118134
+ 1e+09Hz 0.991874 -0.0131252
+ 1.1e+09Hz 0.991846 -0.0144368
+ 1.2e+09Hz 0.991816 -0.0157481
+ 1.3e+09Hz 0.991784 -0.0170591
+ 1.4e+09Hz 0.991748 -0.0183698
+ 1.5e+09Hz 0.991711 -0.0196802
+ 1.6e+09Hz 0.99167 -0.0209902
+ 1.7e+09Hz 0.991627 -0.0222998
+ 1.8e+09Hz 0.991582 -0.023609
+ 1.9e+09Hz 0.991534 -0.0249178
+ 2e+09Hz 0.991483 -0.0262261
+ 2.1e+09Hz 0.99143 -0.027534
+ 2.2e+09Hz 0.991374 -0.0288414
+ 2.3e+09Hz 0.991316 -0.0301482
+ 2.4e+09Hz 0.991256 -0.0314545
+ 2.5e+09Hz 0.991193 -0.0327603
+ 2.6e+09Hz 0.991127 -0.0340654
+ 2.7e+09Hz 0.991059 -0.03537
+ 2.8e+09Hz 0.990989 -0.036674
+ 2.9e+09Hz 0.990916 -0.0379773
+ 3e+09Hz 0.990841 -0.03928
+ 3.1e+09Hz 0.990763 -0.040582
+ 3.2e+09Hz 0.990683 -0.0418833
+ 3.3e+09Hz 0.990601 -0.043184
+ 3.4e+09Hz 0.990516 -0.0444839
+ 3.5e+09Hz 0.990429 -0.045783
+ 3.6e+09Hz 0.99034 -0.0470814
+ 3.7e+09Hz 0.990249 -0.048379
+ 3.8e+09Hz 0.990155 -0.0496759
+ 3.9e+09Hz 0.990059 -0.050972
+ 4e+09Hz 0.989961 -0.0522672
+ 4.1e+09Hz 0.98986 -0.0535616
+ 4.2e+09Hz 0.989757 -0.0548552
+ 4.3e+09Hz 0.989652 -0.0561479
+ 4.4e+09Hz 0.989545 -0.0574397
+ 4.5e+09Hz 0.989436 -0.0587307
+ 4.6e+09Hz 0.989325 -0.0600208
+ 4.7e+09Hz 0.989211 -0.06131
+ 4.8e+09Hz 0.989096 -0.0625983
+ 4.9e+09Hz 0.988978 -0.0638857
+ 5e+09Hz 0.988858 -0.0651721
+ 5.1e+09Hz 0.988737 -0.0664576
+ 5.2e+09Hz 0.988613 -0.0677422
+ 5.3e+09Hz 0.988487 -0.0690258
+ 5.4e+09Hz 0.98836 -0.0703084
+ 5.5e+09Hz 0.98823 -0.0715902
+ 5.6e+09Hz 0.988099 -0.0728709
+ 5.7e+09Hz 0.987965 -0.0741506
+ 5.8e+09Hz 0.98783 -0.0754294
+ 5.9e+09Hz 0.987693 -0.0767072
+ 6e+09Hz 0.987554 -0.077984
+ 6.1e+09Hz 0.987413 -0.0792599
+ 6.2e+09Hz 0.98727 -0.0805347
+ 6.3e+09Hz 0.987126 -0.0818085
+ 6.4e+09Hz 0.986979 -0.0830813
+ 6.5e+09Hz 0.986831 -0.0843532
+ 6.6e+09Hz 0.986682 -0.085624
+ 6.7e+09Hz 0.98653 -0.0868939
+ 6.8e+09Hz 0.986377 -0.0881627
+ 6.9e+09Hz 0.986222 -0.0894306
+ 7e+09Hz 0.986066 -0.0906974
+ 7.1e+09Hz 0.985908 -0.0919633
+ 7.2e+09Hz 0.985748 -0.0932281
+ 7.3e+09Hz 0.985587 -0.094492
+ 7.4e+09Hz 0.985424 -0.0957549
+ 7.5e+09Hz 0.985259 -0.0970168
+ 7.6e+09Hz 0.985093 -0.0982777
+ 7.7e+09Hz 0.984926 -0.0995376
+ 7.8e+09Hz 0.984757 -0.100797
+ 7.9e+09Hz 0.984586 -0.102055
+ 8e+09Hz 0.984414 -0.103312
+ 8.1e+09Hz 0.984241 -0.104568
+ 8.2e+09Hz 0.984066 -0.105823
+ 8.3e+09Hz 0.98389 -0.107077
+ 8.4e+09Hz 0.983712 -0.10833
+ 8.5e+09Hz 0.983533 -0.109582
+ 8.6e+09Hz 0.983352 -0.110834
+ 8.7e+09Hz 0.98317 -0.112084
+ 8.8e+09Hz 0.982987 -0.113334
+ 8.9e+09Hz 0.982802 -0.114583
+ 9e+09Hz 0.982616 -0.11583
+ 9.1e+09Hz 0.982429 -0.117077
+ 9.2e+09Hz 0.982241 -0.118323
+ 9.3e+09Hz 0.982051 -0.119568
+ 9.4e+09Hz 0.98186 -0.120813
+ 9.5e+09Hz 0.981667 -0.122056
+ 9.6e+09Hz 0.981473 -0.123299
+ 9.7e+09Hz 0.981279 -0.12454
+ 9.8e+09Hz 0.981082 -0.125781
+ 9.9e+09Hz 0.980885 -0.127021
+ 1e+10Hz 0.980687 -0.128261
+ 1.01e+10Hz 0.980487 -0.129499
+ 1.02e+10Hz 0.980286 -0.130737
+ 1.03e+10Hz 0.980084 -0.131974
+ 1.04e+10Hz 0.97988 -0.13321
+ 1.05e+10Hz 0.979676 -0.134446
+ 1.06e+10Hz 0.97947 -0.135681
+ 1.07e+10Hz 0.979263 -0.136915
+ 1.08e+10Hz 0.979055 -0.138148
+ 1.09e+10Hz 0.978846 -0.139381
+ 1.1e+10Hz 0.978636 -0.140613
+ 1.11e+10Hz 0.978425 -0.141844
+ 1.12e+10Hz 0.978212 -0.143075
+ 1.13e+10Hz 0.977999 -0.144305
+ 1.14e+10Hz 0.977784 -0.145534
+ 1.15e+10Hz 0.977568 -0.146763
+ 1.16e+10Hz 0.977351 -0.147991
+ 1.17e+10Hz 0.977133 -0.149218
+ 1.18e+10Hz 0.976914 -0.150445
+ 1.19e+10Hz 0.976694 -0.151671
+ 1.2e+10Hz 0.976472 -0.152897
+ 1.21e+10Hz 0.97625 -0.154122
+ 1.22e+10Hz 0.976027 -0.155347
+ 1.23e+10Hz 0.975802 -0.156571
+ 1.24e+10Hz 0.975576 -0.157795
+ 1.25e+10Hz 0.975349 -0.159018
+ 1.26e+10Hz 0.975122 -0.160241
+ 1.27e+10Hz 0.974893 -0.161463
+ 1.28e+10Hz 0.974663 -0.162684
+ 1.29e+10Hz 0.974432 -0.163905
+ 1.3e+10Hz 0.974199 -0.165126
+ 1.31e+10Hz 0.973966 -0.166346
+ 1.32e+10Hz 0.973732 -0.167566
+ 1.33e+10Hz 0.973496 -0.168786
+ 1.34e+10Hz 0.97326 -0.170005
+ 1.35e+10Hz 0.973022 -0.171223
+ 1.36e+10Hz 0.972783 -0.172441
+ 1.37e+10Hz 0.972543 -0.173659
+ 1.38e+10Hz 0.972302 -0.174876
+ 1.39e+10Hz 0.97206 -0.176093
+ 1.4e+10Hz 0.971817 -0.17731
+ 1.41e+10Hz 0.971573 -0.178526
+ 1.42e+10Hz 0.971328 -0.179742
+ 1.43e+10Hz 0.971081 -0.180958
+ 1.44e+10Hz 0.970833 -0.182173
+ 1.45e+10Hz 0.970585 -0.183388
+ 1.46e+10Hz 0.970335 -0.184603
+ 1.47e+10Hz 0.970084 -0.185817
+ 1.48e+10Hz 0.969831 -0.187031
+ 1.49e+10Hz 0.969578 -0.188245
+ 1.5e+10Hz 0.969324 -0.189459
+ 1.51e+10Hz 0.969068 -0.190672
+ 1.52e+10Hz 0.968811 -0.191885
+ 1.53e+10Hz 0.968553 -0.193098
+ 1.54e+10Hz 0.968294 -0.19431
+ 1.55e+10Hz 0.968034 -0.195522
+ 1.56e+10Hz 0.967772 -0.196734
+ 1.57e+10Hz 0.967509 -0.197946
+ 1.58e+10Hz 0.967245 -0.199157
+ 1.59e+10Hz 0.96698 -0.200369
+ 1.6e+10Hz 0.966714 -0.201579
+ 1.61e+10Hz 0.966446 -0.20279
+ 1.62e+10Hz 0.966177 -0.204001
+ 1.63e+10Hz 0.965907 -0.205211
+ 1.64e+10Hz 0.965636 -0.206421
+ 1.65e+10Hz 0.965363 -0.207631
+ 1.66e+10Hz 0.96509 -0.208841
+ 1.67e+10Hz 0.964815 -0.210051
+ 1.68e+10Hz 0.964538 -0.21126
+ 1.69e+10Hz 0.96426 -0.212469
+ 1.7e+10Hz 0.963982 -0.213678
+ 1.71e+10Hz 0.963701 -0.214887
+ 1.72e+10Hz 0.96342 -0.216095
+ 1.73e+10Hz 0.963137 -0.217304
+ 1.74e+10Hz 0.962853 -0.218512
+ 1.75e+10Hz 0.962567 -0.21972
+ 1.76e+10Hz 0.96228 -0.220927
+ 1.77e+10Hz 0.961992 -0.222135
+ 1.78e+10Hz 0.961703 -0.223343
+ 1.79e+10Hz 0.961412 -0.22455
+ 1.8e+10Hz 0.96112 -0.225757
+ 1.81e+10Hz 0.960826 -0.226964
+ 1.82e+10Hz 0.960531 -0.22817
+ 1.83e+10Hz 0.960235 -0.229377
+ 1.84e+10Hz 0.959937 -0.230583
+ 1.85e+10Hz 0.959638 -0.231789
+ 1.86e+10Hz 0.959337 -0.232995
+ 1.87e+10Hz 0.959035 -0.234201
+ 1.88e+10Hz 0.958732 -0.235406
+ 1.89e+10Hz 0.958427 -0.236612
+ 1.9e+10Hz 0.958121 -0.237817
+ 1.91e+10Hz 0.957813 -0.239022
+ 1.92e+10Hz 0.957504 -0.240227
+ 1.93e+10Hz 0.957193 -0.241431
+ 1.94e+10Hz 0.956881 -0.242635
+ 1.95e+10Hz 0.956568 -0.243839
+ 1.96e+10Hz 0.956253 -0.245043
+ 1.97e+10Hz 0.955936 -0.246247
+ 1.98e+10Hz 0.955619 -0.24745
+ 1.99e+10Hz 0.955299 -0.248653
+ 2e+10Hz 0.954978 -0.249856
+ 2.01e+10Hz 0.954656 -0.251059
+ 2.02e+10Hz 0.954332 -0.252262
+ 2.03e+10Hz 0.954007 -0.253464
+ 2.04e+10Hz 0.95368 -0.254666
+ 2.05e+10Hz 0.953351 -0.255867
+ 2.06e+10Hz 0.953021 -0.257069
+ 2.07e+10Hz 0.95269 -0.25827
+ 2.08e+10Hz 0.952357 -0.259471
+ 2.09e+10Hz 0.952022 -0.260672
+ 2.1e+10Hz 0.951686 -0.261872
+ 2.11e+10Hz 0.951349 -0.263072
+ 2.12e+10Hz 0.95101 -0.264272
+ 2.13e+10Hz 0.950669 -0.265471
+ 2.14e+10Hz 0.950327 -0.26667
+ 2.15e+10Hz 0.949983 -0.267869
+ 2.16e+10Hz 0.949637 -0.269068
+ 2.17e+10Hz 0.949291 -0.270266
+ 2.18e+10Hz 0.948942 -0.271464
+ 2.19e+10Hz 0.948592 -0.272662
+ 2.2e+10Hz 0.94824 -0.273859
+ 2.21e+10Hz 0.947887 -0.275056
+ 2.22e+10Hz 0.947532 -0.276253
+ 2.23e+10Hz 0.947176 -0.277449
+ 2.24e+10Hz 0.946818 -0.278645
+ 2.25e+10Hz 0.946459 -0.27984
+ 2.26e+10Hz 0.946098 -0.281035
+ 2.27e+10Hz 0.945735 -0.28223
+ 2.28e+10Hz 0.945371 -0.283424
+ 2.29e+10Hz 0.945005 -0.284618
+ 2.3e+10Hz 0.944637 -0.285812
+ 2.31e+10Hz 0.944268 -0.287005
+ 2.32e+10Hz 0.943898 -0.288198
+ 2.33e+10Hz 0.943525 -0.28939
+ 2.34e+10Hz 0.943152 -0.290582
+ 2.35e+10Hz 0.942776 -0.291774
+ 2.36e+10Hz 0.942399 -0.292965
+ 2.37e+10Hz 0.942021 -0.294156
+ 2.38e+10Hz 0.94164 -0.295346
+ 2.39e+10Hz 0.941259 -0.296536
+ 2.4e+10Hz 0.940875 -0.297725
+ 2.41e+10Hz 0.940491 -0.298914
+ 2.42e+10Hz 0.940104 -0.300102
+ 2.43e+10Hz 0.939716 -0.30129
+ 2.44e+10Hz 0.939326 -0.302477
+ 2.45e+10Hz 0.938935 -0.303664
+ 2.46e+10Hz 0.938542 -0.304851
+ 2.47e+10Hz 0.938148 -0.306037
+ 2.48e+10Hz 0.937751 -0.307222
+ 2.49e+10Hz 0.937354 -0.308407
+ 2.5e+10Hz 0.936955 -0.309592
+ 2.51e+10Hz 0.936554 -0.310776
+ 2.52e+10Hz 0.936152 -0.311959
+ 2.53e+10Hz 0.935748 -0.313142
+ 2.54e+10Hz 0.935342 -0.314324
+ 2.55e+10Hz 0.934935 -0.315506
+ 2.56e+10Hz 0.934526 -0.316687
+ 2.57e+10Hz 0.934116 -0.317868
+ 2.58e+10Hz 0.933704 -0.319048
+ 2.59e+10Hz 0.933291 -0.320228
+ 2.6e+10Hz 0.932876 -0.321407
+ 2.61e+10Hz 0.93246 -0.322585
+ 2.62e+10Hz 0.932042 -0.323763
+ 2.63e+10Hz 0.931622 -0.324941
+ 2.64e+10Hz 0.931201 -0.326117
+ 2.65e+10Hz 0.930778 -0.327294
+ 2.66e+10Hz 0.930354 -0.328469
+ 2.67e+10Hz 0.929928 -0.329644
+ 2.68e+10Hz 0.929501 -0.330819
+ 2.69e+10Hz 0.929072 -0.331992
+ 2.7e+10Hz 0.928642 -0.333166
+ 2.71e+10Hz 0.92821 -0.334338
+ 2.72e+10Hz 0.927777 -0.33551
+ 2.73e+10Hz 0.927342 -0.336682
+ 2.74e+10Hz 0.926905 -0.337852
+ 2.75e+10Hz 0.926467 -0.339022
+ 2.76e+10Hz 0.926028 -0.340192
+ 2.77e+10Hz 0.925587 -0.341361
+ 2.78e+10Hz 0.925144 -0.342529
+ 2.79e+10Hz 0.9247 -0.343697
+ 2.8e+10Hz 0.924255 -0.344864
+ 2.81e+10Hz 0.923808 -0.34603
+ 2.82e+10Hz 0.923359 -0.347196
+ 2.83e+10Hz 0.922909 -0.348361
+ 2.84e+10Hz 0.922458 -0.349525
+ 2.85e+10Hz 0.922005 -0.350689
+ 2.86e+10Hz 0.92155 -0.351852
+ 2.87e+10Hz 0.921094 -0.353015
+ 2.88e+10Hz 0.920637 -0.354176
+ 2.89e+10Hz 0.920178 -0.355337
+ 2.9e+10Hz 0.919718 -0.356498
+ 2.91e+10Hz 0.919256 -0.357658
+ 2.92e+10Hz 0.918793 -0.358817
+ 2.93e+10Hz 0.918328 -0.359975
+ 2.94e+10Hz 0.917862 -0.361133
+ 2.95e+10Hz 0.917394 -0.36229
+ 2.96e+10Hz 0.916925 -0.363447
+ 2.97e+10Hz 0.916455 -0.364603
+ 2.98e+10Hz 0.915983 -0.365758
+ 2.99e+10Hz 0.91551 -0.366912
+ 3e+10Hz 0.915035 -0.368066
+ 3.01e+10Hz 0.914559 -0.369219
+ 3.02e+10Hz 0.914081 -0.370372
+ 3.03e+10Hz 0.913602 -0.371524
+ 3.04e+10Hz 0.913121 -0.372675
+ 3.05e+10Hz 0.912639 -0.373825
+ 3.06e+10Hz 0.912156 -0.374975
+ 3.07e+10Hz 0.911671 -0.376124
+ 3.08e+10Hz 0.911185 -0.377272
+ 3.09e+10Hz 0.910698 -0.37842
+ 3.1e+10Hz 0.910209 -0.379567
+ 3.11e+10Hz 0.909718 -0.380713
+ 3.12e+10Hz 0.909227 -0.381859
+ 3.13e+10Hz 0.908733 -0.383004
+ 3.14e+10Hz 0.908239 -0.384148
+ 3.15e+10Hz 0.907743 -0.385292
+ 3.16e+10Hz 0.907246 -0.386435
+ 3.17e+10Hz 0.906747 -0.387577
+ 3.18e+10Hz 0.906247 -0.388719
+ 3.19e+10Hz 0.905745 -0.38986
+ 3.2e+10Hz 0.905242 -0.391
+ 3.21e+10Hz 0.904738 -0.392139
+ 3.22e+10Hz 0.904233 -0.393278
+ 3.23e+10Hz 0.903726 -0.394416
+ 3.24e+10Hz 0.903217 -0.395554
+ 3.25e+10Hz 0.902708 -0.396691
+ 3.26e+10Hz 0.902196 -0.397827
+ 3.27e+10Hz 0.901684 -0.398962
+ 3.28e+10Hz 0.90117 -0.400097
+ 3.29e+10Hz 0.900655 -0.401231
+ 3.3e+10Hz 0.900138 -0.402364
+ 3.31e+10Hz 0.899621 -0.403497
+ 3.32e+10Hz 0.899101 -0.404629
+ 3.33e+10Hz 0.898581 -0.405761
+ 3.34e+10Hz 0.898059 -0.406891
+ 3.35e+10Hz 0.897535 -0.408021
+ 3.36e+10Hz 0.897011 -0.40915
+ 3.37e+10Hz 0.896485 -0.410279
+ 3.38e+10Hz 0.895957 -0.411407
+ 3.39e+10Hz 0.895429 -0.412534
+ 3.4e+10Hz 0.894899 -0.413661
+ 3.41e+10Hz 0.894367 -0.414787
+ 3.42e+10Hz 0.893834 -0.415912
+ 3.43e+10Hz 0.8933 -0.417037
+ 3.44e+10Hz 0.892765 -0.418161
+ 3.45e+10Hz 0.892228 -0.419284
+ 3.46e+10Hz 0.89169 -0.420406
+ 3.47e+10Hz 0.89115 -0.421528
+ 3.48e+10Hz 0.890609 -0.42265
+ 3.49e+10Hz 0.890067 -0.42377
+ 3.5e+10Hz 0.889524 -0.42489
+ 3.51e+10Hz 0.888979 -0.426009
+ 3.52e+10Hz 0.888433 -0.427128
+ 3.53e+10Hz 0.887885 -0.428245
+ 3.54e+10Hz 0.887336 -0.429363
+ 3.55e+10Hz 0.886786 -0.430479
+ 3.56e+10Hz 0.886234 -0.431595
+ 3.57e+10Hz 0.885682 -0.43271
+ 3.58e+10Hz 0.885127 -0.433825
+ 3.59e+10Hz 0.884572 -0.434938
+ 3.6e+10Hz 0.884015 -0.436051
+ 3.61e+10Hz 0.883456 -0.437164
+ 3.62e+10Hz 0.882897 -0.438276
+ 3.63e+10Hz 0.882336 -0.439387
+ 3.64e+10Hz 0.881773 -0.440497
+ 3.65e+10Hz 0.88121 -0.441607
+ 3.66e+10Hz 0.880645 -0.442716
+ 3.67e+10Hz 0.880078 -0.443825
+ 3.68e+10Hz 0.879511 -0.444932
+ 3.69e+10Hz 0.878942 -0.446039
+ 3.7e+10Hz 0.878371 -0.447146
+ 3.71e+10Hz 0.8778 -0.448251
+ 3.72e+10Hz 0.877227 -0.449356
+ 3.73e+10Hz 0.876652 -0.450461
+ 3.74e+10Hz 0.876076 -0.451564
+ 3.75e+10Hz 0.875499 -0.452668
+ 3.76e+10Hz 0.874921 -0.45377
+ 3.77e+10Hz 0.874341 -0.454871
+ 3.78e+10Hz 0.87376 -0.455973
+ 3.79e+10Hz 0.873177 -0.457073
+ 3.8e+10Hz 0.872593 -0.458172
+ 3.81e+10Hz 0.872008 -0.459271
+ 3.82e+10Hz 0.871421 -0.46037
+ 3.83e+10Hz 0.870833 -0.461467
+ 3.84e+10Hz 0.870244 -0.462564
+ 3.85e+10Hz 0.869653 -0.46366
+ 3.86e+10Hz 0.869061 -0.464756
+ 3.87e+10Hz 0.868468 -0.465851
+ 3.88e+10Hz 0.867873 -0.466945
+ 3.89e+10Hz 0.867277 -0.468038
+ 3.9e+10Hz 0.86668 -0.469131
+ 3.91e+10Hz 0.866081 -0.470223
+ 3.92e+10Hz 0.865481 -0.471314
+ 3.93e+10Hz 0.864879 -0.472405
+ 3.94e+10Hz 0.864276 -0.473495
+ 3.95e+10Hz 0.863672 -0.474584
+ 3.96e+10Hz 0.863066 -0.475672
+ 3.97e+10Hz 0.862459 -0.47676
+ 3.98e+10Hz 0.861851 -0.477847
+ 3.99e+10Hz 0.861241 -0.478934
+ 4e+10Hz 0.86063 -0.48002
+ 4.01e+10Hz 0.860017 -0.481104
+ 4.02e+10Hz 0.859403 -0.482189
+ 4.03e+10Hz 0.858788 -0.483272
+ 4.04e+10Hz 0.858172 -0.484355
+ 4.05e+10Hz 0.857554 -0.485437
+ 4.06e+10Hz 0.856934 -0.486519
+ 4.07e+10Hz 0.856313 -0.487599
+ 4.08e+10Hz 0.855691 -0.488679
+ 4.09e+10Hz 0.855068 -0.489758
+ 4.1e+10Hz 0.854443 -0.490837
+ 4.11e+10Hz 0.853817 -0.491915
+ 4.12e+10Hz 0.853189 -0.492992
+ 4.13e+10Hz 0.85256 -0.494068
+ 4.14e+10Hz 0.85193 -0.495144
+ 4.15e+10Hz 0.851298 -0.496218
+ 4.16e+10Hz 0.850665 -0.497292
+ 4.17e+10Hz 0.85003 -0.498366
+ 4.18e+10Hz 0.849394 -0.499438
+ 4.19e+10Hz 0.848757 -0.50051
+ 4.2e+10Hz 0.848118 -0.501581
+ 4.21e+10Hz 0.847478 -0.502651
+ 4.22e+10Hz 0.846837 -0.503721
+ 4.23e+10Hz 0.846194 -0.504789
+ 4.24e+10Hz 0.84555 -0.505857
+ 4.25e+10Hz 0.844904 -0.506925
+ 4.26e+10Hz 0.844257 -0.507991
+ 4.27e+10Hz 0.843609 -0.509057
+ 4.28e+10Hz 0.842959 -0.510122
+ 4.29e+10Hz 0.842308 -0.511185
+ 4.3e+10Hz 0.841655 -0.512249
+ 4.31e+10Hz 0.841001 -0.513311
+ 4.32e+10Hz 0.840346 -0.514373
+ 4.33e+10Hz 0.839689 -0.515434
+ 4.34e+10Hz 0.839031 -0.516494
+ 4.35e+10Hz 0.838372 -0.517553
+ 4.36e+10Hz 0.837711 -0.518612
+ 4.37e+10Hz 0.837049 -0.51967
+ 4.38e+10Hz 0.836385 -0.520726
+ 4.39e+10Hz 0.83572 -0.521782
+ 4.4e+10Hz 0.835054 -0.522838
+ 4.41e+10Hz 0.834386 -0.523892
+ 4.42e+10Hz 0.833717 -0.524946
+ 4.43e+10Hz 0.833047 -0.525998
+ 4.44e+10Hz 0.832375 -0.52705
+ 4.45e+10Hz 0.831702 -0.528102
+ 4.46e+10Hz 0.831027 -0.529152
+ 4.47e+10Hz 0.830351 -0.530201
+ 4.48e+10Hz 0.829674 -0.53125
+ 4.49e+10Hz 0.828995 -0.532297
+ 4.5e+10Hz 0.828315 -0.533344
+ 4.51e+10Hz 0.827633 -0.53439
+ 4.52e+10Hz 0.826951 -0.535436
+ 4.53e+10Hz 0.826266 -0.53648
+ 4.54e+10Hz 0.825581 -0.537523
+ 4.55e+10Hz 0.824894 -0.538566
+ 4.56e+10Hz 0.824205 -0.539608
+ 4.57e+10Hz 0.823516 -0.540649
+ 4.58e+10Hz 0.822825 -0.541689
+ 4.59e+10Hz 0.822132 -0.542728
+ 4.6e+10Hz 0.821438 -0.543766
+ 4.61e+10Hz 0.820743 -0.544803
+ 4.62e+10Hz 0.820047 -0.54584
+ 4.63e+10Hz 0.819349 -0.546875
+ 4.64e+10Hz 0.81865 -0.54791
+ 4.65e+10Hz 0.817949 -0.548944
+ 4.66e+10Hz 0.817247 -0.549977
+ 4.67e+10Hz 0.816544 -0.551009
+ 4.68e+10Hz 0.815839 -0.55204
+ 4.69e+10Hz 0.815133 -0.55307
+ 4.7e+10Hz 0.814426 -0.554099
+ 4.71e+10Hz 0.813717 -0.555127
+ 4.72e+10Hz 0.813007 -0.556155
+ 4.73e+10Hz 0.812296 -0.557181
+ 4.74e+10Hz 0.811583 -0.558207
+ 4.75e+10Hz 0.810869 -0.559232
+ 4.76e+10Hz 0.810154 -0.560256
+ 4.77e+10Hz 0.809437 -0.561278
+ 4.78e+10Hz 0.808719 -0.5623
+ 4.79e+10Hz 0.808 -0.563321
+ 4.8e+10Hz 0.807279 -0.564341
+ 4.81e+10Hz 0.806557 -0.56536
+ 4.82e+10Hz 0.805834 -0.566378
+ 4.83e+10Hz 0.805109 -0.567396
+ 4.84e+10Hz 0.804383 -0.568412
+ 4.85e+10Hz 0.803656 -0.569427
+ 4.86e+10Hz 0.802927 -0.570441
+ 4.87e+10Hz 0.802198 -0.571455
+ 4.88e+10Hz 0.801466 -0.572467
+ 4.89e+10Hz 0.800734 -0.573479
+ 4.9e+10Hz 0.8 -0.574489
+ 4.91e+10Hz 0.799265 -0.575499
+ 4.92e+10Hz 0.798528 -0.576507
+ 4.93e+10Hz 0.797791 -0.577515
+ 4.94e+10Hz 0.797052 -0.578522
+ 4.95e+10Hz 0.796311 -0.579527
+ 4.96e+10Hz 0.79557 -0.580532
+ 4.97e+10Hz 0.794827 -0.581536
+ 4.98e+10Hz 0.794083 -0.582538
+ 4.99e+10Hz 0.793337 -0.58354
+ 5e+10Hz 0.79259 -0.584541
+ 5.01e+10Hz 0.791842 -0.585541
+ 5.02e+10Hz 0.791093 -0.58654
+ 5.03e+10Hz 0.790342 -0.587537
+ 5.04e+10Hz 0.78959 -0.588534
+ 5.05e+10Hz 0.788837 -0.58953
+ 5.06e+10Hz 0.788083 -0.590525
+ 5.07e+10Hz 0.787327 -0.591519
+ 5.08e+10Hz 0.78657 -0.592512
+ 5.09e+10Hz 0.785812 -0.593503
+ 5.1e+10Hz 0.785053 -0.594494
+ 5.11e+10Hz 0.784292 -0.595484
+ 5.12e+10Hz 0.78353 -0.596473
+ 5.13e+10Hz 0.782767 -0.597461
+ 5.14e+10Hz 0.782002 -0.598448
+ 5.15e+10Hz 0.781236 -0.599434
+ 5.16e+10Hz 0.780469 -0.600418
+ 5.17e+10Hz 0.779701 -0.601402
+ 5.18e+10Hz 0.778932 -0.602385
+ 5.19e+10Hz 0.778161 -0.603367
+ 5.2e+10Hz 0.777389 -0.604348
+ 5.21e+10Hz 0.776616 -0.605328
+ 5.22e+10Hz 0.775841 -0.606306
+ 5.23e+10Hz 0.775066 -0.607284
+ 5.24e+10Hz 0.774289 -0.608261
+ 5.25e+10Hz 0.773511 -0.609236
+ 5.26e+10Hz 0.772732 -0.610211
+ 5.27e+10Hz 0.771951 -0.611185
+ 5.28e+10Hz 0.771169 -0.612157
+ 5.29e+10Hz 0.770386 -0.613129
+ 5.3e+10Hz 0.769602 -0.6141
+ 5.31e+10Hz 0.768817 -0.615069
+ 5.32e+10Hz 0.76803 -0.616038
+ 5.33e+10Hz 0.767242 -0.617005
+ 5.34e+10Hz 0.766453 -0.617972
+ 5.35e+10Hz 0.765663 -0.618937
+ 5.36e+10Hz 0.764871 -0.619902
+ 5.37e+10Hz 0.764079 -0.620865
+ 5.38e+10Hz 0.763285 -0.621827
+ 5.39e+10Hz 0.76249 -0.622789
+ 5.4e+10Hz 0.761694 -0.623749
+ 5.41e+10Hz 0.760896 -0.624708
+ 5.42e+10Hz 0.760097 -0.625667
+ 5.43e+10Hz 0.759298 -0.626624
+ 5.44e+10Hz 0.758497 -0.62758
+ 5.45e+10Hz 0.757695 -0.628535
+ 5.46e+10Hz 0.756891 -0.629489
+ 5.47e+10Hz 0.756086 -0.630442
+ 5.48e+10Hz 0.755281 -0.631394
+ 5.49e+10Hz 0.754474 -0.632345
+ 5.5e+10Hz 0.753666 -0.633295
+ 5.51e+10Hz 0.752856 -0.634244
+ 5.52e+10Hz 0.752046 -0.635192
+ 5.53e+10Hz 0.751234 -0.636139
+ 5.54e+10Hz 0.750421 -0.637085
+ 5.55e+10Hz 0.749607 -0.638029
+ 5.56e+10Hz 0.748792 -0.638973
+ 5.57e+10Hz 0.747976 -0.639916
+ 5.58e+10Hz 0.747159 -0.640857
+ 5.59e+10Hz 0.74634 -0.641798
+ 5.6e+10Hz 0.74552 -0.642737
+ 5.61e+10Hz 0.744699 -0.643676
+ 5.62e+10Hz 0.743877 -0.644613
+ 5.63e+10Hz 0.743054 -0.64555
+ 5.64e+10Hz 0.742229 -0.646485
+ 5.65e+10Hz 0.741404 -0.647419
+ 5.66e+10Hz 0.740577 -0.648352
+ 5.67e+10Hz 0.739749 -0.649285
+ 5.68e+10Hz 0.73892 -0.650216
+ 5.69e+10Hz 0.73809 -0.651146
+ 5.7e+10Hz 0.737258 -0.652075
+ 5.71e+10Hz 0.736426 -0.653003
+ 5.72e+10Hz 0.735592 -0.65393
+ 5.73e+10Hz 0.734757 -0.654856
+ 5.74e+10Hz 0.733921 -0.65578
+ 5.75e+10Hz 0.733084 -0.656704
+ 5.76e+10Hz 0.732246 -0.657627
+ 5.77e+10Hz 0.731406 -0.658549
+ 5.78e+10Hz 0.730566 -0.659469
+ 5.79e+10Hz 0.729724 -0.660389
+ 5.8e+10Hz 0.728881 -0.661307
+ 5.81e+10Hz 0.728037 -0.662225
+ 5.82e+10Hz 0.727192 -0.663141
+ 5.83e+10Hz 0.726346 -0.664056
+ 5.84e+10Hz 0.725498 -0.664971
+ 5.85e+10Hz 0.72465 -0.665884
+ 5.86e+10Hz 0.7238 -0.666796
+ 5.87e+10Hz 0.722949 -0.667707
+ 5.88e+10Hz 0.722097 -0.668617
+ 5.89e+10Hz 0.721244 -0.669526
+ 5.9e+10Hz 0.72039 -0.670434
+ 5.91e+10Hz 0.719535 -0.67134
+ 5.92e+10Hz 0.718678 -0.672246
+ 5.93e+10Hz 0.71782 -0.673151
+ 5.94e+10Hz 0.716962 -0.674054
+ 5.95e+10Hz 0.716102 -0.674957
+ 5.96e+10Hz 0.715241 -0.675858
+ 5.97e+10Hz 0.714379 -0.676759
+ 5.98e+10Hz 0.713515 -0.677658
+ 5.99e+10Hz 0.712651 -0.678556
+ 6e+10Hz 0.711785 -0.679453
+ 6.01e+10Hz 0.710919 -0.680349
+ 6.02e+10Hz 0.710051 -0.681244
+ 6.03e+10Hz 0.709182 -0.682138
+ 6.04e+10Hz 0.708312 -0.683031
+ 6.05e+10Hz 0.707441 -0.683923
+ 6.06e+10Hz 0.706568 -0.684813
+ 6.07e+10Hz 0.705695 -0.685703
+ 6.08e+10Hz 0.70482 -0.686592
+ 6.09e+10Hz 0.703944 -0.687479
+ 6.1e+10Hz 0.703068 -0.688365
+ 6.11e+10Hz 0.70219 -0.68925
+ 6.12e+10Hz 0.701311 -0.690135
+ 6.13e+10Hz 0.70043 -0.691018
+ 6.14e+10Hz 0.699549 -0.6919
+ 6.15e+10Hz 0.698667 -0.69278
+ 6.16e+10Hz 0.697783 -0.69366
+ 6.17e+10Hz 0.696899 -0.694539
+ 6.18e+10Hz 0.696013 -0.695416
+ 6.19e+10Hz 0.695126 -0.696293
+ 6.2e+10Hz 0.694238 -0.697168
+ 6.21e+10Hz 0.693349 -0.698042
+ 6.22e+10Hz 0.692458 -0.698916
+ 6.23e+10Hz 0.691567 -0.699788
+ 6.24e+10Hz 0.690674 -0.700658
+ 6.25e+10Hz 0.689781 -0.701528
+ 6.26e+10Hz 0.688886 -0.702397
+ 6.27e+10Hz 0.68799 -0.703264
+ 6.28e+10Hz 0.687093 -0.704131
+ 6.29e+10Hz 0.686195 -0.704996
+ 6.3e+10Hz 0.685296 -0.705861
+ 6.31e+10Hz 0.684396 -0.706724
+ 6.32e+10Hz 0.683494 -0.707586
+ 6.33e+10Hz 0.682592 -0.708446
+ 6.34e+10Hz 0.681688 -0.709306
+ 6.35e+10Hz 0.680783 -0.710165
+ 6.36e+10Hz 0.679878 -0.711022
+ 6.37e+10Hz 0.678971 -0.711878
+ 6.38e+10Hz 0.678063 -0.712734
+ 6.39e+10Hz 0.677153 -0.713588
+ 6.4e+10Hz 0.676243 -0.714441
+ 6.41e+10Hz 0.675332 -0.715292
+ 6.42e+10Hz 0.674419 -0.716143
+ 6.43e+10Hz 0.673506 -0.716992
+ 6.44e+10Hz 0.672591 -0.717841
+ 6.45e+10Hz 0.671675 -0.718688
+ 6.46e+10Hz 0.670758 -0.719534
+ 6.47e+10Hz 0.66984 -0.720379
+ 6.48e+10Hz 0.668921 -0.721222
+ 6.49e+10Hz 0.668001 -0.722065
+ 6.5e+10Hz 0.66708 -0.722907
+ 6.51e+10Hz 0.666157 -0.723747
+ 6.52e+10Hz 0.665234 -0.724586
+ 6.53e+10Hz 0.664309 -0.725424
+ 6.54e+10Hz 0.663384 -0.72626
+ 6.55e+10Hz 0.662457 -0.727096
+ 6.56e+10Hz 0.661529 -0.72793
+ 6.57e+10Hz 0.6606 -0.728764
+ 6.58e+10Hz 0.65967 -0.729595
+ 6.59e+10Hz 0.658739 -0.730426
+ 6.6e+10Hz 0.657807 -0.731256
+ 6.61e+10Hz 0.656874 -0.732085
+ 6.62e+10Hz 0.655939 -0.732912
+ 6.63e+10Hz 0.655004 -0.733738
+ 6.64e+10Hz 0.654067 -0.734563
+ 6.65e+10Hz 0.65313 -0.735387
+ 6.66e+10Hz 0.652191 -0.736209
+ 6.67e+10Hz 0.651251 -0.73703
+ 6.68e+10Hz 0.650311 -0.73785
+ 6.69e+10Hz 0.649369 -0.738669
+ 6.7e+10Hz 0.648426 -0.739487
+ 6.71e+10Hz 0.647482 -0.740304
+ 6.72e+10Hz 0.646536 -0.741119
+ 6.73e+10Hz 0.64559 -0.741933
+ 6.74e+10Hz 0.644643 -0.742746
+ 6.75e+10Hz 0.643695 -0.743558
+ 6.76e+10Hz 0.642745 -0.744368
+ 6.77e+10Hz 0.641795 -0.745177
+ 6.78e+10Hz 0.640844 -0.745985
+ 6.79e+10Hz 0.639891 -0.746792
+ 6.8e+10Hz 0.638937 -0.747598
+ 6.81e+10Hz 0.637983 -0.748402
+ 6.82e+10Hz 0.637027 -0.749205
+ 6.83e+10Hz 0.63607 -0.750007
+ 6.84e+10Hz 0.635113 -0.750807
+ 6.85e+10Hz 0.634154 -0.751607
+ 6.86e+10Hz 0.633194 -0.752405
+ 6.87e+10Hz 0.632233 -0.753202
+ 6.88e+10Hz 0.631271 -0.753997
+ 6.89e+10Hz 0.630308 -0.754792
+ 6.9e+10Hz 0.629344 -0.755585
+ 6.91e+10Hz 0.628379 -0.756377
+ 6.92e+10Hz 0.627413 -0.757168
+ 6.93e+10Hz 0.626446 -0.757957
+ 6.94e+10Hz 0.625478 -0.758745
+ 6.95e+10Hz 0.624508 -0.759532
+ 6.96e+10Hz 0.623538 -0.760318
+ 6.97e+10Hz 0.622567 -0.761102
+ 6.98e+10Hz 0.621595 -0.761885
+ 6.99e+10Hz 0.620621 -0.762667
+ 7e+10Hz 0.619647 -0.763448
+ 7.01e+10Hz 0.618672 -0.764227
+ 7.02e+10Hz 0.617696 -0.765005
+ 7.03e+10Hz 0.616718 -0.765782
+ 7.04e+10Hz 0.61574 -0.766557
+ 7.05e+10Hz 0.614761 -0.767331
+ 7.06e+10Hz 0.61378 -0.768104
+ 7.07e+10Hz 0.612799 -0.768876
+ 7.08e+10Hz 0.611817 -0.769646
+ 7.09e+10Hz 0.610834 -0.770415
+ 7.1e+10Hz 0.609849 -0.771183
+ 7.11e+10Hz 0.608864 -0.77195
+ 7.12e+10Hz 0.607878 -0.772715
+ 7.13e+10Hz 0.60689 -0.773479
+ 7.14e+10Hz 0.605902 -0.774242
+ 7.15e+10Hz 0.604913 -0.775003
+ 7.16e+10Hz 0.603923 -0.775763
+ 7.17e+10Hz 0.602932 -0.776522
+ 7.18e+10Hz 0.601939 -0.777279
+ 7.19e+10Hz 0.600946 -0.778035
+ 7.2e+10Hz 0.599952 -0.77879
+ 7.21e+10Hz 0.598957 -0.779544
+ 7.22e+10Hz 0.597961 -0.780296
+ 7.23e+10Hz 0.596964 -0.781047
+ 7.24e+10Hz 0.595966 -0.781796
+ 7.25e+10Hz 0.594968 -0.782545
+ 7.26e+10Hz 0.593968 -0.783292
+ 7.27e+10Hz 0.592967 -0.784038
+ 7.28e+10Hz 0.591965 -0.784782
+ 7.29e+10Hz 0.590963 -0.785525
+ 7.3e+10Hz 0.589959 -0.786267
+ 7.31e+10Hz 0.588954 -0.787007
+ 7.32e+10Hz 0.587949 -0.787746
+ 7.33e+10Hz 0.586943 -0.788484
+ 7.34e+10Hz 0.585935 -0.789221
+ 7.35e+10Hz 0.584927 -0.789956
+ 7.36e+10Hz 0.583918 -0.79069
+ 7.37e+10Hz 0.582908 -0.791422
+ 7.38e+10Hz 0.581897 -0.792153
+ 7.39e+10Hz 0.580885 -0.792883
+ 7.4e+10Hz 0.579872 -0.793612
+ 7.41e+10Hz 0.578858 -0.794339
+ 7.42e+10Hz 0.577843 -0.795065
+ 7.43e+10Hz 0.576828 -0.79579
+ 7.44e+10Hz 0.575811 -0.796513
+ 7.45e+10Hz 0.574793 -0.797235
+ 7.46e+10Hz 0.573775 -0.797956
+ 7.47e+10Hz 0.572756 -0.798675
+ 7.48e+10Hz 0.571736 -0.799393
+ 7.49e+10Hz 0.570715 -0.80011
+ 7.5e+10Hz 0.569693 -0.800825
+ 7.51e+10Hz 0.56867 -0.801539
+ 7.52e+10Hz 0.567646 -0.802251
+ 7.53e+10Hz 0.566622 -0.802963
+ 7.54e+10Hz 0.565596 -0.803673
+ 7.55e+10Hz 0.56457 -0.804381
+ 7.56e+10Hz 0.563542 -0.805089
+ 7.57e+10Hz 0.562514 -0.805795
+ 7.58e+10Hz 0.561485 -0.806499
+ 7.59e+10Hz 0.560455 -0.807203
+ 7.6e+10Hz 0.559425 -0.807904
+ 7.61e+10Hz 0.558393 -0.808605
+ 7.62e+10Hz 0.557361 -0.809304
+ 7.63e+10Hz 0.556327 -0.810002
+ 7.64e+10Hz 0.555293 -0.810699
+ 7.65e+10Hz 0.554258 -0.811394
+ 7.66e+10Hz 0.553222 -0.812088
+ 7.67e+10Hz 0.552185 -0.812781
+ 7.68e+10Hz 0.551147 -0.813472
+ 7.69e+10Hz 0.550109 -0.814162
+ 7.7e+10Hz 0.54907 -0.81485
+ 7.71e+10Hz 0.548029 -0.815537
+ 7.72e+10Hz 0.546988 -0.816223
+ 7.73e+10Hz 0.545946 -0.816908
+ 7.74e+10Hz 0.544904 -0.817591
+ 7.75e+10Hz 0.54386 -0.818273
+ 7.76e+10Hz 0.542816 -0.818953
+ 7.77e+10Hz 0.54177 -0.819632
+ 7.78e+10Hz 0.540724 -0.82031
+ 7.79e+10Hz 0.539677 -0.820987
+ 7.8e+10Hz 0.53863 -0.821662
+ 7.81e+10Hz 0.537581 -0.822335
+ 7.82e+10Hz 0.536532 -0.823008
+ 7.83e+10Hz 0.535481 -0.823679
+ 7.84e+10Hz 0.53443 -0.824349
+ 7.85e+10Hz 0.533378 -0.825017
+ 7.86e+10Hz 0.532326 -0.825684
+ 7.87e+10Hz 0.531272 -0.82635
+ 7.88e+10Hz 0.530218 -0.827014
+ 7.89e+10Hz 0.529163 -0.827677
+ 7.9e+10Hz 0.528107 -0.828339
+ 7.91e+10Hz 0.52705 -0.828999
+ 7.92e+10Hz 0.525992 -0.829658
+ 7.93e+10Hz 0.524934 -0.830315
+ 7.94e+10Hz 0.523875 -0.830972
+ 7.95e+10Hz 0.522815 -0.831627
+ 7.96e+10Hz 0.521754 -0.83228
+ 7.97e+10Hz 0.520692 -0.832932
+ 7.98e+10Hz 0.51963 -0.833583
+ 7.99e+10Hz 0.518567 -0.834233
+ 8e+10Hz 0.517502 -0.834881
+ 8.01e+10Hz 0.516438 -0.835527
+ 8.02e+10Hz 0.515372 -0.836173
+ 8.03e+10Hz 0.514305 -0.836817
+ 8.04e+10Hz 0.513238 -0.83746
+ 8.05e+10Hz 0.51217 -0.838101
+ 8.06e+10Hz 0.511101 -0.838741
+ 8.07e+10Hz 0.510032 -0.83938
+ 8.08e+10Hz 0.508961 -0.840017
+ 8.09e+10Hz 0.50789 -0.840653
+ 8.1e+10Hz 0.506818 -0.841287
+ 8.11e+10Hz 0.505746 -0.841921
+ 8.12e+10Hz 0.504672 -0.842553
+ 8.13e+10Hz 0.503598 -0.843183
+ 8.14e+10Hz 0.502523 -0.843812
+ 8.15e+10Hz 0.501447 -0.84444
+ 8.16e+10Hz 0.50037 -0.845066
+ 8.17e+10Hz 0.499293 -0.845692
+ 8.18e+10Hz 0.498214 -0.846315
+ 8.19e+10Hz 0.497135 -0.846938
+ 8.2e+10Hz 0.496056 -0.847559
+ 8.21e+10Hz 0.494975 -0.848178
+ 8.22e+10Hz 0.493894 -0.848796
+ 8.23e+10Hz 0.492812 -0.849413
+ 8.24e+10Hz 0.491729 -0.850029
+ 8.25e+10Hz 0.490645 -0.850643
+ 8.26e+10Hz 0.489561 -0.851256
+ 8.27e+10Hz 0.488476 -0.851867
+ 8.28e+10Hz 0.48739 -0.852477
+ 8.29e+10Hz 0.486303 -0.853086
+ 8.3e+10Hz 0.485216 -0.853693
+ 8.31e+10Hz 0.484127 -0.854299
+ 8.32e+10Hz 0.483038 -0.854904
+ 8.33e+10Hz 0.481949 -0.855507
+ 8.34e+10Hz 0.480858 -0.856109
+ 8.35e+10Hz 0.479767 -0.85671
+ 8.36e+10Hz 0.478675 -0.857309
+ 8.37e+10Hz 0.477582 -0.857907
+ 8.38e+10Hz 0.476488 -0.858503
+ 8.39e+10Hz 0.475394 -0.859098
+ 8.4e+10Hz 0.474299 -0.859691
+ 8.41e+10Hz 0.473203 -0.860284
+ 8.42e+10Hz 0.472107 -0.860874
+ 8.43e+10Hz 0.47101 -0.861464
+ 8.44e+10Hz 0.469911 -0.862052
+ 8.45e+10Hz 0.468813 -0.862639
+ 8.46e+10Hz 0.467713 -0.863224
+ 8.47e+10Hz 0.466613 -0.863808
+ 8.48e+10Hz 0.465512 -0.864391
+ 8.49e+10Hz 0.46441 -0.864972
+ 8.5e+10Hz 0.463307 -0.865552
+ 8.51e+10Hz 0.462204 -0.86613
+ 8.52e+10Hz 0.4611 -0.866707
+ 8.53e+10Hz 0.459996 -0.867282
+ 8.54e+10Hz 0.45889 -0.867857
+ 8.55e+10Hz 0.457784 -0.868429
+ 8.56e+10Hz 0.456677 -0.869001
+ 8.57e+10Hz 0.455569 -0.869571
+ 8.58e+10Hz 0.454461 -0.870139
+ 8.59e+10Hz 0.453352 -0.870707
+ 8.6e+10Hz 0.452242 -0.871273
+ 8.61e+10Hz 0.451131 -0.871837
+ 8.62e+10Hz 0.45002 -0.8724
+ 8.63e+10Hz 0.448908 -0.872962
+ 8.64e+10Hz 0.447795 -0.873522
+ 8.65e+10Hz 0.446681 -0.874081
+ 8.66e+10Hz 0.445567 -0.874638
+ 8.67e+10Hz 0.444452 -0.875194
+ 8.68e+10Hz 0.443336 -0.875748
+ 8.69e+10Hz 0.44222 -0.876302
+ 8.7e+10Hz 0.441103 -0.876853
+ 8.71e+10Hz 0.439985 -0.877404
+ 8.72e+10Hz 0.438866 -0.877953
+ 8.73e+10Hz 0.437747 -0.8785
+ 8.74e+10Hz 0.436627 -0.879046
+ 8.75e+10Hz 0.435506 -0.879591
+ 8.76e+10Hz 0.434385 -0.880134
+ 8.77e+10Hz 0.433262 -0.880676
+ 8.78e+10Hz 0.43214 -0.881216
+ 8.79e+10Hz 0.431016 -0.881755
+ 8.8e+10Hz 0.429892 -0.882292
+ 8.81e+10Hz 0.428767 -0.882828
+ 8.82e+10Hz 0.427641 -0.883363
+ 8.83e+10Hz 0.426515 -0.883896
+ 8.84e+10Hz 0.425388 -0.884428
+ 8.85e+10Hz 0.42426 -0.884958
+ 8.86e+10Hz 0.423132 -0.885487
+ 8.87e+10Hz 0.422003 -0.886015
+ 8.88e+10Hz 0.420873 -0.88654
+ 8.89e+10Hz 0.419742 -0.887065
+ 8.9e+10Hz 0.418611 -0.887588
+ 8.91e+10Hz 0.417479 -0.88811
+ 8.92e+10Hz 0.416346 -0.88863
+ 8.93e+10Hz 0.415213 -0.889149
+ 8.94e+10Hz 0.414079 -0.889666
+ 8.95e+10Hz 0.412945 -0.890182
+ 8.96e+10Hz 0.411809 -0.890696
+ 8.97e+10Hz 0.410673 -0.891209
+ 8.98e+10Hz 0.409537 -0.89172
+ 8.99e+10Hz 0.408399 -0.89223
+ 9e+10Hz 0.407261 -0.892739
+ 9.01e+10Hz 0.406123 -0.893246
+ 9.02e+10Hz 0.404983 -0.893751
+ 9.03e+10Hz 0.403843 -0.894255
+ 9.04e+10Hz 0.402703 -0.894758
+ 9.05e+10Hz 0.401562 -0.895259
+ 9.06e+10Hz 0.40042 -0.895759
+ 9.07e+10Hz 0.399277 -0.896257
+ 9.08e+10Hz 0.398134 -0.896754
+ 9.09e+10Hz 0.39699 -0.897249
+ 9.1e+10Hz 0.395845 -0.897743
+ 9.11e+10Hz 0.3947 -0.898235
+ 9.12e+10Hz 0.393554 -0.898726
+ 9.13e+10Hz 0.392408 -0.899215
+ 9.14e+10Hz 0.391261 -0.899703
+ 9.15e+10Hz 0.390113 -0.90019
+ 9.16e+10Hz 0.388965 -0.900675
+ 9.17e+10Hz 0.387816 -0.901158
+ 9.18e+10Hz 0.386666 -0.90164
+ 9.19e+10Hz 0.385516 -0.90212
+ 9.2e+10Hz 0.384365 -0.902599
+ 9.21e+10Hz 0.383213 -0.903077
+ 9.22e+10Hz 0.382061 -0.903552
+ 9.23e+10Hz 0.380908 -0.904027
+ 9.24e+10Hz 0.379755 -0.9045
+ 9.25e+10Hz 0.378601 -0.904971
+ 9.26e+10Hz 0.377447 -0.905441
+ 9.27e+10Hz 0.376292 -0.90591
+ 9.28e+10Hz 0.375136 -0.906377
+ 9.29e+10Hz 0.373979 -0.906842
+ 9.3e+10Hz 0.372822 -0.907306
+ 9.31e+10Hz 0.371665 -0.907768
+ 9.32e+10Hz 0.370507 -0.908229
+ 9.33e+10Hz 0.369348 -0.908689
+ 9.34e+10Hz 0.368189 -0.909146
+ 9.35e+10Hz 0.367029 -0.909603
+ 9.36e+10Hz 0.365868 -0.910057
+ 9.37e+10Hz 0.364707 -0.910511
+ 9.38e+10Hz 0.363546 -0.910963
+ 9.39e+10Hz 0.362383 -0.911413
+ 9.4e+10Hz 0.361221 -0.911862
+ 9.41e+10Hz 0.360057 -0.912309
+ 9.42e+10Hz 0.358893 -0.912755
+ 9.43e+10Hz 0.357729 -0.913199
+ 9.44e+10Hz 0.356564 -0.913642
+ 9.45e+10Hz 0.355398 -0.914083
+ 9.46e+10Hz 0.354232 -0.914523
+ 9.47e+10Hz 0.353066 -0.914961
+ 9.48e+10Hz 0.351898 -0.915397
+ 9.49e+10Hz 0.350731 -0.915833
+ 9.5e+10Hz 0.349562 -0.916266
+ 9.51e+10Hz 0.348394 -0.916698
+ 9.52e+10Hz 0.347224 -0.917129
+ 9.53e+10Hz 0.346054 -0.917558
+ 9.54e+10Hz 0.344884 -0.917985
+ 9.55e+10Hz 0.343713 -0.918411
+ 9.56e+10Hz 0.342541 -0.918836
+ 9.57e+10Hz 0.341369 -0.919258
+ 9.58e+10Hz 0.340197 -0.91968
+ 9.59e+10Hz 0.339024 -0.9201
+ 9.6e+10Hz 0.33785 -0.920518
+ 9.61e+10Hz 0.336676 -0.920935
+ 9.62e+10Hz 0.335502 -0.92135
+ 9.63e+10Hz 0.334326 -0.921764
+ 9.64e+10Hz 0.333151 -0.922176
+ 9.65e+10Hz 0.331975 -0.922586
+ 9.66e+10Hz 0.330798 -0.922996
+ 9.67e+10Hz 0.329621 -0.923403
+ 9.68e+10Hz 0.328444 -0.923809
+ 9.69e+10Hz 0.327266 -0.924214
+ 9.7e+10Hz 0.326087 -0.924617
+ 9.71e+10Hz 0.324908 -0.925018
+ 9.72e+10Hz 0.323728 -0.925418
+ 9.73e+10Hz 0.322549 -0.925817
+ 9.74e+10Hz 0.321368 -0.926214
+ 9.75e+10Hz 0.320187 -0.926609
+ 9.76e+10Hz 0.319006 -0.927003
+ 9.77e+10Hz 0.317824 -0.927395
+ 9.78e+10Hz 0.316642 -0.927786
+ 9.79e+10Hz 0.315459 -0.928175
+ 9.8e+10Hz 0.314276 -0.928563
+ 9.81e+10Hz 0.313092 -0.928949
+ 9.82e+10Hz 0.311908 -0.929334
+ 9.83e+10Hz 0.310723 -0.929717
+ 9.84e+10Hz 0.309538 -0.930098
+ 9.85e+10Hz 0.308353 -0.930478
+ 9.86e+10Hz 0.307167 -0.930857
+ 9.87e+10Hz 0.30598 -0.931234
+ 9.88e+10Hz 0.304794 -0.931609
+ 9.89e+10Hz 0.303606 -0.931983
+ 9.9e+10Hz 0.302419 -0.932356
+ 9.91e+10Hz 0.301231 -0.932727
+ 9.92e+10Hz 0.300042 -0.933096
+ 9.93e+10Hz 0.298853 -0.933464
+ 9.94e+10Hz 0.297664 -0.93383
+ 9.95e+10Hz 0.296474 -0.934195
+ 9.96e+10Hz 0.295284 -0.934558
+ 9.97e+10Hz 0.294093 -0.93492
+ 9.98e+10Hz 0.292902 -0.93528
+ 9.99e+10Hz 0.29171 -0.935639
+ 1e+11Hz 0.290519 -0.935996
+ 1.001e+11Hz 0.289326 -0.936352
+ 1.002e+11Hz 0.288133 -0.936706
+ 1.003e+11Hz 0.28694 -0.937059
+ 1.004e+11Hz 0.285747 -0.93741
+ 1.005e+11Hz 0.284553 -0.937759
+ 1.006e+11Hz 0.283359 -0.938107
+ 1.007e+11Hz 0.282164 -0.938454
+ 1.008e+11Hz 0.280969 -0.938799
+ 1.009e+11Hz 0.279773 -0.939142
+ 1.01e+11Hz 0.278577 -0.939484
+ 1.011e+11Hz 0.277381 -0.939825
+ 1.012e+11Hz 0.276184 -0.940164
+ 1.013e+11Hz 0.274987 -0.940501
+ 1.014e+11Hz 0.27379 -0.940837
+ 1.015e+11Hz 0.272592 -0.941171
+ 1.016e+11Hz 0.271394 -0.941504
+ 1.017e+11Hz 0.270195 -0.941835
+ 1.018e+11Hz 0.268996 -0.942165
+ 1.019e+11Hz 0.267797 -0.942494
+ 1.02e+11Hz 0.266597 -0.94282
+ 1.021e+11Hz 0.265397 -0.943146
+ 1.022e+11Hz 0.264197 -0.943469
+ 1.023e+11Hz 0.262996 -0.943792
+ 1.024e+11Hz 0.261794 -0.944112
+ 1.025e+11Hz 0.260593 -0.944432
+ 1.026e+11Hz 0.259391 -0.944749
+ 1.027e+11Hz 0.258189 -0.945066
+ 1.028e+11Hz 0.256986 -0.94538
+ 1.029e+11Hz 0.255783 -0.945693
+ 1.03e+11Hz 0.25458 -0.946005
+ 1.031e+11Hz 0.253376 -0.946315
+ 1.032e+11Hz 0.252172 -0.946624
+ 1.033e+11Hz 0.250967 -0.946931
+ 1.034e+11Hz 0.249762 -0.947237
+ 1.035e+11Hz 0.248557 -0.947541
+ 1.036e+11Hz 0.247352 -0.947844
+ 1.037e+11Hz 0.246146 -0.948145
+ 1.038e+11Hz 0.24494 -0.948444
+ 1.039e+11Hz 0.243733 -0.948743
+ 1.04e+11Hz 0.242526 -0.949039
+ 1.041e+11Hz 0.241319 -0.949334
+ 1.042e+11Hz 0.240111 -0.949628
+ 1.043e+11Hz 0.238903 -0.94992
+ 1.044e+11Hz 0.237695 -0.95021
+ 1.045e+11Hz 0.236486 -0.9505
+ 1.046e+11Hz 0.235277 -0.950787
+ 1.047e+11Hz 0.234068 -0.951073
+ 1.048e+11Hz 0.232858 -0.951358
+ 1.049e+11Hz 0.231648 -0.951641
+ 1.05e+11Hz 0.230438 -0.951922
+ 1.051e+11Hz 0.229227 -0.952202
+ 1.052e+11Hz 0.228016 -0.952481
+ 1.053e+11Hz 0.226805 -0.952758
+ 1.054e+11Hz 0.225593 -0.953033
+ 1.055e+11Hz 0.224381 -0.953307
+ 1.056e+11Hz 0.223168 -0.95358
+ 1.057e+11Hz 0.221956 -0.953851
+ 1.058e+11Hz 0.220743 -0.954121
+ 1.059e+11Hz 0.219529 -0.954388
+ 1.06e+11Hz 0.218316 -0.954655
+ 1.061e+11Hz 0.217102 -0.95492
+ 1.062e+11Hz 0.215887 -0.955183
+ 1.063e+11Hz 0.214673 -0.955445
+ 1.064e+11Hz 0.213458 -0.955706
+ 1.065e+11Hz 0.212242 -0.955965
+ 1.066e+11Hz 0.211027 -0.956222
+ 1.067e+11Hz 0.209811 -0.956478
+ 1.068e+11Hz 0.208594 -0.956732
+ 1.069e+11Hz 0.207378 -0.956985
+ 1.07e+11Hz 0.206161 -0.957237
+ 1.071e+11Hz 0.204944 -0.957487
+ 1.072e+11Hz 0.203726 -0.957735
+ 1.073e+11Hz 0.202508 -0.957982
+ 1.074e+11Hz 0.20129 -0.958227
+ 1.075e+11Hz 0.200071 -0.958471
+ 1.076e+11Hz 0.198852 -0.958713
+ 1.077e+11Hz 0.197633 -0.958954
+ 1.078e+11Hz 0.196414 -0.959193
+ 1.079e+11Hz 0.195194 -0.959431
+ 1.08e+11Hz 0.193974 -0.959667
+ 1.081e+11Hz 0.192754 -0.959902
+ 1.082e+11Hz 0.191533 -0.960135
+ 1.083e+11Hz 0.190312 -0.960367
+ 1.084e+11Hz 0.189091 -0.960597
+ 1.085e+11Hz 0.187869 -0.960825
+ 1.086e+11Hz 0.186647 -0.961052
+ 1.087e+11Hz 0.185425 -0.961278
+ 1.088e+11Hz 0.184202 -0.961502
+ 1.089e+11Hz 0.182979 -0.961724
+ 1.09e+11Hz 0.181756 -0.961945
+ 1.091e+11Hz 0.180533 -0.962165
+ 1.092e+11Hz 0.179309 -0.962383
+ 1.093e+11Hz 0.178085 -0.962599
+ 1.094e+11Hz 0.176861 -0.962814
+ 1.095e+11Hz 0.175636 -0.963027
+ 1.096e+11Hz 0.174411 -0.963239
+ 1.097e+11Hz 0.173186 -0.963449
+ 1.098e+11Hz 0.171961 -0.963658
+ 1.099e+11Hz 0.170735 -0.963865
+ 1.1e+11Hz 0.169509 -0.964071
+ 1.101e+11Hz 0.168283 -0.964275
+ 1.102e+11Hz 0.167056 -0.964477
+ 1.103e+11Hz 0.165829 -0.964678
+ 1.104e+11Hz 0.164602 -0.964877
+ 1.105e+11Hz 0.163374 -0.965075
+ 1.106e+11Hz 0.162147 -0.965272
+ 1.107e+11Hz 0.160919 -0.965466
+ 1.108e+11Hz 0.15969 -0.96566
+ 1.109e+11Hz 0.158462 -0.965851
+ 1.11e+11Hz 0.157233 -0.966041
+ 1.111e+11Hz 0.156004 -0.96623
+ 1.112e+11Hz 0.154774 -0.966417
+ 1.113e+11Hz 0.153545 -0.966602
+ 1.114e+11Hz 0.152315 -0.966786
+ 1.115e+11Hz 0.151085 -0.966968
+ 1.116e+11Hz 0.149854 -0.967149
+ 1.117e+11Hz 0.148624 -0.967328
+ 1.118e+11Hz 0.147393 -0.967506
+ 1.119e+11Hz 0.146161 -0.967682
+ 1.12e+11Hz 0.14493 -0.967856
+ 1.121e+11Hz 0.143698 -0.968029
+ 1.122e+11Hz 0.142466 -0.968201
+ 1.123e+11Hz 0.141234 -0.96837
+ 1.124e+11Hz 0.140002 -0.968538
+ 1.125e+11Hz 0.138769 -0.968705
+ 1.126e+11Hz 0.137536 -0.96887
+ 1.127e+11Hz 0.136303 -0.969033
+ 1.128e+11Hz 0.13507 -0.969195
+ 1.129e+11Hz 0.133836 -0.969356
+ 1.13e+11Hz 0.132602 -0.969514
+ 1.131e+11Hz 0.131368 -0.969672
+ 1.132e+11Hz 0.130134 -0.969827
+ 1.133e+11Hz 0.1289 -0.969981
+ 1.134e+11Hz 0.127665 -0.970133
+ 1.135e+11Hz 0.12643 -0.970284
+ 1.136e+11Hz 0.125195 -0.970433
+ 1.137e+11Hz 0.12396 -0.970581
+ 1.138e+11Hz 0.122724 -0.970727
+ 1.139e+11Hz 0.121488 -0.970871
+ 1.14e+11Hz 0.120252 -0.971014
+ 1.141e+11Hz 0.119016 -0.971155
+ 1.142e+11Hz 0.11778 -0.971295
+ 1.143e+11Hz 0.116543 -0.971433
+ 1.144e+11Hz 0.115306 -0.971569
+ 1.145e+11Hz 0.11407 -0.971704
+ 1.146e+11Hz 0.112832 -0.971837
+ 1.147e+11Hz 0.111595 -0.971968
+ 1.148e+11Hz 0.110358 -0.972098
+ 1.149e+11Hz 0.10912 -0.972227
+ 1.15e+11Hz 0.107882 -0.972353
+ 1.151e+11Hz 0.106644 -0.972479
+ 1.152e+11Hz 0.105406 -0.972602
+ 1.153e+11Hz 0.104168 -0.972724
+ 1.154e+11Hz 0.102929 -0.972844
+ 1.155e+11Hz 0.101691 -0.972963
+ 1.156e+11Hz 0.100452 -0.97308
+ 1.157e+11Hz 0.0992128 -0.973196
+ 1.158e+11Hz 0.0979737 -0.973309
+ 1.159e+11Hz 0.0967344 -0.973422
+ 1.16e+11Hz 0.095495 -0.973532
+ 1.161e+11Hz 0.0942555 -0.973641
+ 1.162e+11Hz 0.0930159 -0.973749
+ 1.163e+11Hz 0.0917761 -0.973854
+ 1.164e+11Hz 0.0905362 -0.973959
+ 1.165e+11Hz 0.0892962 -0.974061
+ 1.166e+11Hz 0.088056 -0.974162
+ 1.167e+11Hz 0.0868157 -0.974261
+ 1.168e+11Hz 0.0855754 -0.974359
+ 1.169e+11Hz 0.0843349 -0.974455
+ 1.17e+11Hz 0.0830943 -0.97455
+ 1.171e+11Hz 0.0818536 -0.974642
+ 1.172e+11Hz 0.0806128 -0.974734
+ 1.173e+11Hz 0.0793719 -0.974823
+ 1.174e+11Hz 0.0781309 -0.974911
+ 1.175e+11Hz 0.0768898 -0.974997
+ 1.176e+11Hz 0.0756486 -0.975082
+ 1.177e+11Hz 0.0744074 -0.975165
+ 1.178e+11Hz 0.073166 -0.975247
+ 1.179e+11Hz 0.0719246 -0.975327
+ 1.18e+11Hz 0.0706832 -0.975405
+ 1.181e+11Hz 0.0694416 -0.975482
+ 1.182e+11Hz 0.0682 -0.975557
+ 1.183e+11Hz 0.0669583 -0.97563
+ 1.184e+11Hz 0.0657166 -0.975702
+ 1.185e+11Hz 0.0644748 -0.975772
+ 1.186e+11Hz 0.0632329 -0.975841
+ 1.187e+11Hz 0.061991 -0.975908
+ 1.188e+11Hz 0.0607491 -0.975973
+ 1.189e+11Hz 0.0595071 -0.976037
+ 1.19e+11Hz 0.0582651 -0.976099
+ 1.191e+11Hz 0.057023 -0.976159
+ 1.192e+11Hz 0.055781 -0.976218
+ 1.193e+11Hz 0.0545388 -0.976275
+ 1.194e+11Hz 0.0532967 -0.976331
+ 1.195e+11Hz 0.0520545 -0.976385
+ 1.196e+11Hz 0.0508123 -0.976437
+ 1.197e+11Hz 0.0495702 -0.976488
+ 1.198e+11Hz 0.0483279 -0.976537
+ 1.199e+11Hz 0.0470857 -0.976585
+ 1.2e+11Hz 0.0458435 -0.976631
+ 1.201e+11Hz 0.0446013 -0.976676
+ 1.202e+11Hz 0.043359 -0.976718
+ 1.203e+11Hz 0.0421168 -0.97676
+ 1.204e+11Hz 0.0408746 -0.976799
+ 1.205e+11Hz 0.0396323 -0.976837
+ 1.206e+11Hz 0.0383901 -0.976873
+ 1.207e+11Hz 0.037148 -0.976908
+ 1.208e+11Hz 0.0359058 -0.976942
+ 1.209e+11Hz 0.0346636 -0.976973
+ 1.21e+11Hz 0.0334215 -0.977003
+ 1.211e+11Hz 0.0321794 -0.977032
+ 1.212e+11Hz 0.0309373 -0.977059
+ 1.213e+11Hz 0.0296953 -0.977084
+ 1.214e+11Hz 0.0284533 -0.977108
+ 1.215e+11Hz 0.0272113 -0.97713
+ 1.216e+11Hz 0.0259693 -0.97715
+ 1.217e+11Hz 0.0247275 -0.977169
+ 1.218e+11Hz 0.0234856 -0.977186
+ 1.219e+11Hz 0.0222438 -0.977202
+ 1.22e+11Hz 0.0210021 -0.977216
+ 1.221e+11Hz 0.0197603 -0.977229
+ 1.222e+11Hz 0.0185187 -0.97724
+ 1.223e+11Hz 0.0172771 -0.97725
+ 1.224e+11Hz 0.0160355 -0.977258
+ 1.225e+11Hz 0.0147941 -0.977264
+ 1.226e+11Hz 0.0135526 -0.977269
+ 1.227e+11Hz 0.0123113 -0.977272
+ 1.228e+11Hz 0.01107 -0.977274
+ 1.229e+11Hz 0.00982877 -0.977274
+ 1.23e+11Hz 0.00858762 -0.977272
+ 1.231e+11Hz 0.00734654 -0.977269
+ 1.232e+11Hz 0.00610553 -0.977265
+ 1.233e+11Hz 0.00486459 -0.977259
+ 1.234e+11Hz 0.00362373 -0.977251
+ 1.235e+11Hz 0.00238295 -0.977242
+ 1.236e+11Hz 0.00114225 -0.977231
+ 1.237e+11Hz -9.83727e-05 -0.977219
+ 1.238e+11Hz -0.00133891 -0.977205
+ 1.239e+11Hz -0.00257937 -0.97719
+ 1.24e+11Hz -0.00381974 -0.977173
+ 1.241e+11Hz -0.00506002 -0.977154
+ 1.242e+11Hz -0.00630022 -0.977134
+ 1.243e+11Hz -0.00754032 -0.977113
+ 1.244e+11Hz -0.00878034 -0.97709
+ 1.245e+11Hz -0.0100203 -0.977065
+ 1.246e+11Hz -0.0112601 -0.977039
+ 1.247e+11Hz -0.0124998 -0.977011
+ 1.248e+11Hz -0.0137395 -0.976982
+ 1.249e+11Hz -0.0149791 -0.976951
+ 1.25e+11Hz -0.0162185 -0.976919
+ 1.251e+11Hz -0.0174579 -0.976886
+ 1.252e+11Hz -0.0186971 -0.97685
+ 1.253e+11Hz -0.0199363 -0.976814
+ 1.254e+11Hz -0.0211754 -0.976775
+ 1.255e+11Hz -0.0224143 -0.976735
+ 1.256e+11Hz -0.0236532 -0.976694
+ 1.257e+11Hz -0.024892 -0.976651
+ 1.258e+11Hz -0.0261306 -0.976607
+ 1.259e+11Hz -0.0273692 -0.976561
+ 1.26e+11Hz -0.0286077 -0.976514
+ 1.261e+11Hz -0.029846 -0.976465
+ 1.262e+11Hz -0.0310843 -0.976415
+ 1.263e+11Hz -0.0323225 -0.976363
+ 1.264e+11Hz -0.0335605 -0.97631
+ 1.265e+11Hz -0.0347985 -0.976255
+ 1.266e+11Hz -0.0360364 -0.976198
+ 1.267e+11Hz -0.0372741 -0.976141
+ 1.268e+11Hz -0.0385117 -0.976081
+ 1.269e+11Hz -0.0397493 -0.976021
+ 1.27e+11Hz -0.0409868 -0.975958
+ 1.271e+11Hz -0.0422241 -0.975894
+ 1.272e+11Hz -0.0434613 -0.975829
+ 1.273e+11Hz -0.0446985 -0.975762
+ 1.274e+11Hz -0.0459355 -0.975694
+ 1.275e+11Hz -0.0471724 -0.975624
+ 1.276e+11Hz -0.0484093 -0.975553
+ 1.277e+11Hz -0.049646 -0.97548
+ 1.278e+11Hz -0.0508826 -0.975406
+ 1.279e+11Hz -0.0521192 -0.97533
+ 1.28e+11Hz -0.0533556 -0.975253
+ 1.281e+11Hz -0.0545919 -0.975175
+ 1.282e+11Hz -0.0558281 -0.975094
+ 1.283e+11Hz -0.0570643 -0.975013
+ 1.284e+11Hz -0.0583003 -0.97493
+ 1.285e+11Hz -0.0595362 -0.974845
+ 1.286e+11Hz -0.0607721 -0.974759
+ 1.287e+11Hz -0.0620078 -0.974671
+ 1.288e+11Hz -0.0632434 -0.974582
+ 1.289e+11Hz -0.064479 -0.974491
+ 1.29e+11Hz -0.0657144 -0.974399
+ 1.291e+11Hz -0.0669498 -0.974306
+ 1.292e+11Hz -0.068185 -0.974211
+ 1.293e+11Hz -0.0694202 -0.974114
+ 1.294e+11Hz -0.0706552 -0.974016
+ 1.295e+11Hz -0.0718902 -0.973917
+ 1.296e+11Hz -0.073125 -0.973816
+ 1.297e+11Hz -0.0743598 -0.973713
+ 1.298e+11Hz -0.0755945 -0.973609
+ 1.299e+11Hz -0.0768291 -0.973504
+ 1.3e+11Hz -0.0780636 -0.973397
+ 1.301e+11Hz -0.079298 -0.973289
+ 1.302e+11Hz -0.0805323 -0.973178
+ 1.303e+11Hz -0.0817665 -0.973067
+ 1.304e+11Hz -0.0830006 -0.972954
+ 1.305e+11Hz -0.0842346 -0.97284
+ 1.306e+11Hz -0.0854685 -0.972724
+ 1.307e+11Hz -0.0867024 -0.972606
+ 1.308e+11Hz -0.0879361 -0.972487
+ 1.309e+11Hz -0.0891698 -0.972367
+ 1.31e+11Hz -0.0904033 -0.972245
+ 1.311e+11Hz -0.0916368 -0.972122
+ 1.312e+11Hz -0.0928702 -0.971997
+ 1.313e+11Hz -0.0941035 -0.97187
+ 1.314e+11Hz -0.0953367 -0.971742
+ 1.315e+11Hz -0.0965698 -0.971613
+ 1.316e+11Hz -0.0978028 -0.971482
+ 1.317e+11Hz -0.0990357 -0.971349
+ 1.318e+11Hz -0.100268 -0.971215
+ 1.319e+11Hz -0.101501 -0.97108
+ 1.32e+11Hz -0.102734 -0.970943
+ 1.321e+11Hz -0.103966 -0.970804
+ 1.322e+11Hz -0.105199 -0.970664
+ 1.323e+11Hz -0.106431 -0.970523
+ 1.324e+11Hz -0.107663 -0.970379
+ 1.325e+11Hz -0.108896 -0.970235
+ 1.326e+11Hz -0.110128 -0.970089
+ 1.327e+11Hz -0.11136 -0.969941
+ 1.328e+11Hz -0.112591 -0.969792
+ 1.329e+11Hz -0.113823 -0.969641
+ 1.33e+11Hz -0.115055 -0.969488
+ 1.331e+11Hz -0.116287 -0.969334
+ 1.332e+11Hz -0.117518 -0.969179
+ 1.333e+11Hz -0.118749 -0.969022
+ 1.334e+11Hz -0.119981 -0.968863
+ 1.335e+11Hz -0.121212 -0.968703
+ 1.336e+11Hz -0.122443 -0.968542
+ 1.337e+11Hz -0.123674 -0.968378
+ 1.338e+11Hz -0.124904 -0.968213
+ 1.339e+11Hz -0.126135 -0.968047
+ 1.34e+11Hz -0.127366 -0.967879
+ 1.341e+11Hz -0.128596 -0.96771
+ 1.342e+11Hz -0.129826 -0.967538
+ 1.343e+11Hz -0.131057 -0.967366
+ 1.344e+11Hz -0.132287 -0.967192
+ 1.345e+11Hz -0.133517 -0.967016
+ 1.346e+11Hz -0.134746 -0.966838
+ 1.347e+11Hz -0.135976 -0.966659
+ 1.348e+11Hz -0.137206 -0.966479
+ 1.349e+11Hz -0.138435 -0.966297
+ 1.35e+11Hz -0.139664 -0.966113
+ 1.351e+11Hz -0.140894 -0.965928
+ 1.352e+11Hz -0.142123 -0.965741
+ 1.353e+11Hz -0.143351 -0.965552
+ 1.354e+11Hz -0.14458 -0.965362
+ 1.355e+11Hz -0.145809 -0.96517
+ 1.356e+11Hz -0.147037 -0.964977
+ 1.357e+11Hz -0.148265 -0.964782
+ 1.358e+11Hz -0.149494 -0.964585
+ 1.359e+11Hz -0.150721 -0.964387
+ 1.36e+11Hz -0.151949 -0.964187
+ 1.361e+11Hz -0.153177 -0.963986
+ 1.362e+11Hz -0.154404 -0.963782
+ 1.363e+11Hz -0.155631 -0.963578
+ 1.364e+11Hz -0.156858 -0.963371
+ 1.365e+11Hz -0.158085 -0.963163
+ 1.366e+11Hz -0.159312 -0.962954
+ 1.367e+11Hz -0.160538 -0.962742
+ 1.368e+11Hz -0.161765 -0.96253
+ 1.369e+11Hz -0.162991 -0.962315
+ 1.37e+11Hz -0.164217 -0.962099
+ 1.371e+11Hz -0.165442 -0.961881
+ 1.372e+11Hz -0.166668 -0.961662
+ 1.373e+11Hz -0.167893 -0.961441
+ 1.374e+11Hz -0.169118 -0.961218
+ 1.375e+11Hz -0.170343 -0.960993
+ 1.376e+11Hz -0.171567 -0.960767
+ 1.377e+11Hz -0.172791 -0.96054
+ 1.378e+11Hz -0.174015 -0.96031
+ 1.379e+11Hz -0.175239 -0.960079
+ 1.38e+11Hz -0.176463 -0.959847
+ 1.381e+11Hz -0.177686 -0.959612
+ 1.382e+11Hz -0.178909 -0.959376
+ 1.383e+11Hz -0.180132 -0.959139
+ 1.384e+11Hz -0.181354 -0.958899
+ 1.385e+11Hz -0.182576 -0.958658
+ 1.386e+11Hz -0.183798 -0.958415
+ 1.387e+11Hz -0.18502 -0.958171
+ 1.388e+11Hz -0.186241 -0.957925
+ 1.389e+11Hz -0.187462 -0.957678
+ 1.39e+11Hz -0.188683 -0.957428
+ 1.391e+11Hz -0.189903 -0.957177
+ 1.392e+11Hz -0.191124 -0.956925
+ 1.393e+11Hz -0.192343 -0.95667
+ 1.394e+11Hz -0.193563 -0.956414
+ 1.395e+11Hz -0.194782 -0.956157
+ 1.396e+11Hz -0.196001 -0.955897
+ 1.397e+11Hz -0.197219 -0.955636
+ 1.398e+11Hz -0.198437 -0.955374
+ 1.399e+11Hz -0.199655 -0.95511
+ 1.4e+11Hz -0.200872 -0.954844
+ 1.401e+11Hz -0.202089 -0.954576
+ 1.402e+11Hz -0.203306 -0.954307
+ 1.403e+11Hz -0.204522 -0.954036
+ 1.404e+11Hz -0.205738 -0.953763
+ 1.405e+11Hz -0.206954 -0.953489
+ 1.406e+11Hz -0.208169 -0.953213
+ 1.407e+11Hz -0.209383 -0.952935
+ 1.408e+11Hz -0.210598 -0.952656
+ 1.409e+11Hz -0.211812 -0.952375
+ 1.41e+11Hz -0.213025 -0.952093
+ 1.411e+11Hz -0.214238 -0.951809
+ 1.412e+11Hz -0.215451 -0.951523
+ 1.413e+11Hz -0.216663 -0.951235
+ 1.414e+11Hz -0.217875 -0.950946
+ 1.415e+11Hz -0.219086 -0.950655
+ 1.416e+11Hz -0.220297 -0.950363
+ 1.417e+11Hz -0.221507 -0.950069
+ 1.418e+11Hz -0.222717 -0.949773
+ 1.419e+11Hz -0.223927 -0.949476
+ 1.42e+11Hz -0.225136 -0.949177
+ 1.421e+11Hz -0.226344 -0.948877
+ 1.422e+11Hz -0.227552 -0.948574
+ 1.423e+11Hz -0.22876 -0.948271
+ 1.424e+11Hz -0.229967 -0.947965
+ 1.425e+11Hz -0.231174 -0.947658
+ 1.426e+11Hz -0.23238 -0.94735
+ 1.427e+11Hz -0.233585 -0.94704
+ 1.428e+11Hz -0.23479 -0.946728
+ 1.429e+11Hz -0.235995 -0.946415
+ 1.43e+11Hz -0.237199 -0.946099
+ 1.431e+11Hz -0.238402 -0.945783
+ 1.432e+11Hz -0.239605 -0.945465
+ 1.433e+11Hz -0.240808 -0.945145
+ 1.434e+11Hz -0.24201 -0.944824
+ 1.435e+11Hz -0.243211 -0.944501
+ 1.436e+11Hz -0.244412 -0.944176
+ 1.437e+11Hz -0.245613 -0.943851
+ 1.438e+11Hz -0.246812 -0.943523
+ 1.439e+11Hz -0.248012 -0.943194
+ 1.44e+11Hz -0.24921 -0.942863
+ 1.441e+11Hz -0.250408 -0.942531
+ 1.442e+11Hz -0.251606 -0.942197
+ 1.443e+11Hz -0.252803 -0.941862
+ 1.444e+11Hz -0.253999 -0.941525
+ 1.445e+11Hz -0.255195 -0.941187
+ 1.446e+11Hz -0.256391 -0.940847
+ 1.447e+11Hz -0.257585 -0.940506
+ 1.448e+11Hz -0.25878 -0.940163
+ 1.449e+11Hz -0.259973 -0.939819
+ 1.45e+11Hz -0.261166 -0.939473
+ 1.451e+11Hz -0.262358 -0.939126
+ 1.452e+11Hz -0.26355 -0.938777
+ 1.453e+11Hz -0.264742 -0.938427
+ 1.454e+11Hz -0.265932 -0.938075
+ 1.455e+11Hz -0.267122 -0.937722
+ 1.456e+11Hz -0.268312 -0.937367
+ 1.457e+11Hz -0.269501 -0.937011
+ 1.458e+11Hz -0.270689 -0.936654
+ 1.459e+11Hz -0.271877 -0.936295
+ 1.46e+11Hz -0.273064 -0.935934
+ 1.461e+11Hz -0.27425 -0.935572
+ 1.462e+11Hz -0.275436 -0.935209
+ 1.463e+11Hz -0.276622 -0.934844
+ 1.464e+11Hz -0.277806 -0.934478
+ 1.465e+11Hz -0.27899 -0.934111
+ 1.466e+11Hz -0.280174 -0.933742
+ 1.467e+11Hz -0.281357 -0.933372
+ 1.468e+11Hz -0.282539 -0.933
+ 1.469e+11Hz -0.283721 -0.932627
+ 1.47e+11Hz -0.284902 -0.932252
+ 1.471e+11Hz -0.286083 -0.931876
+ 1.472e+11Hz -0.287263 -0.931499
+ 1.473e+11Hz -0.288442 -0.931121
+ 1.474e+11Hz -0.289621 -0.93074
+ 1.475e+11Hz -0.290799 -0.930359
+ 1.476e+11Hz -0.291977 -0.929976
+ 1.477e+11Hz -0.293154 -0.929593
+ 1.478e+11Hz -0.29433 -0.929207
+ 1.479e+11Hz -0.295507 -0.928821
+ 1.48e+11Hz -0.296682 -0.928432
+ 1.481e+11Hz -0.297857 -0.928043
+ 1.482e+11Hz -0.299031 -0.927652
+ 1.483e+11Hz -0.300204 -0.927261
+ 1.484e+11Hz -0.301378 -0.926867
+ 1.485e+11Hz -0.30255 -0.926473
+ 1.486e+11Hz -0.303722 -0.926077
+ 1.487e+11Hz -0.304894 -0.925679
+ 1.488e+11Hz -0.306065 -0.925281
+ 1.489e+11Hz -0.307235 -0.924881
+ 1.49e+11Hz -0.308405 -0.92448
+ 1.491e+11Hz -0.309574 -0.924078
+ 1.492e+11Hz -0.310743 -0.923674
+ 1.493e+11Hz -0.311911 -0.923269
+ 1.494e+11Hz -0.313079 -0.922863
+ 1.495e+11Hz -0.314246 -0.922455
+ 1.496e+11Hz -0.315412 -0.922047
+ 1.497e+11Hz -0.316579 -0.921637
+ 1.498e+11Hz -0.317744 -0.921225
+ 1.499e+11Hz -0.318909 -0.920813
+ 1.5e+11Hz -0.320074 -0.920399
+ ]

A22 %vd(20 3) %vd(22, 3) xfer4
.model xfer4 xfer R_I=true table=[
+ 0Hz 0.00814086 0
+ 1e+08Hz 0.00814138 1.81109e-05
+ 2e+08Hz 0.00814294 3.62035e-05
+ 3e+08Hz 0.00814553 5.42595e-05
+ 4e+08Hz 0.00814916 7.22604e-05
+ 5e+08Hz 0.00815382 9.01881e-05
+ 6e+08Hz 0.00815952 0.000108024
+ 7e+08Hz 0.00816625 0.000125751
+ 8e+08Hz 0.008174 0.00014335
+ 9e+08Hz 0.00818278 0.000160803
+ 1e+09Hz 0.00819258 0.000178092
+ 1.1e+09Hz 0.0082034 0.000195199
+ 1.2e+09Hz 0.00821522 0.000212108
+ 1.3e+09Hz 0.00822806 0.000228799
+ 1.4e+09Hz 0.0082419 0.000245256
+ 1.5e+09Hz 0.00825673 0.000261462
+ 1.6e+09Hz 0.00827256 0.000277398
+ 1.7e+09Hz 0.00828937 0.000293049
+ 1.8e+09Hz 0.00830716 0.000308397
+ 1.9e+09Hz 0.00832592 0.000323426
+ 2e+09Hz 0.00834564 0.000338119
+ 2.1e+09Hz 0.00836631 0.00035246
+ 2.2e+09Hz 0.00838794 0.000366432
+ 2.3e+09Hz 0.0084105 0.000380021
+ 2.4e+09Hz 0.00843399 0.00039321
+ 2.5e+09Hz 0.0084584 0.000405985
+ 2.6e+09Hz 0.00848372 0.000418329
+ 2.7e+09Hz 0.00850994 0.000430229
+ 2.8e+09Hz 0.00853705 0.00044167
+ 2.9e+09Hz 0.00856504 0.000452636
+ 3e+09Hz 0.0085939 0.000463115
+ 3.1e+09Hz 0.00862361 0.000473093
+ 3.2e+09Hz 0.00865417 0.000482556
+ 3.3e+09Hz 0.00868557 0.00049149
+ 3.4e+09Hz 0.00871779 0.000499884
+ 3.5e+09Hz 0.00875082 0.000507725
+ 3.6e+09Hz 0.00878464 0.000514999
+ 3.7e+09Hz 0.00881925 0.000521697
+ 3.8e+09Hz 0.00885463 0.000527805
+ 3.9e+09Hz 0.00889078 0.000533313
+ 4e+09Hz 0.00892766 0.000538209
+ 4.1e+09Hz 0.00896528 0.000542485
+ 4.2e+09Hz 0.00900361 0.000546128
+ 4.3e+09Hz 0.00904265 0.000549129
+ 4.4e+09Hz 0.00908238 0.000551479
+ 4.5e+09Hz 0.00912278 0.000553169
+ 4.6e+09Hz 0.00916385 0.00055419
+ 4.7e+09Hz 0.00920556 0.000554533
+ 4.8e+09Hz 0.0092479 0.000554191
+ 4.9e+09Hz 0.00929085 0.000553155
+ 5e+09Hz 0.00933441 0.000551419
+ 5.1e+09Hz 0.00937856 0.000548975
+ 5.2e+09Hz 0.00942327 0.000545817
+ 5.3e+09Hz 0.00946854 0.000541939
+ 5.4e+09Hz 0.00951435 0.000537335
+ 5.5e+09Hz 0.00956069 0.000532
+ 5.6e+09Hz 0.00960754 0.000525927
+ 5.7e+09Hz 0.00965488 0.000519114
+ 5.8e+09Hz 0.00970269 0.000511555
+ 5.9e+09Hz 0.00975098 0.000503247
+ 6e+09Hz 0.0097997 0.000494185
+ 6.1e+09Hz 0.00984886 0.000484367
+ 6.2e+09Hz 0.00989844 0.00047379
+ 6.3e+09Hz 0.00994842 0.000462452
+ 6.4e+09Hz 0.00999878 0.000450349
+ 6.5e+09Hz 0.0100495 0.000437481
+ 6.6e+09Hz 0.0101006 0.000423846
+ 6.7e+09Hz 0.010152 0.000409443
+ 6.8e+09Hz 0.0102038 0.000394272
+ 6.9e+09Hz 0.0102558 0.000378331
+ 7e+09Hz 0.0103082 0.000361622
+ 7.1e+09Hz 0.0103608 0.000344143
+ 7.2e+09Hz 0.0104137 0.000325897
+ 7.3e+09Hz 0.0104668 0.000306884
+ 7.4e+09Hz 0.0105202 0.000287105
+ 7.5e+09Hz 0.0105738 0.000266562
+ 7.6e+09Hz 0.0106275 0.000245258
+ 7.7e+09Hz 0.0106815 0.000223193
+ 7.8e+09Hz 0.0107357 0.000200372
+ 7.9e+09Hz 0.01079 0.000176796
+ 8e+09Hz 0.0108445 0.000152469
+ 8.1e+09Hz 0.010899 0.000127395
+ 8.2e+09Hz 0.0109537 0.000101576
+ 8.3e+09Hz 0.0110086 7.50187e-05
+ 8.4e+09Hz 0.0110635 4.77256e-05
+ 8.5e+09Hz 0.0111185 1.97018e-05
+ 8.6e+09Hz 0.0111735 -9.04791e-06
+ 8.7e+09Hz 0.0112286 -3.85183e-05
+ 8.8e+09Hz 0.0112838 -6.87042e-05
+ 8.9e+09Hz 0.0113389 -9.95998e-05
+ 9e+09Hz 0.0113941 -0.000131199
+ 9.1e+09Hz 0.0114493 -0.000163497
+ 9.2e+09Hz 0.0115045 -0.000196486
+ 9.3e+09Hz 0.0115597 -0.00023016
+ 9.4e+09Hz 0.0116148 -0.000264512
+ 9.5e+09Hz 0.0116699 -0.000299536
+ 9.6e+09Hz 0.011725 -0.000335224
+ 9.7e+09Hz 0.01178 -0.000371569
+ 9.8e+09Hz 0.0118349 -0.000408563
+ 9.9e+09Hz 0.0118897 -0.0004462
+ 1e+10Hz 0.0119444 -0.00048447
+ 1.01e+10Hz 0.0119991 -0.000523366
+ 1.02e+10Hz 0.0120536 -0.000562881
+ 1.03e+10Hz 0.012108 -0.000603005
+ 1.04e+10Hz 0.0121622 -0.00064373
+ 1.05e+10Hz 0.0122164 -0.000685048
+ 1.06e+10Hz 0.0122703 -0.00072695
+ 1.07e+10Hz 0.0123242 -0.000769427
+ 1.08e+10Hz 0.0123778 -0.00081247
+ 1.09e+10Hz 0.0124314 -0.000856071
+ 1.1e+10Hz 0.0124847 -0.00090022
+ 1.11e+10Hz 0.0125378 -0.000944909
+ 1.12e+10Hz 0.0125907 -0.000990126
+ 1.13e+10Hz 0.0126435 -0.00103586
+ 1.14e+10Hz 0.012696 -0.00108212
+ 1.15e+10Hz 0.0127484 -0.00112887
+ 1.16e+10Hz 0.0128005 -0.00117611
+ 1.17e+10Hz 0.0128524 -0.00122384
+ 1.18e+10Hz 0.0129041 -0.00127203
+ 1.19e+10Hz 0.0129555 -0.0013207
+ 1.2e+10Hz 0.0130067 -0.00136981
+ 1.21e+10Hz 0.0130577 -0.00141937
+ 1.22e+10Hz 0.0131084 -0.00146937
+ 1.23e+10Hz 0.0131589 -0.00151979
+ 1.24e+10Hz 0.0132091 -0.00157062
+ 1.25e+10Hz 0.0132591 -0.00162186
+ 1.26e+10Hz 0.0133088 -0.0016735
+ 1.27e+10Hz 0.0133582 -0.00172552
+ 1.28e+10Hz 0.0134074 -0.00177791
+ 1.29e+10Hz 0.0134563 -0.00183068
+ 1.3e+10Hz 0.013505 -0.0018838
+ 1.31e+10Hz 0.0135533 -0.00193727
+ 1.32e+10Hz 0.0136014 -0.00199108
+ 1.33e+10Hz 0.0136493 -0.00204521
+ 1.34e+10Hz 0.0136968 -0.00209967
+ 1.35e+10Hz 0.0137441 -0.00215443
+ 1.36e+10Hz 0.0137911 -0.0022095
+ 1.37e+10Hz 0.0138379 -0.00226486
+ 1.38e+10Hz 0.0138843 -0.00232049
+ 1.39e+10Hz 0.0139305 -0.00237641
+ 1.4e+10Hz 0.0139764 -0.00243258
+ 1.41e+10Hz 0.014022 -0.00248901
+ 1.42e+10Hz 0.0140673 -0.00254569
+ 1.43e+10Hz 0.0141124 -0.00260261
+ 1.44e+10Hz 0.0141572 -0.00265976
+ 1.45e+10Hz 0.0142017 -0.00271712
+ 1.46e+10Hz 0.0142459 -0.0027747
+ 1.47e+10Hz 0.0142899 -0.00283249
+ 1.48e+10Hz 0.0143336 -0.00289047
+ 1.49e+10Hz 0.014377 -0.00294863
+ 1.5e+10Hz 0.0144202 -0.00300698
+ 1.51e+10Hz 0.0144631 -0.0030655
+ 1.52e+10Hz 0.0145057 -0.00312418
+ 1.53e+10Hz 0.0145481 -0.00318303
+ 1.54e+10Hz 0.0145902 -0.00324202
+ 1.55e+10Hz 0.0146321 -0.00330115
+ 1.56e+10Hz 0.0146737 -0.00336042
+ 1.57e+10Hz 0.014715 -0.00341982
+ 1.58e+10Hz 0.0147561 -0.00347933
+ 1.59e+10Hz 0.014797 -0.00353896
+ 1.6e+10Hz 0.0148376 -0.0035987
+ 1.61e+10Hz 0.014878 -0.00365855
+ 1.62e+10Hz 0.0149182 -0.00371848
+ 1.63e+10Hz 0.0149581 -0.00377851
+ 1.64e+10Hz 0.0149978 -0.00383862
+ 1.65e+10Hz 0.0150373 -0.0038988
+ 1.66e+10Hz 0.0150765 -0.00395906
+ 1.67e+10Hz 0.0151156 -0.00401939
+ 1.68e+10Hz 0.0151544 -0.00407977
+ 1.69e+10Hz 0.0151931 -0.00414021
+ 1.7e+10Hz 0.0152315 -0.0042007
+ 1.71e+10Hz 0.0152698 -0.00426123
+ 1.72e+10Hz 0.0153078 -0.00432181
+ 1.73e+10Hz 0.0153457 -0.00438242
+ 1.74e+10Hz 0.0153834 -0.00444307
+ 1.75e+10Hz 0.0154208 -0.00450374
+ 1.76e+10Hz 0.0154582 -0.00456443
+ 1.77e+10Hz 0.0154953 -0.00462514
+ 1.78e+10Hz 0.0155323 -0.00468587
+ 1.79e+10Hz 0.0155692 -0.00474661
+ 1.8e+10Hz 0.0156058 -0.00480736
+ 1.81e+10Hz 0.0156424 -0.00486811
+ 1.82e+10Hz 0.0156788 -0.00492887
+ 1.83e+10Hz 0.015715 -0.00498962
+ 1.84e+10Hz 0.0157511 -0.00505037
+ 1.85e+10Hz 0.0157871 -0.00511111
+ 1.86e+10Hz 0.015823 -0.00517184
+ 1.87e+10Hz 0.0158587 -0.00523256
+ 1.88e+10Hz 0.0158944 -0.00529327
+ 1.89e+10Hz 0.0159299 -0.00535395
+ 1.9e+10Hz 0.0159653 -0.00541463
+ 1.91e+10Hz 0.0160006 -0.00547528
+ 1.92e+10Hz 0.0160359 -0.0055359
+ 1.93e+10Hz 0.016071 -0.00559651
+ 1.94e+10Hz 0.0161061 -0.00565709
+ 1.95e+10Hz 0.016141 -0.00571764
+ 1.96e+10Hz 0.0161759 -0.00577817
+ 1.97e+10Hz 0.0162108 -0.00583867
+ 1.98e+10Hz 0.0162455 -0.00589914
+ 1.99e+10Hz 0.0162802 -0.00595958
+ 2e+10Hz 0.0163149 -0.00601999
+ 2.01e+10Hz 0.0163495 -0.00608036
+ 2.02e+10Hz 0.0163841 -0.00614071
+ 2.03e+10Hz 0.0164186 -0.00620102
+ 2.04e+10Hz 0.0164531 -0.00626131
+ 2.05e+10Hz 0.0164875 -0.00632156
+ 2.06e+10Hz 0.016522 -0.00638178
+ 2.07e+10Hz 0.0165564 -0.00644197
+ 2.08e+10Hz 0.0165908 -0.00650213
+ 2.09e+10Hz 0.0166252 -0.00656226
+ 2.1e+10Hz 0.0166595 -0.00662236
+ 2.11e+10Hz 0.0166939 -0.00668243
+ 2.12e+10Hz 0.0167283 -0.00674247
+ 2.13e+10Hz 0.0167627 -0.00680248
+ 2.14e+10Hz 0.016797 -0.00686247
+ 2.15e+10Hz 0.0168314 -0.00692244
+ 2.16e+10Hz 0.0168659 -0.00698237
+ 2.17e+10Hz 0.0169003 -0.00704229
+ 2.18e+10Hz 0.0169347 -0.00710219
+ 2.19e+10Hz 0.0169692 -0.00716206
+ 2.2e+10Hz 0.0170038 -0.00722192
+ 2.21e+10Hz 0.0170383 -0.00728176
+ 2.22e+10Hz 0.0170729 -0.00734159
+ 2.23e+10Hz 0.0171076 -0.0074014
+ 2.24e+10Hz 0.0171422 -0.00746121
+ 2.25e+10Hz 0.017177 -0.007521
+ 2.26e+10Hz 0.0172118 -0.00758079
+ 2.27e+10Hz 0.0172466 -0.00764057
+ 2.28e+10Hz 0.0172815 -0.00770035
+ 2.29e+10Hz 0.0173165 -0.00776013
+ 2.3e+10Hz 0.0173515 -0.00781991
+ 2.31e+10Hz 0.0173866 -0.00787969
+ 2.32e+10Hz 0.0174218 -0.00793948
+ 2.33e+10Hz 0.017457 -0.00799928
+ 2.34e+10Hz 0.0174923 -0.00805909
+ 2.35e+10Hz 0.0175277 -0.00811891
+ 2.36e+10Hz 0.0175632 -0.00817875
+ 2.37e+10Hz 0.0175988 -0.0082386
+ 2.38e+10Hz 0.0176344 -0.00829848
+ 2.39e+10Hz 0.0176701 -0.00835838
+ 2.4e+10Hz 0.017706 -0.00841832
+ 2.41e+10Hz 0.0177419 -0.00847827
+ 2.42e+10Hz 0.0177779 -0.00853826
+ 2.43e+10Hz 0.017814 -0.00859829
+ 2.44e+10Hz 0.0178501 -0.00865835
+ 2.45e+10Hz 0.0178864 -0.00871846
+ 2.46e+10Hz 0.0179228 -0.0087786
+ 2.47e+10Hz 0.0179593 -0.0088388
+ 2.48e+10Hz 0.0179959 -0.00889904
+ 2.49e+10Hz 0.0180326 -0.00895933
+ 2.5e+10Hz 0.0180694 -0.00901968
+ 2.51e+10Hz 0.0181063 -0.00908008
+ 2.52e+10Hz 0.0181433 -0.00914055
+ 2.53e+10Hz 0.0181804 -0.00920108
+ 2.54e+10Hz 0.0182176 -0.00926168
+ 2.55e+10Hz 0.0182549 -0.00932234
+ 2.56e+10Hz 0.0182924 -0.00938308
+ 2.57e+10Hz 0.0183299 -0.00944389
+ 2.58e+10Hz 0.0183675 -0.00950478
+ 2.59e+10Hz 0.0184053 -0.00956575
+ 2.6e+10Hz 0.0184432 -0.0096268
+ 2.61e+10Hz 0.0184812 -0.00968794
+ 2.62e+10Hz 0.0185193 -0.00974917
+ 2.63e+10Hz 0.0185575 -0.00981049
+ 2.64e+10Hz 0.0185958 -0.0098719
+ 2.65e+10Hz 0.0186342 -0.00993341
+ 2.66e+10Hz 0.0186727 -0.00999502
+ 2.67e+10Hz 0.0187114 -0.0100567
+ 2.68e+10Hz 0.0187501 -0.0101186
+ 2.69e+10Hz 0.018789 -0.0101805
+ 2.7e+10Hz 0.0188279 -0.0102425
+ 2.71e+10Hz 0.018867 -0.0103047
+ 2.72e+10Hz 0.0189062 -0.0103669
+ 2.73e+10Hz 0.0189455 -0.0104293
+ 2.74e+10Hz 0.0189849 -0.0104918
+ 2.75e+10Hz 0.0190244 -0.0105544
+ 2.76e+10Hz 0.019064 -0.0106172
+ 2.77e+10Hz 0.0191037 -0.0106801
+ 2.78e+10Hz 0.0191435 -0.0107431
+ 2.79e+10Hz 0.0191835 -0.0108062
+ 2.8e+10Hz 0.0192235 -0.0108695
+ 2.81e+10Hz 0.0192636 -0.0109329
+ 2.82e+10Hz 0.0193038 -0.0109965
+ 2.83e+10Hz 0.0193441 -0.0110602
+ 2.84e+10Hz 0.0193845 -0.011124
+ 2.85e+10Hz 0.019425 -0.011188
+ 2.86e+10Hz 0.0194657 -0.0112521
+ 2.87e+10Hz 0.0195063 -0.0113164
+ 2.88e+10Hz 0.0195471 -0.0113808
+ 2.89e+10Hz 0.019588 -0.0114454
+ 2.9e+10Hz 0.019629 -0.0115101
+ 2.91e+10Hz 0.01967 -0.011575
+ 2.92e+10Hz 0.0197111 -0.0116401
+ 2.93e+10Hz 0.0197523 -0.0117053
+ 2.94e+10Hz 0.0197936 -0.0117707
+ 2.95e+10Hz 0.019835 -0.0118362
+ 2.96e+10Hz 0.0198765 -0.0119019
+ 2.97e+10Hz 0.019918 -0.0119678
+ 2.98e+10Hz 0.0199596 -0.0120338
+ 2.99e+10Hz 0.0200013 -0.0121
+ 3e+10Hz 0.0200431 -0.0121664
+ 3.01e+10Hz 0.0200849 -0.0122329
+ 3.02e+10Hz 0.0201268 -0.0122996
+ 3.03e+10Hz 0.0201688 -0.0123665
+ 3.04e+10Hz 0.0202108 -0.0124336
+ 3.05e+10Hz 0.0202529 -0.0125008
+ 3.06e+10Hz 0.020295 -0.0125682
+ 3.07e+10Hz 0.0203372 -0.0126358
+ 3.08e+10Hz 0.0203795 -0.0127036
+ 3.09e+10Hz 0.0204218 -0.0127715
+ 3.1e+10Hz 0.0204642 -0.0128397
+ 3.11e+10Hz 0.0205066 -0.012908
+ 3.12e+10Hz 0.0205491 -0.0129765
+ 3.13e+10Hz 0.0205916 -0.0130451
+ 3.14e+10Hz 0.0206342 -0.013114
+ 3.15e+10Hz 0.0206768 -0.013183
+ 3.16e+10Hz 0.0207195 -0.0132522
+ 3.17e+10Hz 0.0207622 -0.0133216
+ 3.18e+10Hz 0.0208049 -0.0133912
+ 3.19e+10Hz 0.0208477 -0.013461
+ 3.2e+10Hz 0.0208905 -0.0135309
+ 3.21e+10Hz 0.0209333 -0.0136011
+ 3.22e+10Hz 0.0209762 -0.0136714
+ 3.23e+10Hz 0.0210191 -0.0137419
+ 3.24e+10Hz 0.021062 -0.0138126
+ 3.25e+10Hz 0.021105 -0.0138835
+ 3.26e+10Hz 0.0211479 -0.0139546
+ 3.27e+10Hz 0.0211909 -0.0140258
+ 3.28e+10Hz 0.021234 -0.0140973
+ 3.29e+10Hz 0.021277 -0.0141689
+ 3.3e+10Hz 0.0213201 -0.0142407
+ 3.31e+10Hz 0.0213631 -0.0143127
+ 3.32e+10Hz 0.0214062 -0.0143849
+ 3.33e+10Hz 0.0214493 -0.0144572
+ 3.34e+10Hz 0.0214924 -0.0145298
+ 3.35e+10Hz 0.0215355 -0.0146025
+ 3.36e+10Hz 0.0215786 -0.0146754
+ 3.37e+10Hz 0.0216218 -0.0147485
+ 3.38e+10Hz 0.0216649 -0.0148218
+ 3.39e+10Hz 0.021708 -0.0148953
+ 3.4e+10Hz 0.0217511 -0.0149689
+ 3.41e+10Hz 0.0217943 -0.0150428
+ 3.42e+10Hz 0.0218374 -0.0151168
+ 3.43e+10Hz 0.0218805 -0.015191
+ 3.44e+10Hz 0.0219236 -0.0152653
+ 3.45e+10Hz 0.0219667 -0.0153399
+ 3.46e+10Hz 0.0220098 -0.0154146
+ 3.47e+10Hz 0.0220529 -0.0154895
+ 3.48e+10Hz 0.022096 -0.0155646
+ 3.49e+10Hz 0.0221391 -0.0156399
+ 3.5e+10Hz 0.0221821 -0.0157153
+ 3.51e+10Hz 0.0222251 -0.0157909
+ 3.52e+10Hz 0.0222682 -0.0158667
+ 3.53e+10Hz 0.0223112 -0.0159426
+ 3.54e+10Hz 0.0223541 -0.0160188
+ 3.55e+10Hz 0.0223971 -0.0160951
+ 3.56e+10Hz 0.02244 -0.0161715
+ 3.57e+10Hz 0.022483 -0.0162482
+ 3.58e+10Hz 0.0225259 -0.016325
+ 3.59e+10Hz 0.0225687 -0.016402
+ 3.6e+10Hz 0.0226116 -0.0164791
+ 3.61e+10Hz 0.0226544 -0.0165564
+ 3.62e+10Hz 0.0226972 -0.0166339
+ 3.63e+10Hz 0.02274 -0.0167115
+ 3.64e+10Hz 0.0227827 -0.0167893
+ 3.65e+10Hz 0.0228254 -0.0168673
+ 3.66e+10Hz 0.0228681 -0.0169454
+ 3.67e+10Hz 0.0229107 -0.0170237
+ 3.68e+10Hz 0.0229534 -0.0171021
+ 3.69e+10Hz 0.0229959 -0.0171808
+ 3.7e+10Hz 0.0230385 -0.0172595
+ 3.71e+10Hz 0.023081 -0.0173384
+ 3.72e+10Hz 0.0231235 -0.0174175
+ 3.73e+10Hz 0.0231659 -0.0174967
+ 3.74e+10Hz 0.0232083 -0.0175761
+ 3.75e+10Hz 0.0232507 -0.0176556
+ 3.76e+10Hz 0.023293 -0.0177353
+ 3.77e+10Hz 0.0233354 -0.0178151
+ 3.78e+10Hz 0.0233776 -0.0178951
+ 3.79e+10Hz 0.0234198 -0.0179753
+ 3.8e+10Hz 0.023462 -0.0180555
+ 3.81e+10Hz 0.0235042 -0.018136
+ 3.82e+10Hz 0.0235463 -0.0182165
+ 3.83e+10Hz 0.0235884 -0.0182972
+ 3.84e+10Hz 0.0236304 -0.0183781
+ 3.85e+10Hz 0.0236724 -0.0184591
+ 3.86e+10Hz 0.0237143 -0.0185402
+ 3.87e+10Hz 0.0237562 -0.0186215
+ 3.88e+10Hz 0.0237981 -0.0187029
+ 3.89e+10Hz 0.0238399 -0.0187845
+ 3.9e+10Hz 0.0238817 -0.0188662
+ 3.91e+10Hz 0.0239235 -0.018948
+ 3.92e+10Hz 0.0239652 -0.01903
+ 3.93e+10Hz 0.0240069 -0.0191121
+ 3.94e+10Hz 0.0240485 -0.0191943
+ 3.95e+10Hz 0.0240901 -0.0192767
+ 3.96e+10Hz 0.0241316 -0.0193592
+ 3.97e+10Hz 0.0241731 -0.0194418
+ 3.98e+10Hz 0.0242146 -0.0195246
+ 3.99e+10Hz 0.024256 -0.0196075
+ 4e+10Hz 0.0242974 -0.0196905
+ 4.01e+10Hz 0.0243387 -0.0197737
+ 4.02e+10Hz 0.02438 -0.0198569
+ 4.03e+10Hz 0.0244213 -0.0199403
+ 4.04e+10Hz 0.0244625 -0.0200239
+ 4.05e+10Hz 0.0245037 -0.0201075
+ 4.06e+10Hz 0.0245449 -0.0201913
+ 4.07e+10Hz 0.024586 -0.0202752
+ 4.08e+10Hz 0.024627 -0.0203593
+ 4.09e+10Hz 0.0246681 -0.0204434
+ 4.1e+10Hz 0.024709 -0.0205277
+ 4.11e+10Hz 0.02475 -0.0206121
+ 4.12e+10Hz 0.0247909 -0.0206966
+ 4.13e+10Hz 0.0248318 -0.0207813
+ 4.14e+10Hz 0.0248726 -0.020866
+ 4.15e+10Hz 0.0249134 -0.0209509
+ 4.16e+10Hz 0.0249542 -0.0210359
+ 4.17e+10Hz 0.0249949 -0.021121
+ 4.18e+10Hz 0.0250356 -0.0212063
+ 4.19e+10Hz 0.0250763 -0.0212916
+ 4.2e+10Hz 0.0251169 -0.0213771
+ 4.21e+10Hz 0.0251575 -0.0214627
+ 4.22e+10Hz 0.025198 -0.0215484
+ 4.23e+10Hz 0.0252385 -0.0216342
+ 4.24e+10Hz 0.025279 -0.0217202
+ 4.25e+10Hz 0.0253195 -0.0218062
+ 4.26e+10Hz 0.0253599 -0.0218924
+ 4.27e+10Hz 0.0254003 -0.0219787
+ 4.28e+10Hz 0.0254406 -0.0220651
+ 4.29e+10Hz 0.0254809 -0.0221516
+ 4.3e+10Hz 0.0255212 -0.0222383
+ 4.31e+10Hz 0.0255615 -0.022325
+ 4.32e+10Hz 0.0256017 -0.0224119
+ 4.33e+10Hz 0.0256419 -0.0224989
+ 4.34e+10Hz 0.0256821 -0.022586
+ 4.35e+10Hz 0.0257222 -0.0226732
+ 4.36e+10Hz 0.0257623 -0.0227605
+ 4.37e+10Hz 0.0258024 -0.0228479
+ 4.38e+10Hz 0.0258425 -0.0229355
+ 4.39e+10Hz 0.0258825 -0.0230231
+ 4.4e+10Hz 0.0259225 -0.0231109
+ 4.41e+10Hz 0.0259625 -0.0231988
+ 4.42e+10Hz 0.0260024 -0.0232868
+ 4.43e+10Hz 0.0260423 -0.023375
+ 4.44e+10Hz 0.0260822 -0.0234632
+ 4.45e+10Hz 0.0261221 -0.0235516
+ 4.46e+10Hz 0.0261619 -0.02364
+ 4.47e+10Hz 0.0262017 -0.0237286
+ 4.48e+10Hz 0.0262415 -0.0238173
+ 4.49e+10Hz 0.0262813 -0.0239061
+ 4.5e+10Hz 0.026321 -0.0239951
+ 4.51e+10Hz 0.0263607 -0.0240841
+ 4.52e+10Hz 0.0264004 -0.0241733
+ 4.53e+10Hz 0.0264401 -0.0242626
+ 4.54e+10Hz 0.0264797 -0.024352
+ 4.55e+10Hz 0.0265194 -0.0244415
+ 4.56e+10Hz 0.026559 -0.0245311
+ 4.57e+10Hz 0.0265985 -0.0246209
+ 4.58e+10Hz 0.0266381 -0.0247107
+ 4.59e+10Hz 0.0266776 -0.0248007
+ 4.6e+10Hz 0.0267171 -0.0248908
+ 4.61e+10Hz 0.0267566 -0.024981
+ 4.62e+10Hz 0.0267961 -0.0250714
+ 4.63e+10Hz 0.0268355 -0.0251618
+ 4.64e+10Hz 0.0268749 -0.0252524
+ 4.65e+10Hz 0.0269143 -0.0253431
+ 4.66e+10Hz 0.0269537 -0.025434
+ 4.67e+10Hz 0.0269931 -0.0255249
+ 4.68e+10Hz 0.0270324 -0.025616
+ 4.69e+10Hz 0.0270717 -0.0257072
+ 4.7e+10Hz 0.027111 -0.0257985
+ 4.71e+10Hz 0.0271503 -0.0258899
+ 4.72e+10Hz 0.0271895 -0.0259815
+ 4.73e+10Hz 0.0272288 -0.0260732
+ 4.74e+10Hz 0.027268 -0.026165
+ 4.75e+10Hz 0.0273072 -0.0262569
+ 4.76e+10Hz 0.0273463 -0.026349
+ 4.77e+10Hz 0.0273855 -0.0264412
+ 4.78e+10Hz 0.0274246 -0.0265335
+ 4.79e+10Hz 0.0274637 -0.0266259
+ 4.8e+10Hz 0.0275028 -0.0267185
+ 4.81e+10Hz 0.0275419 -0.0268112
+ 4.82e+10Hz 0.0275809 -0.026904
+ 4.83e+10Hz 0.0276199 -0.026997
+ 4.84e+10Hz 0.0276589 -0.0270901
+ 4.85e+10Hz 0.0276979 -0.0271833
+ 4.86e+10Hz 0.0277368 -0.0272767
+ 4.87e+10Hz 0.0277757 -0.0273702
+ 4.88e+10Hz 0.0278146 -0.0274638
+ 4.89e+10Hz 0.0278535 -0.0275575
+ 4.9e+10Hz 0.0278924 -0.0276514
+ 4.91e+10Hz 0.0279312 -0.0277454
+ 4.92e+10Hz 0.02797 -0.0278396
+ 4.93e+10Hz 0.0280088 -0.0279339
+ 4.94e+10Hz 0.0280475 -0.0280283
+ 4.95e+10Hz 0.0280862 -0.0281228
+ 4.96e+10Hz 0.0281249 -0.0282175
+ 4.97e+10Hz 0.0281636 -0.0283124
+ 4.98e+10Hz 0.0282023 -0.0284073
+ 4.99e+10Hz 0.0282409 -0.0285024
+ 5e+10Hz 0.0282795 -0.0285977
+ 5.01e+10Hz 0.028318 -0.0286931
+ 5.02e+10Hz 0.0283566 -0.0287886
+ 5.03e+10Hz 0.028395 -0.0288843
+ 5.04e+10Hz 0.0284335 -0.0289801
+ 5.05e+10Hz 0.0284719 -0.029076
+ 5.06e+10Hz 0.0285104 -0.0291721
+ 5.07e+10Hz 0.0285487 -0.0292683
+ 5.08e+10Hz 0.0285871 -0.0293647
+ 5.09e+10Hz 0.0286254 -0.0294612
+ 5.1e+10Hz 0.0286637 -0.0295579
+ 5.11e+10Hz 0.0287019 -0.0296547
+ 5.12e+10Hz 0.0287401 -0.0297517
+ 5.13e+10Hz 0.0287783 -0.0298488
+ 5.14e+10Hz 0.0288164 -0.029946
+ 5.15e+10Hz 0.0288545 -0.0300434
+ 5.16e+10Hz 0.0288925 -0.0301409
+ 5.17e+10Hz 0.0289306 -0.0302386
+ 5.18e+10Hz 0.0289685 -0.0303364
+ 5.19e+10Hz 0.0290065 -0.0304344
+ 5.2e+10Hz 0.0290444 -0.0305325
+ 5.21e+10Hz 0.0290822 -0.0306308
+ 5.22e+10Hz 0.0291201 -0.0307292
+ 5.23e+10Hz 0.0291578 -0.0308278
+ 5.24e+10Hz 0.0291955 -0.0309265
+ 5.25e+10Hz 0.0292332 -0.0310253
+ 5.26e+10Hz 0.0292709 -0.0311243
+ 5.27e+10Hz 0.0293084 -0.0312235
+ 5.28e+10Hz 0.029346 -0.0313228
+ 5.29e+10Hz 0.0293835 -0.0314223
+ 5.3e+10Hz 0.0294209 -0.0315219
+ 5.31e+10Hz 0.0294583 -0.0316216
+ 5.32e+10Hz 0.0294957 -0.0317215
+ 5.33e+10Hz 0.0295329 -0.0318216
+ 5.34e+10Hz 0.0295702 -0.0319218
+ 5.35e+10Hz 0.0296074 -0.0320222
+ 5.36e+10Hz 0.0296445 -0.0321227
+ 5.37e+10Hz 0.0296816 -0.0322234
+ 5.38e+10Hz 0.0297186 -0.0323242
+ 5.39e+10Hz 0.0297555 -0.0324251
+ 5.4e+10Hz 0.0297924 -0.0325263
+ 5.41e+10Hz 0.0298293 -0.0326275
+ 5.42e+10Hz 0.0298661 -0.032729
+ 5.43e+10Hz 0.0299028 -0.0328305
+ 5.44e+10Hz 0.0299394 -0.0329323
+ 5.45e+10Hz 0.029976 -0.0330341
+ 5.46e+10Hz 0.0300126 -0.0331362
+ 5.47e+10Hz 0.030049 -0.0332383
+ 5.48e+10Hz 0.0300854 -0.0333407
+ 5.49e+10Hz 0.0301218 -0.0334432
+ 5.5e+10Hz 0.030158 -0.0335458
+ 5.51e+10Hz 0.0301942 -0.0336486
+ 5.52e+10Hz 0.0302304 -0.0337515
+ 5.53e+10Hz 0.0302664 -0.0338546
+ 5.54e+10Hz 0.0303024 -0.0339579
+ 5.55e+10Hz 0.0303384 -0.0340613
+ 5.56e+10Hz 0.0303742 -0.0341648
+ 5.57e+10Hz 0.03041 -0.0342685
+ 5.58e+10Hz 0.0304457 -0.0343723
+ 5.59e+10Hz 0.0304813 -0.0344763
+ 5.6e+10Hz 0.0305168 -0.0345805
+ 5.61e+10Hz 0.0305523 -0.0346848
+ 5.62e+10Hz 0.0305877 -0.0347892
+ 5.63e+10Hz 0.030623 -0.0348938
+ 5.64e+10Hz 0.0306582 -0.0349986
+ 5.65e+10Hz 0.0306934 -0.0351034
+ 5.66e+10Hz 0.0307284 -0.0352085
+ 5.67e+10Hz 0.0307634 -0.0353137
+ 5.68e+10Hz 0.0307983 -0.035419
+ 5.69e+10Hz 0.0308331 -0.0355245
+ 5.7e+10Hz 0.0308678 -0.0356301
+ 5.71e+10Hz 0.0309025 -0.0357359
+ 5.72e+10Hz 0.030937 -0.0358418
+ 5.73e+10Hz 0.0309715 -0.0359479
+ 5.74e+10Hz 0.0310059 -0.0360541
+ 5.75e+10Hz 0.0310402 -0.0361604
+ 5.76e+10Hz 0.0310744 -0.0362669
+ 5.77e+10Hz 0.0311085 -0.0363736
+ 5.78e+10Hz 0.0311425 -0.0364804
+ 5.79e+10Hz 0.0311764 -0.0365873
+ 5.8e+10Hz 0.0312102 -0.0366944
+ 5.81e+10Hz 0.0312439 -0.0368016
+ 5.82e+10Hz 0.0312776 -0.036909
+ 5.83e+10Hz 0.0313111 -0.0370165
+ 5.84e+10Hz 0.0313446 -0.0371241
+ 5.85e+10Hz 0.0313779 -0.0372319
+ 5.86e+10Hz 0.0314111 -0.0373398
+ 5.87e+10Hz 0.0314443 -0.0374479
+ 5.88e+10Hz 0.0314773 -0.0375561
+ 5.89e+10Hz 0.0315103 -0.0376644
+ 5.9e+10Hz 0.0315431 -0.0377729
+ 5.91e+10Hz 0.0315759 -0.0378815
+ 5.92e+10Hz 0.0316085 -0.0379903
+ 5.93e+10Hz 0.031641 -0.0380992
+ 5.94e+10Hz 0.0316734 -0.0382082
+ 5.95e+10Hz 0.0317058 -0.0383174
+ 5.96e+10Hz 0.031738 -0.0384266
+ 5.97e+10Hz 0.0317701 -0.0385361
+ 5.98e+10Hz 0.0318021 -0.0386456
+ 5.99e+10Hz 0.031834 -0.0387553
+ 6e+10Hz 0.0318658 -0.0388651
+ 6.01e+10Hz 0.0318974 -0.0389751
+ 6.02e+10Hz 0.031929 -0.0390852
+ 6.03e+10Hz 0.0319605 -0.0391954
+ 6.04e+10Hz 0.0319918 -0.0393057
+ 6.05e+10Hz 0.032023 -0.0394162
+ 6.06e+10Hz 0.0320542 -0.0395268
+ 6.07e+10Hz 0.0320852 -0.0396375
+ 6.08e+10Hz 0.0321161 -0.0397484
+ 6.09e+10Hz 0.0321469 -0.0398594
+ 6.1e+10Hz 0.0321775 -0.0399705
+ 6.11e+10Hz 0.0322081 -0.0400817
+ 6.12e+10Hz 0.0322385 -0.0401931
+ 6.13e+10Hz 0.0322689 -0.0403045
+ 6.14e+10Hz 0.0322991 -0.0404161
+ 6.15e+10Hz 0.0323292 -0.0405278
+ 6.16e+10Hz 0.0323592 -0.0406397
+ 6.17e+10Hz 0.032389 -0.0407517
+ 6.18e+10Hz 0.0324188 -0.0408637
+ 6.19e+10Hz 0.0324484 -0.0409759
+ 6.2e+10Hz 0.0324779 -0.0410883
+ 6.21e+10Hz 0.0325073 -0.0412007
+ 6.22e+10Hz 0.0325366 -0.0413133
+ 6.23e+10Hz 0.0325657 -0.0414259
+ 6.24e+10Hz 0.0325948 -0.0415387
+ 6.25e+10Hz 0.0326237 -0.0416516
+ 6.26e+10Hz 0.0326525 -0.0417647
+ 6.27e+10Hz 0.0326812 -0.0418778
+ 6.28e+10Hz 0.0327097 -0.041991
+ 6.29e+10Hz 0.0327382 -0.0421044
+ 6.3e+10Hz 0.0327665 -0.0422179
+ 6.31e+10Hz 0.0327947 -0.0423314
+ 6.32e+10Hz 0.0328227 -0.0424451
+ 6.33e+10Hz 0.0328507 -0.0425589
+ 6.34e+10Hz 0.0328785 -0.0426729
+ 6.35e+10Hz 0.0329062 -0.0427869
+ 6.36e+10Hz 0.0329338 -0.042901
+ 6.37e+10Hz 0.0329612 -0.0430152
+ 6.38e+10Hz 0.0329885 -0.0431296
+ 6.39e+10Hz 0.0330158 -0.043244
+ 6.4e+10Hz 0.0330428 -0.0433586
+ 6.41e+10Hz 0.0330698 -0.0434733
+ 6.42e+10Hz 0.0330966 -0.043588
+ 6.43e+10Hz 0.0331234 -0.0437029
+ 6.44e+10Hz 0.0331499 -0.0438179
+ 6.45e+10Hz 0.0331764 -0.043933
+ 6.46e+10Hz 0.0332028 -0.0440482
+ 6.47e+10Hz 0.033229 -0.0441634
+ 6.48e+10Hz 0.0332551 -0.0442788
+ 6.49e+10Hz 0.033281 -0.0443943
+ 6.5e+10Hz 0.0333069 -0.0445099
+ 6.51e+10Hz 0.0333326 -0.0446256
+ 6.52e+10Hz 0.0333582 -0.0447414
+ 6.53e+10Hz 0.0333836 -0.0448573
+ 6.54e+10Hz 0.033409 -0.0449732
+ 6.55e+10Hz 0.0334342 -0.0450893
+ 6.56e+10Hz 0.0334593 -0.0452055
+ 6.57e+10Hz 0.0334842 -0.0453218
+ 6.58e+10Hz 0.0335091 -0.0454381
+ 6.59e+10Hz 0.0335338 -0.0455546
+ 6.6e+10Hz 0.0335584 -0.0456712
+ 6.61e+10Hz 0.0335828 -0.0457878
+ 6.62e+10Hz 0.0336071 -0.0459046
+ 6.63e+10Hz 0.0336313 -0.0460214
+ 6.64e+10Hz 0.0336554 -0.0461383
+ 6.65e+10Hz 0.0336794 -0.0462554
+ 6.66e+10Hz 0.0337032 -0.0463725
+ 6.67e+10Hz 0.0337269 -0.0464897
+ 6.68e+10Hz 0.0337505 -0.046607
+ 6.69e+10Hz 0.0337739 -0.0467244
+ 6.7e+10Hz 0.0337972 -0.0468419
+ 6.71e+10Hz 0.0338204 -0.0469595
+ 6.72e+10Hz 0.0338435 -0.0470771
+ 6.73e+10Hz 0.0338664 -0.0471949
+ 6.74e+10Hz 0.0338893 -0.0473128
+ 6.75e+10Hz 0.0339119 -0.0474307
+ 6.76e+10Hz 0.0339345 -0.0475487
+ 6.77e+10Hz 0.0339569 -0.0476668
+ 6.78e+10Hz 0.0339792 -0.047785
+ 6.79e+10Hz 0.0340014 -0.0479033
+ 6.8e+10Hz 0.0340234 -0.0480217
+ 6.81e+10Hz 0.0340454 -0.0481401
+ 6.82e+10Hz 0.0340672 -0.0482587
+ 6.83e+10Hz 0.0340888 -0.0483773
+ 6.84e+10Hz 0.0341104 -0.0484961
+ 6.85e+10Hz 0.0341318 -0.0486149
+ 6.86e+10Hz 0.0341531 -0.0487338
+ 6.87e+10Hz 0.0341743 -0.0488527
+ 6.88e+10Hz 0.0341953 -0.0489718
+ 6.89e+10Hz 0.0342162 -0.049091
+ 6.9e+10Hz 0.034237 -0.0492102
+ 6.91e+10Hz 0.0342576 -0.0493295
+ 6.92e+10Hz 0.0342781 -0.0494489
+ 6.93e+10Hz 0.0342985 -0.0495684
+ 6.94e+10Hz 0.0343188 -0.049688
+ 6.95e+10Hz 0.0343389 -0.0498076
+ 6.96e+10Hz 0.0343589 -0.0499274
+ 6.97e+10Hz 0.0343788 -0.0500472
+ 6.98e+10Hz 0.0343986 -0.0501671
+ 6.99e+10Hz 0.0344182 -0.050287
+ 7e+10Hz 0.0344377 -0.0504071
+ 7.01e+10Hz 0.0344571 -0.0505273
+ 7.02e+10Hz 0.0344763 -0.0506475
+ 7.03e+10Hz 0.0344954 -0.0507678
+ 7.04e+10Hz 0.0345144 -0.0508882
+ 7.05e+10Hz 0.0345333 -0.0510087
+ 7.06e+10Hz 0.034552 -0.0511292
+ 7.07e+10Hz 0.0345706 -0.0512499
+ 7.08e+10Hz 0.0345891 -0.0513706
+ 7.09e+10Hz 0.0346074 -0.0514914
+ 7.1e+10Hz 0.0346256 -0.0516123
+ 7.11e+10Hz 0.0346437 -0.0517332
+ 7.12e+10Hz 0.0346616 -0.0518543
+ 7.13e+10Hz 0.0346795 -0.0519754
+ 7.14e+10Hz 0.0346971 -0.0520966
+ 7.15e+10Hz 0.0347147 -0.0522179
+ 7.16e+10Hz 0.0347321 -0.0523392
+ 7.17e+10Hz 0.0347494 -0.0524607
+ 7.18e+10Hz 0.0347666 -0.0525822
+ 7.19e+10Hz 0.0347836 -0.0527038
+ 7.2e+10Hz 0.0348005 -0.0528255
+ 7.21e+10Hz 0.0348173 -0.0529472
+ 7.22e+10Hz 0.0348339 -0.0530691
+ 7.23e+10Hz 0.0348504 -0.053191
+ 7.24e+10Hz 0.0348668 -0.053313
+ 7.25e+10Hz 0.0348831 -0.053435
+ 7.26e+10Hz 0.0348992 -0.0535572
+ 7.27e+10Hz 0.0349151 -0.0536794
+ 7.28e+10Hz 0.034931 -0.0538017
+ 7.29e+10Hz 0.0349467 -0.0539241
+ 7.3e+10Hz 0.0349623 -0.0540466
+ 7.31e+10Hz 0.0349777 -0.0541691
+ 7.32e+10Hz 0.034993 -0.0542917
+ 7.33e+10Hz 0.0350082 -0.0544144
+ 7.34e+10Hz 0.0350232 -0.0545372
+ 7.35e+10Hz 0.0350381 -0.0546601
+ 7.36e+10Hz 0.0350529 -0.054783
+ 7.37e+10Hz 0.0350675 -0.054906
+ 7.38e+10Hz 0.035082 -0.0550291
+ 7.39e+10Hz 0.0350964 -0.0551522
+ 7.4e+10Hz 0.0351106 -0.0552755
+ 7.41e+10Hz 0.0351247 -0.0553988
+ 7.42e+10Hz 0.0351386 -0.0555222
+ 7.43e+10Hz 0.0351524 -0.0556456
+ 7.44e+10Hz 0.0351661 -0.0557692
+ 7.45e+10Hz 0.0351796 -0.0558928
+ 7.46e+10Hz 0.035193 -0.0560165
+ 7.47e+10Hz 0.0352062 -0.0561403
+ 7.48e+10Hz 0.0352194 -0.0562641
+ 7.49e+10Hz 0.0352323 -0.056388
+ 7.5e+10Hz 0.0352451 -0.056512
+ 7.51e+10Hz 0.0352578 -0.0566361
+ 7.52e+10Hz 0.0352704 -0.0567602
+ 7.53e+10Hz 0.0352828 -0.0568844
+ 7.54e+10Hz 0.035295 -0.0570087
+ 7.55e+10Hz 0.0353071 -0.0571331
+ 7.56e+10Hz 0.0353191 -0.0572575
+ 7.57e+10Hz 0.0353309 -0.057382
+ 7.58e+10Hz 0.0353426 -0.0575066
+ 7.59e+10Hz 0.0353542 -0.0576313
+ 7.6e+10Hz 0.0353656 -0.057756
+ 7.61e+10Hz 0.0353768 -0.0578808
+ 7.62e+10Hz 0.0353879 -0.0580057
+ 7.63e+10Hz 0.0353989 -0.0581307
+ 7.64e+10Hz 0.0354097 -0.0582557
+ 7.65e+10Hz 0.0354203 -0.0583808
+ 7.66e+10Hz 0.0354308 -0.058506
+ 7.67e+10Hz 0.0354412 -0.0586312
+ 7.68e+10Hz 0.0354514 -0.0587565
+ 7.69e+10Hz 0.0354615 -0.0588819
+ 7.7e+10Hz 0.0354714 -0.0590073
+ 7.71e+10Hz 0.0354812 -0.0591328
+ 7.72e+10Hz 0.0354908 -0.0592584
+ 7.73e+10Hz 0.0355002 -0.0593841
+ 7.74e+10Hz 0.0355095 -0.0595098
+ 7.75e+10Hz 0.0355187 -0.0596356
+ 7.76e+10Hz 0.0355277 -0.0597615
+ 7.77e+10Hz 0.0355365 -0.0598874
+ 7.78e+10Hz 0.0355452 -0.0600134
+ 7.79e+10Hz 0.0355538 -0.0601394
+ 7.8e+10Hz 0.0355622 -0.0602656
+ 7.81e+10Hz 0.0355704 -0.0603918
+ 7.82e+10Hz 0.0355784 -0.060518
+ 7.83e+10Hz 0.0355864 -0.0606443
+ 7.84e+10Hz 0.0355941 -0.0607707
+ 7.85e+10Hz 0.0356017 -0.0608972
+ 7.86e+10Hz 0.0356092 -0.0610237
+ 7.87e+10Hz 0.0356165 -0.0611503
+ 7.88e+10Hz 0.0356236 -0.0612769
+ 7.89e+10Hz 0.0356305 -0.0614036
+ 7.9e+10Hz 0.0356373 -0.0615304
+ 7.91e+10Hz 0.035644 -0.0616573
+ 7.92e+10Hz 0.0356505 -0.0617842
+ 7.93e+10Hz 0.0356568 -0.0619111
+ 7.94e+10Hz 0.0356629 -0.0620381
+ 7.95e+10Hz 0.0356689 -0.0621652
+ 7.96e+10Hz 0.0356748 -0.0622923
+ 7.97e+10Hz 0.0356805 -0.0624195
+ 7.98e+10Hz 0.035686 -0.0625468
+ 7.99e+10Hz 0.0356913 -0.0626741
+ 8e+10Hz 0.0356965 -0.0628015
+ 8.01e+10Hz 0.0357015 -0.0629289
+ 8.02e+10Hz 0.0357063 -0.0630564
+ 8.03e+10Hz 0.035711 -0.0631839
+ 8.04e+10Hz 0.0357155 -0.0633115
+ 8.05e+10Hz 0.0357198 -0.0634391
+ 8.06e+10Hz 0.035724 -0.0635668
+ 8.07e+10Hz 0.035728 -0.0636946
+ 8.08e+10Hz 0.0357319 -0.0638224
+ 8.09e+10Hz 0.0357355 -0.0639502
+ 8.1e+10Hz 0.035739 -0.0640781
+ 8.11e+10Hz 0.0357423 -0.0642061
+ 8.12e+10Hz 0.0357455 -0.0643341
+ 8.13e+10Hz 0.0357485 -0.0644622
+ 8.14e+10Hz 0.0357513 -0.0645903
+ 8.15e+10Hz 0.0357539 -0.0647184
+ 8.16e+10Hz 0.0357564 -0.0648466
+ 8.17e+10Hz 0.0357587 -0.0649749
+ 8.18e+10Hz 0.0357608 -0.0651031
+ 8.19e+10Hz 0.0357628 -0.0652315
+ 8.2e+10Hz 0.0357645 -0.0653599
+ 8.21e+10Hz 0.0357661 -0.0654883
+ 8.22e+10Hz 0.0357676 -0.0656167
+ 8.23e+10Hz 0.0357688 -0.0657453
+ 8.24e+10Hz 0.0357699 -0.0658738
+ 8.25e+10Hz 0.0357708 -0.0660024
+ 8.26e+10Hz 0.0357715 -0.066131
+ 8.27e+10Hz 0.035772 -0.0662597
+ 8.28e+10Hz 0.0357724 -0.0663884
+ 8.29e+10Hz 0.0357726 -0.0665171
+ 8.3e+10Hz 0.0357726 -0.0666459
+ 8.31e+10Hz 0.0357724 -0.0667747
+ 8.32e+10Hz 0.0357721 -0.0669036
+ 8.33e+10Hz 0.0357716 -0.0670325
+ 8.34e+10Hz 0.0357709 -0.0671614
+ 8.35e+10Hz 0.03577 -0.0672904
+ 8.36e+10Hz 0.0357689 -0.0674194
+ 8.37e+10Hz 0.0357677 -0.0675484
+ 8.38e+10Hz 0.0357663 -0.0676774
+ 8.39e+10Hz 0.0357647 -0.0678065
+ 8.4e+10Hz 0.0357629 -0.0679356
+ 8.41e+10Hz 0.0357609 -0.0680648
+ 8.42e+10Hz 0.0357588 -0.0681939
+ 8.43e+10Hz 0.0357565 -0.0683231
+ 8.44e+10Hz 0.035754 -0.0684523
+ 8.45e+10Hz 0.0357513 -0.0685816
+ 8.46e+10Hz 0.0357484 -0.0687108
+ 8.47e+10Hz 0.0357454 -0.0688401
+ 8.48e+10Hz 0.0357422 -0.0689695
+ 8.49e+10Hz 0.0357388 -0.0690988
+ 8.5e+10Hz 0.0357352 -0.0692281
+ 8.51e+10Hz 0.0357314 -0.0693575
+ 8.52e+10Hz 0.0357274 -0.0694869
+ 8.53e+10Hz 0.0357233 -0.0696163
+ 8.54e+10Hz 0.035719 -0.0697458
+ 8.55e+10Hz 0.0357145 -0.0698752
+ 8.56e+10Hz 0.0357098 -0.0700047
+ 8.57e+10Hz 0.0357049 -0.0701342
+ 8.58e+10Hz 0.0356999 -0.0702636
+ 8.59e+10Hz 0.0356946 -0.0703932
+ 8.6e+10Hz 0.0356892 -0.0705227
+ 8.61e+10Hz 0.0356836 -0.0706522
+ 8.62e+10Hz 0.0356778 -0.0707818
+ 8.63e+10Hz 0.0356719 -0.0709113
+ 8.64e+10Hz 0.0356657 -0.0710409
+ 8.65e+10Hz 0.0356594 -0.0711705
+ 8.66e+10Hz 0.0356529 -0.0713
+ 8.67e+10Hz 0.0356462 -0.0714296
+ 8.68e+10Hz 0.0356393 -0.0715592
+ 8.69e+10Hz 0.0356322 -0.0716888
+ 8.7e+10Hz 0.035625 -0.0718184
+ 8.71e+10Hz 0.0356176 -0.071948
+ 8.72e+10Hz 0.03561 -0.0720776
+ 8.73e+10Hz 0.0356022 -0.0722073
+ 8.74e+10Hz 0.0355942 -0.0723369
+ 8.75e+10Hz 0.035586 -0.0724665
+ 8.76e+10Hz 0.0355777 -0.0725961
+ 8.77e+10Hz 0.0355692 -0.0727257
+ 8.78e+10Hz 0.0355604 -0.0728553
+ 8.79e+10Hz 0.0355516 -0.072985
+ 8.8e+10Hz 0.0355425 -0.0731146
+ 8.81e+10Hz 0.0355332 -0.0732442
+ 8.82e+10Hz 0.0355238 -0.0733738
+ 8.83e+10Hz 0.0355142 -0.0735034
+ 8.84e+10Hz 0.0355044 -0.073633
+ 8.85e+10Hz 0.0354944 -0.0737625
+ 8.86e+10Hz 0.0354842 -0.0738921
+ 8.87e+10Hz 0.0354739 -0.0740217
+ 8.88e+10Hz 0.0354634 -0.0741512
+ 8.89e+10Hz 0.0354527 -0.0742808
+ 8.9e+10Hz 0.0354418 -0.0744103
+ 8.91e+10Hz 0.0354307 -0.0745398
+ 8.92e+10Hz 0.0354195 -0.0746693
+ 8.93e+10Hz 0.035408 -0.0747989
+ 8.94e+10Hz 0.0353964 -0.0749283
+ 8.95e+10Hz 0.0353846 -0.0750578
+ 8.96e+10Hz 0.0353727 -0.0751873
+ 8.97e+10Hz 0.0353605 -0.0753167
+ 8.98e+10Hz 0.0353482 -0.0754461
+ 8.99e+10Hz 0.0353357 -0.0755755
+ 9e+10Hz 0.035323 -0.0757049
+ 9.01e+10Hz 0.0353102 -0.0758343
+ 9.02e+10Hz 0.0352971 -0.0759637
+ 9.03e+10Hz 0.0352839 -0.076093
+ 9.04e+10Hz 0.0352705 -0.0762223
+ 9.05e+10Hz 0.035257 -0.0763516
+ 9.06e+10Hz 0.0352432 -0.0764809
+ 9.07e+10Hz 0.0352293 -0.0766101
+ 9.08e+10Hz 0.0352152 -0.0767394
+ 9.09e+10Hz 0.0352009 -0.0768686
+ 9.1e+10Hz 0.0351865 -0.0769978
+ 9.11e+10Hz 0.0351718 -0.0771269
+ 9.12e+10Hz 0.035157 -0.0772561
+ 9.13e+10Hz 0.0351421 -0.0773852
+ 9.14e+10Hz 0.0351269 -0.0775143
+ 9.15e+10Hz 0.0351116 -0.0776433
+ 9.16e+10Hz 0.0350961 -0.0777723
+ 9.17e+10Hz 0.0350804 -0.0779013
+ 9.18e+10Hz 0.0350645 -0.0780303
+ 9.19e+10Hz 0.0350485 -0.0781593
+ 9.2e+10Hz 0.0350323 -0.0782882
+ 9.21e+10Hz 0.035016 -0.0784171
+ 9.22e+10Hz 0.0349994 -0.0785459
+ 9.23e+10Hz 0.0349827 -0.0786748
+ 9.24e+10Hz 0.0349658 -0.0788035
+ 9.25e+10Hz 0.0349488 -0.0789323
+ 9.26e+10Hz 0.0349315 -0.079061
+ 9.27e+10Hz 0.0349141 -0.0791897
+ 9.28e+10Hz 0.0348966 -0.0793184
+ 9.29e+10Hz 0.0348788 -0.079447
+ 9.3e+10Hz 0.0348609 -0.0795756
+ 9.31e+10Hz 0.0348428 -0.0797042
+ 9.32e+10Hz 0.0348246 -0.0798327
+ 9.33e+10Hz 0.0348061 -0.0799612
+ 9.34e+10Hz 0.0347876 -0.0800897
+ 9.35e+10Hz 0.0347688 -0.0802181
+ 9.36e+10Hz 0.0347499 -0.0803465
+ 9.37e+10Hz 0.0347308 -0.0804749
+ 9.38e+10Hz 0.0347115 -0.0806032
+ 9.39e+10Hz 0.0346921 -0.0807314
+ 9.4e+10Hz 0.0346725 -0.0808597
+ 9.41e+10Hz 0.0346527 -0.0809879
+ 9.42e+10Hz 0.0346327 -0.081116
+ 9.43e+10Hz 0.0346126 -0.0812442
+ 9.44e+10Hz 0.0345924 -0.0813722
+ 9.45e+10Hz 0.0345719 -0.0815003
+ 9.46e+10Hz 0.0345513 -0.0816283
+ 9.47e+10Hz 0.0345306 -0.0817562
+ 9.48e+10Hz 0.0345096 -0.0818842
+ 9.49e+10Hz 0.0344885 -0.082012
+ 9.5e+10Hz 0.0344672 -0.0821399
+ 9.51e+10Hz 0.0344458 -0.0822677
+ 9.52e+10Hz 0.0344242 -0.0823954
+ 9.53e+10Hz 0.0344025 -0.0825231
+ 9.54e+10Hz 0.0343805 -0.0826508
+ 9.55e+10Hz 0.0343584 -0.0827784
+ 9.56e+10Hz 0.0343362 -0.082906
+ 9.57e+10Hz 0.0343137 -0.0830335
+ 9.58e+10Hz 0.0342912 -0.083161
+ 9.59e+10Hz 0.0342684 -0.0832884
+ 9.6e+10Hz 0.0342455 -0.0834158
+ 9.61e+10Hz 0.0342224 -0.0835432
+ 9.62e+10Hz 0.0341992 -0.0836705
+ 9.63e+10Hz 0.0341758 -0.0837978
+ 9.64e+10Hz 0.0341522 -0.083925
+ 9.65e+10Hz 0.0341285 -0.0840522
+ 9.66e+10Hz 0.0341046 -0.0841793
+ 9.67e+10Hz 0.0340805 -0.0843064
+ 9.68e+10Hz 0.0340563 -0.0844334
+ 9.69e+10Hz 0.0340319 -0.0845604
+ 9.7e+10Hz 0.0340074 -0.0846873
+ 9.71e+10Hz 0.0339827 -0.0848142
+ 9.72e+10Hz 0.0339578 -0.084941
+ 9.73e+10Hz 0.0339328 -0.0850678
+ 9.74e+10Hz 0.0339076 -0.0851945
+ 9.75e+10Hz 0.0338823 -0.0853212
+ 9.76e+10Hz 0.0338568 -0.0854479
+ 9.77e+10Hz 0.0338311 -0.0855744
+ 9.78e+10Hz 0.0338053 -0.085701
+ 9.79e+10Hz 0.0337792 -0.0858275
+ 9.8e+10Hz 0.0337531 -0.0859539
+ 9.81e+10Hz 0.0337268 -0.0860803
+ 9.82e+10Hz 0.0337003 -0.0862066
+ 9.83e+10Hz 0.0336736 -0.0863329
+ 9.84e+10Hz 0.0336468 -0.0864591
+ 9.85e+10Hz 0.0336199 -0.0865853
+ 9.86e+10Hz 0.0335928 -0.0867114
+ 9.87e+10Hz 0.0335655 -0.0868375
+ 9.88e+10Hz 0.033538 -0.0869635
+ 9.89e+10Hz 0.0335104 -0.0870894
+ 9.9e+10Hz 0.0334826 -0.0872153
+ 9.91e+10Hz 0.0334547 -0.0873412
+ 9.92e+10Hz 0.0334266 -0.087467
+ 9.93e+10Hz 0.0333984 -0.0875927
+ 9.94e+10Hz 0.03337 -0.0877184
+ 9.95e+10Hz 0.0333414 -0.0878441
+ 9.96e+10Hz 0.0333126 -0.0879696
+ 9.97e+10Hz 0.0332837 -0.0880951
+ 9.98e+10Hz 0.0332547 -0.0882206
+ 9.99e+10Hz 0.0332254 -0.088346
+ 1e+11Hz 0.0331961 -0.0884713
+ 1.001e+11Hz 0.0331665 -0.0885966
+ 1.002e+11Hz 0.0331368 -0.0887218
+ 1.003e+11Hz 0.033107 -0.088847
+ 1.004e+11Hz 0.0330769 -0.0889721
+ 1.005e+11Hz 0.0330467 -0.0890972
+ 1.006e+11Hz 0.0330164 -0.0892221
+ 1.007e+11Hz 0.0329859 -0.0893471
+ 1.008e+11Hz 0.0329552 -0.0894719
+ 1.009e+11Hz 0.0329243 -0.0895967
+ 1.01e+11Hz 0.0328933 -0.0897215
+ 1.011e+11Hz 0.0328622 -0.0898461
+ 1.012e+11Hz 0.0328309 -0.0899708
+ 1.013e+11Hz 0.0327994 -0.0900953
+ 1.014e+11Hz 0.0327677 -0.0902198
+ 1.015e+11Hz 0.0327359 -0.0903442
+ 1.016e+11Hz 0.0327039 -0.0904686
+ 1.017e+11Hz 0.0326718 -0.0905929
+ 1.018e+11Hz 0.0326395 -0.0907171
+ 1.019e+11Hz 0.032607 -0.0908413
+ 1.02e+11Hz 0.0325744 -0.0909654
+ 1.021e+11Hz 0.0325416 -0.0910894
+ 1.022e+11Hz 0.0325087 -0.0912133
+ 1.023e+11Hz 0.0324756 -0.0913372
+ 1.024e+11Hz 0.0324423 -0.0914611
+ 1.025e+11Hz 0.0324089 -0.0915848
+ 1.026e+11Hz 0.0323753 -0.0917085
+ 1.027e+11Hz 0.0323415 -0.0918321
+ 1.028e+11Hz 0.0323075 -0.0919557
+ 1.029e+11Hz 0.0322735 -0.0920791
+ 1.03e+11Hz 0.0322392 -0.0922025
+ 1.031e+11Hz 0.0322048 -0.0923259
+ 1.032e+11Hz 0.0321702 -0.0924491
+ 1.033e+11Hz 0.0321354 -0.0925723
+ 1.034e+11Hz 0.0321005 -0.0926954
+ 1.035e+11Hz 0.0320655 -0.0928184
+ 1.036e+11Hz 0.0320302 -0.0929414
+ 1.037e+11Hz 0.0319948 -0.0930642
+ 1.038e+11Hz 0.0319592 -0.093187
+ 1.039e+11Hz 0.0319235 -0.0933097
+ 1.04e+11Hz 0.0318876 -0.0934324
+ 1.041e+11Hz 0.0318515 -0.093555
+ 1.042e+11Hz 0.0318153 -0.0936774
+ 1.043e+11Hz 0.0317789 -0.0937998
+ 1.044e+11Hz 0.0317424 -0.0939222
+ 1.045e+11Hz 0.0317057 -0.0940444
+ 1.046e+11Hz 0.0316688 -0.0941666
+ 1.047e+11Hz 0.0316317 -0.0942886
+ 1.048e+11Hz 0.0315945 -0.0944106
+ 1.049e+11Hz 0.0315571 -0.0945325
+ 1.05e+11Hz 0.0315196 -0.0946543
+ 1.051e+11Hz 0.0314819 -0.0947761
+ 1.052e+11Hz 0.031444 -0.0948977
+ 1.053e+11Hz 0.031406 -0.0950193
+ 1.054e+11Hz 0.0313678 -0.0951407
+ 1.055e+11Hz 0.0313294 -0.0952621
+ 1.056e+11Hz 0.0312909 -0.0953834
+ 1.057e+11Hz 0.0312522 -0.0955046
+ 1.058e+11Hz 0.0312133 -0.0956257
+ 1.059e+11Hz 0.0311743 -0.0957467
+ 1.06e+11Hz 0.0311351 -0.0958676
+ 1.061e+11Hz 0.0310957 -0.0959885
+ 1.062e+11Hz 0.0310562 -0.0961092
+ 1.063e+11Hz 0.0310165 -0.0962299
+ 1.064e+11Hz 0.0309767 -0.0963504
+ 1.065e+11Hz 0.0309367 -0.0964708
+ 1.066e+11Hz 0.0308965 -0.0965912
+ 1.067e+11Hz 0.0308562 -0.0967114
+ 1.068e+11Hz 0.0308157 -0.0968316
+ 1.069e+11Hz 0.030775 -0.0969516
+ 1.07e+11Hz 0.0307342 -0.0970716
+ 1.071e+11Hz 0.0306932 -0.0971914
+ 1.072e+11Hz 0.030652 -0.0973111
+ 1.073e+11Hz 0.0306107 -0.0974308
+ 1.074e+11Hz 0.0305692 -0.0975503
+ 1.075e+11Hz 0.0305276 -0.0976697
+ 1.076e+11Hz 0.0304858 -0.097789
+ 1.077e+11Hz 0.0304438 -0.0979082
+ 1.078e+11Hz 0.0304017 -0.0980273
+ 1.079e+11Hz 0.0303594 -0.0981463
+ 1.08e+11Hz 0.030317 -0.0982652
+ 1.081e+11Hz 0.0302743 -0.098384
+ 1.082e+11Hz 0.0302316 -0.0985026
+ 1.083e+11Hz 0.0301887 -0.0986212
+ 1.084e+11Hz 0.0301456 -0.0987396
+ 1.085e+11Hz 0.0301023 -0.0988579
+ 1.086e+11Hz 0.0300589 -0.0989761
+ 1.087e+11Hz 0.0300153 -0.0990942
+ 1.088e+11Hz 0.0299716 -0.0992122
+ 1.089e+11Hz 0.0299277 -0.09933
+ 1.09e+11Hz 0.0298837 -0.0994478
+ 1.091e+11Hz 0.0298395 -0.0995654
+ 1.092e+11Hz 0.0297951 -0.0996829
+ 1.093e+11Hz 0.0297506 -0.0998002
+ 1.094e+11Hz 0.0297059 -0.0999175
+ 1.095e+11Hz 0.0296611 -0.100035
+ 1.096e+11Hz 0.0296161 -0.100152
+ 1.097e+11Hz 0.0295709 -0.100268
+ 1.098e+11Hz 0.0295256 -0.100385
+ 1.099e+11Hz 0.0294802 -0.100502
+ 1.1e+11Hz 0.0294346 -0.100618
+ 1.101e+11Hz 0.0293888 -0.100735
+ 1.102e+11Hz 0.0293429 -0.100851
+ 1.103e+11Hz 0.0292968 -0.100967
+ 1.104e+11Hz 0.0292506 -0.101083
+ 1.105e+11Hz 0.0292042 -0.101199
+ 1.106e+11Hz 0.0291577 -0.101315
+ 1.107e+11Hz 0.029111 -0.10143
+ 1.108e+11Hz 0.0290642 -0.101545
+ 1.109e+11Hz 0.0290172 -0.101661
+ 1.11e+11Hz 0.0289701 -0.101776
+ 1.111e+11Hz 0.0289228 -0.101891
+ 1.112e+11Hz 0.0288754 -0.102006
+ 1.113e+11Hz 0.0288279 -0.102121
+ 1.114e+11Hz 0.0287802 -0.102235
+ 1.115e+11Hz 0.0287323 -0.10235
+ 1.116e+11Hz 0.0286843 -0.102464
+ 1.117e+11Hz 0.0286361 -0.102578
+ 1.118e+11Hz 0.0285879 -0.102692
+ 1.119e+11Hz 0.0285394 -0.102806
+ 1.12e+11Hz 0.0284908 -0.10292
+ 1.121e+11Hz 0.0284421 -0.103034
+ 1.122e+11Hz 0.0283933 -0.103147
+ 1.123e+11Hz 0.0283443 -0.10326
+ 1.124e+11Hz 0.0282951 -0.103373
+ 1.125e+11Hz 0.0282458 -0.103486
+ 1.126e+11Hz 0.0281964 -0.103599
+ 1.127e+11Hz 0.0281469 -0.103712
+ 1.128e+11Hz 0.0280972 -0.103825
+ 1.129e+11Hz 0.0280473 -0.103937
+ 1.13e+11Hz 0.0279974 -0.104049
+ 1.131e+11Hz 0.0279473 -0.104161
+ 1.132e+11Hz 0.027897 -0.104273
+ 1.133e+11Hz 0.0278467 -0.104385
+ 1.134e+11Hz 0.0277962 -0.104497
+ 1.135e+11Hz 0.0277456 -0.104608
+ 1.136e+11Hz 0.0276948 -0.10472
+ 1.137e+11Hz 0.0276439 -0.104831
+ 1.138e+11Hz 0.0275929 -0.104942
+ 1.139e+11Hz 0.0275417 -0.105053
+ 1.14e+11Hz 0.0274904 -0.105163
+ 1.141e+11Hz 0.027439 -0.105274
+ 1.142e+11Hz 0.0273875 -0.105384
+ 1.143e+11Hz 0.0273358 -0.105495
+ 1.144e+11Hz 0.0272841 -0.105605
+ 1.145e+11Hz 0.0272322 -0.105715
+ 1.146e+11Hz 0.0271801 -0.105824
+ 1.147e+11Hz 0.027128 -0.105934
+ 1.148e+11Hz 0.0270757 -0.106043
+ 1.149e+11Hz 0.0270233 -0.106153
+ 1.15e+11Hz 0.0269708 -0.106262
+ 1.151e+11Hz 0.0269182 -0.106371
+ 1.152e+11Hz 0.0268654 -0.10648
+ 1.153e+11Hz 0.0268126 -0.106588
+ 1.154e+11Hz 0.0267596 -0.106697
+ 1.155e+11Hz 0.0267065 -0.106805
+ 1.156e+11Hz 0.0266533 -0.106913
+ 1.157e+11Hz 0.0266 -0.107021
+ 1.158e+11Hz 0.0265465 -0.107129
+ 1.159e+11Hz 0.026493 -0.107236
+ 1.16e+11Hz 0.0264393 -0.107344
+ 1.161e+11Hz 0.0263855 -0.107451
+ 1.162e+11Hz 0.0263317 -0.107558
+ 1.163e+11Hz 0.0262777 -0.107665
+ 1.164e+11Hz 0.0262236 -0.107772
+ 1.165e+11Hz 0.0261694 -0.107879
+ 1.166e+11Hz 0.0261151 -0.107985
+ 1.167e+11Hz 0.0260606 -0.108091
+ 1.168e+11Hz 0.0260061 -0.108197
+ 1.169e+11Hz 0.0259515 -0.108303
+ 1.17e+11Hz 0.0258968 -0.108409
+ 1.171e+11Hz 0.0258419 -0.108515
+ 1.172e+11Hz 0.025787 -0.10862
+ 1.173e+11Hz 0.025732 -0.108725
+ 1.174e+11Hz 0.0256769 -0.10883
+ 1.175e+11Hz 0.0256216 -0.108935
+ 1.176e+11Hz 0.0255663 -0.10904
+ 1.177e+11Hz 0.0255109 -0.109145
+ 1.178e+11Hz 0.0254553 -0.109249
+ 1.179e+11Hz 0.0253997 -0.109353
+ 1.18e+11Hz 0.025344 -0.109457
+ 1.181e+11Hz 0.0252882 -0.109561
+ 1.182e+11Hz 0.0252323 -0.109665
+ 1.183e+11Hz 0.0251763 -0.109769
+ 1.184e+11Hz 0.0251202 -0.109872
+ 1.185e+11Hz 0.025064 -0.109975
+ 1.186e+11Hz 0.0250078 -0.110078
+ 1.187e+11Hz 0.0249514 -0.110181
+ 1.188e+11Hz 0.024895 -0.110284
+ 1.189e+11Hz 0.0248384 -0.110386
+ 1.19e+11Hz 0.0247818 -0.110488
+ 1.191e+11Hz 0.0247251 -0.110591
+ 1.192e+11Hz 0.0246683 -0.110693
+ 1.193e+11Hz 0.0246114 -0.110794
+ 1.194e+11Hz 0.0245544 -0.110896
+ 1.195e+11Hz 0.0244974 -0.110997
+ 1.196e+11Hz 0.0244403 -0.111099
+ 1.197e+11Hz 0.024383 -0.1112
+ 1.198e+11Hz 0.0243257 -0.111301
+ 1.199e+11Hz 0.0242683 -0.111402
+ 1.2e+11Hz 0.0242109 -0.111502
+ 1.201e+11Hz 0.0241533 -0.111603
+ 1.202e+11Hz 0.0240957 -0.111703
+ 1.203e+11Hz 0.024038 -0.111803
+ 1.204e+11Hz 0.0239802 -0.111903
+ 1.205e+11Hz 0.0239223 -0.112003
+ 1.206e+11Hz 0.0238644 -0.112102
+ 1.207e+11Hz 0.0238064 -0.112202
+ 1.208e+11Hz 0.0237482 -0.112301
+ 1.209e+11Hz 0.0236901 -0.1124
+ 1.21e+11Hz 0.0236318 -0.112499
+ 1.211e+11Hz 0.0235735 -0.112598
+ 1.212e+11Hz 0.0235151 -0.112696
+ 1.213e+11Hz 0.0234566 -0.112795
+ 1.214e+11Hz 0.023398 -0.112893
+ 1.215e+11Hz 0.0233394 -0.112991
+ 1.216e+11Hz 0.0232807 -0.113089
+ 1.217e+11Hz 0.0232219 -0.113186
+ 1.218e+11Hz 0.0231631 -0.113284
+ 1.219e+11Hz 0.0231041 -0.113381
+ 1.22e+11Hz 0.0230451 -0.113478
+ 1.221e+11Hz 0.0229861 -0.113575
+ 1.222e+11Hz 0.0229269 -0.113672
+ 1.223e+11Hz 0.0228677 -0.113769
+ 1.224e+11Hz 0.0228084 -0.113865
+ 1.225e+11Hz 0.022749 -0.113962
+ 1.226e+11Hz 0.0226896 -0.114058
+ 1.227e+11Hz 0.0226301 -0.114154
+ 1.228e+11Hz 0.0225706 -0.11425
+ 1.229e+11Hz 0.0225109 -0.114345
+ 1.23e+11Hz 0.0224512 -0.114441
+ 1.231e+11Hz 0.0223914 -0.114536
+ 1.232e+11Hz 0.0223316 -0.114631
+ 1.233e+11Hz 0.0222717 -0.114726
+ 1.234e+11Hz 0.0222117 -0.114821
+ 1.235e+11Hz 0.0221516 -0.114915
+ 1.236e+11Hz 0.0220915 -0.11501
+ 1.237e+11Hz 0.0220313 -0.115104
+ 1.238e+11Hz 0.0219711 -0.115198
+ 1.239e+11Hz 0.0219108 -0.115292
+ 1.24e+11Hz 0.0218504 -0.115386
+ 1.241e+11Hz 0.0217899 -0.115479
+ 1.242e+11Hz 0.0217294 -0.115573
+ 1.243e+11Hz 0.0216688 -0.115666
+ 1.244e+11Hz 0.0216081 -0.115759
+ 1.245e+11Hz 0.0215474 -0.115852
+ 1.246e+11Hz 0.0214866 -0.115944
+ 1.247e+11Hz 0.0214257 -0.116037
+ 1.248e+11Hz 0.0213648 -0.116129
+ 1.249e+11Hz 0.0213038 -0.116222
+ 1.25e+11Hz 0.0212428 -0.116314
+ 1.251e+11Hz 0.0211816 -0.116405
+ 1.252e+11Hz 0.0211204 -0.116497
+ 1.253e+11Hz 0.0210592 -0.116588
+ 1.254e+11Hz 0.0209978 -0.11668
+ 1.255e+11Hz 0.0209364 -0.116771
+ 1.256e+11Hz 0.020875 -0.116862
+ 1.257e+11Hz 0.0208135 -0.116953
+ 1.258e+11Hz 0.0207519 -0.117043
+ 1.259e+11Hz 0.0206902 -0.117134
+ 1.26e+11Hz 0.0206285 -0.117224
+ 1.261e+11Hz 0.0205667 -0.117314
+ 1.262e+11Hz 0.0205048 -0.117404
+ 1.263e+11Hz 0.0204429 -0.117494
+ 1.264e+11Hz 0.0203809 -0.117583
+ 1.265e+11Hz 0.0203189 -0.117673
+ 1.266e+11Hz 0.0202567 -0.117762
+ 1.267e+11Hz 0.0201945 -0.117851
+ 1.268e+11Hz 0.0201323 -0.11794
+ 1.269e+11Hz 0.02007 -0.118028
+ 1.27e+11Hz 0.0200076 -0.118117
+ 1.271e+11Hz 0.0199451 -0.118205
+ 1.272e+11Hz 0.0198826 -0.118293
+ 1.273e+11Hz 0.01982 -0.118381
+ 1.274e+11Hz 0.0197574 -0.118469
+ 1.275e+11Hz 0.0196947 -0.118557
+ 1.276e+11Hz 0.0196319 -0.118644
+ 1.277e+11Hz 0.0195691 -0.118731
+ 1.278e+11Hz 0.0195062 -0.118818
+ 1.279e+11Hz 0.0194432 -0.118905
+ 1.28e+11Hz 0.0193801 -0.118992
+ 1.281e+11Hz 0.019317 -0.119078
+ 1.282e+11Hz 0.0192539 -0.119165
+ 1.283e+11Hz 0.0191906 -0.119251
+ 1.284e+11Hz 0.0191273 -0.119337
+ 1.285e+11Hz 0.019064 -0.119422
+ 1.286e+11Hz 0.0190005 -0.119508
+ 1.287e+11Hz 0.018937 -0.119593
+ 1.288e+11Hz 0.0188735 -0.119678
+ 1.289e+11Hz 0.0188099 -0.119763
+ 1.29e+11Hz 0.0187462 -0.119848
+ 1.291e+11Hz 0.0186824 -0.119933
+ 1.292e+11Hz 0.0186186 -0.120017
+ 1.293e+11Hz 0.0185547 -0.120101
+ 1.294e+11Hz 0.0184908 -0.120186
+ 1.295e+11Hz 0.0184268 -0.120269
+ 1.296e+11Hz 0.0183627 -0.120353
+ 1.297e+11Hz 0.0182986 -0.120436
+ 1.298e+11Hz 0.0182344 -0.12052
+ 1.299e+11Hz 0.0181701 -0.120603
+ 1.3e+11Hz 0.0181058 -0.120686
+ 1.301e+11Hz 0.0180415 -0.120768
+ 1.302e+11Hz 0.017977 -0.120851
+ 1.303e+11Hz 0.0179125 -0.120933
+ 1.304e+11Hz 0.017848 -0.121015
+ 1.305e+11Hz 0.0177833 -0.121097
+ 1.306e+11Hz 0.0177186 -0.121178
+ 1.307e+11Hz 0.0176539 -0.12126
+ 1.308e+11Hz 0.0175891 -0.121341
+ 1.309e+11Hz 0.0175243 -0.121422
+ 1.31e+11Hz 0.0174593 -0.121503
+ 1.311e+11Hz 0.0173944 -0.121583
+ 1.312e+11Hz 0.0173293 -0.121664
+ 1.313e+11Hz 0.0172642 -0.121744
+ 1.314e+11Hz 0.0171991 -0.121824
+ 1.315e+11Hz 0.0171339 -0.121904
+ 1.316e+11Hz 0.0170687 -0.121983
+ 1.317e+11Hz 0.0170033 -0.122063
+ 1.318e+11Hz 0.016938 -0.122142
+ 1.319e+11Hz 0.0168726 -0.122221
+ 1.32e+11Hz 0.0168071 -0.122299
+ 1.321e+11Hz 0.0167416 -0.122378
+ 1.322e+11Hz 0.016676 -0.122456
+ 1.323e+11Hz 0.0166104 -0.122534
+ 1.324e+11Hz 0.0165447 -0.122612
+ 1.325e+11Hz 0.016479 -0.122689
+ 1.326e+11Hz 0.0164132 -0.122767
+ 1.327e+11Hz 0.0163474 -0.122844
+ 1.328e+11Hz 0.0162815 -0.122921
+ 1.329e+11Hz 0.0162156 -0.122997
+ 1.33e+11Hz 0.0161497 -0.123074
+ 1.331e+11Hz 0.0160837 -0.12315
+ 1.332e+11Hz 0.0160176 -0.123226
+ 1.333e+11Hz 0.0159515 -0.123302
+ 1.334e+11Hz 0.0158854 -0.123378
+ 1.335e+11Hz 0.0158193 -0.123453
+ 1.336e+11Hz 0.0157531 -0.123528
+ 1.337e+11Hz 0.0156868 -0.123603
+ 1.338e+11Hz 0.0156205 -0.123677
+ 1.339e+11Hz 0.0155542 -0.123752
+ 1.34e+11Hz 0.0154879 -0.123826
+ 1.341e+11Hz 0.0154215 -0.1239
+ 1.342e+11Hz 0.0153551 -0.123974
+ 1.343e+11Hz 0.0152886 -0.124047
+ 1.344e+11Hz 0.0152221 -0.12412
+ 1.345e+11Hz 0.0151556 -0.124193
+ 1.346e+11Hz 0.0150891 -0.124266
+ 1.347e+11Hz 0.0150225 -0.124338
+ 1.348e+11Hz 0.0149559 -0.124411
+ 1.349e+11Hz 0.0148893 -0.124483
+ 1.35e+11Hz 0.0148226 -0.124554
+ 1.351e+11Hz 0.014756 -0.124626
+ 1.352e+11Hz 0.0146893 -0.124697
+ 1.353e+11Hz 0.0146226 -0.124768
+ 1.354e+11Hz 0.0145558 -0.124839
+ 1.355e+11Hz 0.0144891 -0.12491
+ 1.356e+11Hz 0.0144223 -0.12498
+ 1.357e+11Hz 0.0143556 -0.12505
+ 1.358e+11Hz 0.0142888 -0.12512
+ 1.359e+11Hz 0.014222 -0.125189
+ 1.36e+11Hz 0.0141552 -0.125258
+ 1.361e+11Hz 0.0140884 -0.125328
+ 1.362e+11Hz 0.0140216 -0.125396
+ 1.363e+11Hz 0.0139547 -0.125465
+ 1.364e+11Hz 0.0138879 -0.125533
+ 1.365e+11Hz 0.0138211 -0.125601
+ 1.366e+11Hz 0.0137542 -0.125669
+ 1.367e+11Hz 0.0136874 -0.125737
+ 1.368e+11Hz 0.0136206 -0.125804
+ 1.369e+11Hz 0.0135537 -0.125871
+ 1.37e+11Hz 0.0134869 -0.125938
+ 1.371e+11Hz 0.0134201 -0.126004
+ 1.372e+11Hz 0.0133533 -0.12607
+ 1.373e+11Hz 0.0132865 -0.126136
+ 1.374e+11Hz 0.0132197 -0.126202
+ 1.375e+11Hz 0.0131529 -0.126268
+ 1.376e+11Hz 0.0130862 -0.126333
+ 1.377e+11Hz 0.0130194 -0.126398
+ 1.378e+11Hz 0.0129527 -0.126463
+ 1.379e+11Hz 0.012886 -0.126527
+ 1.38e+11Hz 0.0128193 -0.126591
+ 1.381e+11Hz 0.0127527 -0.126655
+ 1.382e+11Hz 0.0126861 -0.126719
+ 1.383e+11Hz 0.0126195 -0.126782
+ 1.384e+11Hz 0.0125529 -0.126846
+ 1.385e+11Hz 0.0124863 -0.126909
+ 1.386e+11Hz 0.0124198 -0.126971
+ 1.387e+11Hz 0.0123533 -0.127034
+ 1.388e+11Hz 0.0122869 -0.127096
+ 1.389e+11Hz 0.0122205 -0.127158
+ 1.39e+11Hz 0.0121541 -0.12722
+ 1.391e+11Hz 0.0120878 -0.127281
+ 1.392e+11Hz 0.0120215 -0.127342
+ 1.393e+11Hz 0.0119553 -0.127403
+ 1.394e+11Hz 0.011889 -0.127464
+ 1.395e+11Hz 0.0118229 -0.127524
+ 1.396e+11Hz 0.0117568 -0.127584
+ 1.397e+11Hz 0.0116907 -0.127644
+ 1.398e+11Hz 0.0116247 -0.127704
+ 1.399e+11Hz 0.0115588 -0.127763
+ 1.4e+11Hz 0.0114929 -0.127822
+ 1.401e+11Hz 0.0114271 -0.127881
+ 1.402e+11Hz 0.0113613 -0.12794
+ 1.403e+11Hz 0.0112956 -0.127998
+ 1.404e+11Hz 0.0112299 -0.128056
+ 1.405e+11Hz 0.0111643 -0.128114
+ 1.406e+11Hz 0.0110988 -0.128172
+ 1.407e+11Hz 0.0110333 -0.128229
+ 1.408e+11Hz 0.0109679 -0.128286
+ 1.409e+11Hz 0.0109026 -0.128343
+ 1.41e+11Hz 0.0108373 -0.1284
+ 1.411e+11Hz 0.0107721 -0.128456
+ 1.412e+11Hz 0.010707 -0.128513
+ 1.413e+11Hz 0.010642 -0.128569
+ 1.414e+11Hz 0.010577 -0.128624
+ 1.415e+11Hz 0.0105122 -0.12868
+ 1.416e+11Hz 0.0104474 -0.128735
+ 1.417e+11Hz 0.0103826 -0.12879
+ 1.418e+11Hz 0.010318 -0.128845
+ 1.419e+11Hz 0.0102534 -0.128899
+ 1.42e+11Hz 0.010189 -0.128953
+ 1.421e+11Hz 0.0101246 -0.129007
+ 1.422e+11Hz 0.0100603 -0.129061
+ 1.423e+11Hz 0.00999607 -0.129115
+ 1.424e+11Hz 0.00993194 -0.129168
+ 1.425e+11Hz 0.00986791 -0.129221
+ 1.426e+11Hz 0.00980397 -0.129274
+ 1.427e+11Hz 0.00974012 -0.129327
+ 1.428e+11Hz 0.00967636 -0.129379
+ 1.429e+11Hz 0.0096127 -0.129432
+ 1.43e+11Hz 0.00954914 -0.129484
+ 1.431e+11Hz 0.00948567 -0.129535
+ 1.432e+11Hz 0.0094223 -0.129587
+ 1.433e+11Hz 0.00935902 -0.129638
+ 1.434e+11Hz 0.00929585 -0.129689
+ 1.435e+11Hz 0.00923278 -0.12974
+ 1.436e+11Hz 0.00916981 -0.129791
+ 1.437e+11Hz 0.00910694 -0.129841
+ 1.438e+11Hz 0.00904417 -0.129892
+ 1.439e+11Hz 0.0089815 -0.129942
+ 1.44e+11Hz 0.00891894 -0.129992
+ 1.441e+11Hz 0.00885649 -0.130041
+ 1.442e+11Hz 0.00879414 -0.130091
+ 1.443e+11Hz 0.00873189 -0.13014
+ 1.444e+11Hz 0.00866975 -0.130189
+ 1.445e+11Hz 0.00860772 -0.130238
+ 1.446e+11Hz 0.0085458 -0.130286
+ 1.447e+11Hz 0.00848398 -0.130335
+ 1.448e+11Hz 0.00842227 -0.130383
+ 1.449e+11Hz 0.00836067 -0.130431
+ 1.45e+11Hz 0.00829918 -0.130479
+ 1.451e+11Hz 0.0082378 -0.130526
+ 1.452e+11Hz 0.00817652 -0.130574
+ 1.453e+11Hz 0.00811536 -0.130621
+ 1.454e+11Hz 0.00805431 -0.130668
+ 1.455e+11Hz 0.00799336 -0.130715
+ 1.456e+11Hz 0.00793253 -0.130762
+ 1.457e+11Hz 0.00787181 -0.130808
+ 1.458e+11Hz 0.00781119 -0.130854
+ 1.459e+11Hz 0.00775069 -0.130901
+ 1.46e+11Hz 0.0076903 -0.130946
+ 1.461e+11Hz 0.00763001 -0.130992
+ 1.462e+11Hz 0.00756984 -0.131038
+ 1.463e+11Hz 0.00750978 -0.131083
+ 1.464e+11Hz 0.00744982 -0.131128
+ 1.465e+11Hz 0.00738998 -0.131173
+ 1.466e+11Hz 0.00733024 -0.131218
+ 1.467e+11Hz 0.00727062 -0.131263
+ 1.468e+11Hz 0.0072111 -0.131307
+ 1.469e+11Hz 0.00715169 -0.131352
+ 1.47e+11Hz 0.00709239 -0.131396
+ 1.471e+11Hz 0.0070332 -0.13144
+ 1.472e+11Hz 0.00697411 -0.131484
+ 1.473e+11Hz 0.00691513 -0.131528
+ 1.474e+11Hz 0.00685626 -0.131571
+ 1.475e+11Hz 0.00679749 -0.131614
+ 1.476e+11Hz 0.00673883 -0.131658
+ 1.477e+11Hz 0.00668027 -0.131701
+ 1.478e+11Hz 0.00662182 -0.131744
+ 1.479e+11Hz 0.00656347 -0.131786
+ 1.48e+11Hz 0.00650522 -0.131829
+ 1.481e+11Hz 0.00644708 -0.131871
+ 1.482e+11Hz 0.00638904 -0.131913
+ 1.483e+11Hz 0.00633109 -0.131955
+ 1.484e+11Hz 0.00627325 -0.131997
+ 1.485e+11Hz 0.00621551 -0.132039
+ 1.486e+11Hz 0.00615786 -0.132081
+ 1.487e+11Hz 0.00610032 -0.132122
+ 1.488e+11Hz 0.00604287 -0.132163
+ 1.489e+11Hz 0.00598551 -0.132204
+ 1.49e+11Hz 0.00592826 -0.132245
+ 1.491e+11Hz 0.00587109 -0.132286
+ 1.492e+11Hz 0.00581402 -0.132327
+ 1.493e+11Hz 0.00575704 -0.132367
+ 1.494e+11Hz 0.00570016 -0.132408
+ 1.495e+11Hz 0.00564336 -0.132448
+ 1.496e+11Hz 0.00558666 -0.132488
+ 1.497e+11Hz 0.00553004 -0.132528
+ 1.498e+11Hz 0.00547352 -0.132568
+ 1.499e+11Hz 0.00541708 -0.132607
+ 1.5e+11Hz 0.00536073 -0.132647
+ ]

.ENDS
.SUBCKT Sub_SPfile_X4 1 2 3
R1N 1 10 -50
R1P 10 11 100
R2N 2 20 -50
R2P 20 21 100

A11 %vd(10 3) %vd(11, 12) xfer1
.model xfer1 xfer R_I=true table=[
+ 0Hz 0.00482376 0
+ 1e+08Hz 0.00482395 1.93737e-06
+ 2e+08Hz 0.00482452 3.86743e-06
+ 3e+08Hz 0.00482548 5.78289e-06
+ 4e+08Hz 0.00482681 7.67645e-06
+ 5e+08Hz 0.00482853 9.54082e-06
+ 6e+08Hz 0.00483063 1.13687e-05
+ 7e+08Hz 0.0048331 1.3153e-05
+ 8e+08Hz 0.00483596 1.48863e-05
+ 9e+08Hz 0.00483919 1.65614e-05
+ 1e+09Hz 0.0048428 1.81712e-05
+ 1.1e+09Hz 0.00484679 1.97086e-05
+ 1.2e+09Hz 0.00485114 2.11664e-05
+ 1.3e+09Hz 0.00485587 2.25375e-05
+ 1.4e+09Hz 0.00486097 2.3815e-05
+ 1.5e+09Hz 0.00486643 2.49917e-05
+ 1.6e+09Hz 0.00487226 2.60609e-05
+ 1.7e+09Hz 0.00487846 2.70156e-05
+ 1.8e+09Hz 0.00488501 2.78489e-05
+ 1.9e+09Hz 0.00489192 2.85541e-05
+ 2e+09Hz 0.00489919 2.91245e-05
+ 2.1e+09Hz 0.00490681 2.95534e-05
+ 2.2e+09Hz 0.00491478 2.98342e-05
+ 2.3e+09Hz 0.00492309 2.99605e-05
+ 2.4e+09Hz 0.00493175 2.99257e-05
+ 2.5e+09Hz 0.00494075 2.97235e-05
+ 2.6e+09Hz 0.00495008 2.93477e-05
+ 2.7e+09Hz 0.00495975 2.87919e-05
+ 2.8e+09Hz 0.00496975 2.80502e-05
+ 2.9e+09Hz 0.00498007 2.71164e-05
+ 3e+09Hz 0.00499071 2.59846e-05
+ 3.1e+09Hz 0.00500167 2.4649e-05
+ 3.2e+09Hz 0.00501294 2.31038e-05
+ 3.3e+09Hz 0.00502452 2.13433e-05
+ 3.4e+09Hz 0.0050364 1.93619e-05
+ 3.5e+09Hz 0.00504859 1.71543e-05
+ 3.6e+09Hz 0.00506107 1.4715e-05
+ 3.7e+09Hz 0.00507383 1.20388e-05
+ 3.8e+09Hz 0.00508689 9.12049e-06
+ 3.9e+09Hz 0.00510022 5.9551e-06
+ 4e+09Hz 0.00511383 2.53768e-06
+ 4.1e+09Hz 0.00512771 -1.13658e-06
+ 4.2e+09Hz 0.00514185 -5.07238e-06
+ 4.3e+09Hz 0.00515626 -9.2743e-06
+ 4.4e+09Hz 0.00517091 -1.37468e-05
+ 4.5e+09Hz 0.00518582 -1.84942e-05
+ 4.6e+09Hz 0.00520097 -2.35208e-05
+ 4.7e+09Hz 0.00521636 -2.88306e-05
+ 4.8e+09Hz 0.00523198 -3.44276e-05
+ 4.9e+09Hz 0.00524782 -4.03157e-05
+ 5e+09Hz 0.00526389 -4.64986e-05
+ 5.1e+09Hz 0.00528017 -5.29798e-05
+ 5.2e+09Hz 0.00529666 -5.97629e-05
+ 5.3e+09Hz 0.00531335 -6.68512e-05
+ 5.4e+09Hz 0.00533024 -7.42479e-05
+ 5.5e+09Hz 0.00534732 -8.1956e-05
+ 5.6e+09Hz 0.00536459 -8.99785e-05
+ 5.7e+09Hz 0.00538203 -9.83183e-05
+ 5.8e+09Hz 0.00539964 -0.000106978
+ 5.9e+09Hz 0.00541742 -0.00011596
+ 6e+09Hz 0.00543536 -0.000125267
+ 6.1e+09Hz 0.00545346 -0.000134901
+ 6.2e+09Hz 0.0054717 -0.000144864
+ 6.3e+09Hz 0.00549008 -0.000155159
+ 6.4e+09Hz 0.00550859 -0.000165787
+ 6.5e+09Hz 0.00552723 -0.00017675
+ 6.6e+09Hz 0.005546 -0.000188049
+ 6.7e+09Hz 0.00556488 -0.000199686
+ 6.8e+09Hz 0.00558387 -0.000211663
+ 6.9e+09Hz 0.00560296 -0.00022398
+ 7e+09Hz 0.00562214 -0.000236638
+ 7.1e+09Hz 0.00564142 -0.000249639
+ 7.2e+09Hz 0.00566077 -0.000262984
+ 7.3e+09Hz 0.00568021 -0.000276673
+ 7.4e+09Hz 0.00569971 -0.000290706
+ 7.5e+09Hz 0.00571928 -0.000305084
+ 7.6e+09Hz 0.00573891 -0.000319807
+ 7.7e+09Hz 0.00575858 -0.000334876
+ 7.8e+09Hz 0.0057783 -0.00035029
+ 7.9e+09Hz 0.00579806 -0.00036605
+ 8e+09Hz 0.00581785 -0.000382155
+ 8.1e+09Hz 0.00583767 -0.000398604
+ 8.2e+09Hz 0.00585751 -0.000415398
+ 8.3e+09Hz 0.00587736 -0.000432536
+ 8.4e+09Hz 0.00589721 -0.000450016
+ 8.5e+09Hz 0.00591707 -0.000467839
+ 8.6e+09Hz 0.00593692 -0.000486003
+ 8.7e+09Hz 0.00595676 -0.000504507
+ 8.8e+09Hz 0.00597658 -0.00052335
+ 8.9e+09Hz 0.00599638 -0.000542531
+ 9e+09Hz 0.00601615 -0.000562048
+ 9.1e+09Hz 0.00603589 -0.0005819
+ 9.2e+09Hz 0.00605558 -0.000602085
+ 9.3e+09Hz 0.00607523 -0.000622601
+ 9.4e+09Hz 0.00609483 -0.000643447
+ 9.5e+09Hz 0.00611437 -0.00066462
+ 9.6e+09Hz 0.00613384 -0.000686119
+ 9.7e+09Hz 0.00615324 -0.000707941
+ 9.8e+09Hz 0.00617257 -0.000730084
+ 9.9e+09Hz 0.00619183 -0.000752546
+ 1e+10Hz 0.00621099 -0.000775324
+ 1.01e+10Hz 0.00623007 -0.000798416
+ 1.02e+10Hz 0.00624905 -0.000821819
+ 1.03e+10Hz 0.00626793 -0.000845531
+ 1.04e+10Hz 0.0062867 -0.000869548
+ 1.05e+10Hz 0.00630536 -0.000893868
+ 1.06e+10Hz 0.00632391 -0.000918487
+ 1.07e+10Hz 0.00634234 -0.000943403
+ 1.08e+10Hz 0.00636064 -0.000968612
+ 1.09e+10Hz 0.00637881 -0.000994112
+ 1.1e+10Hz 0.00639685 -0.0010199
+ 1.11e+10Hz 0.00641475 -0.00104597
+ 1.12e+10Hz 0.00643251 -0.00107232
+ 1.13e+10Hz 0.00645012 -0.00109895
+ 1.14e+10Hz 0.00646758 -0.00112585
+ 1.15e+10Hz 0.00648489 -0.00115302
+ 1.16e+10Hz 0.00650203 -0.00118045
+ 1.17e+10Hz 0.00651902 -0.00120815
+ 1.18e+10Hz 0.00653583 -0.00123611
+ 1.19e+10Hz 0.00655248 -0.00126432
+ 1.2e+10Hz 0.00656895 -0.00129278
+ 1.21e+10Hz 0.00658524 -0.00132148
+ 1.22e+10Hz 0.00660135 -0.00135043
+ 1.23e+10Hz 0.00661728 -0.00137962
+ 1.24e+10Hz 0.00663302 -0.00140904
+ 1.25e+10Hz 0.00664857 -0.00143869
+ 1.26e+10Hz 0.00666392 -0.00146857
+ 1.27e+10Hz 0.00667908 -0.00149867
+ 1.28e+10Hz 0.00669404 -0.00152899
+ 1.29e+10Hz 0.00670879 -0.00155951
+ 1.3e+10Hz 0.00672335 -0.00159025
+ 1.31e+10Hz 0.00673769 -0.00162119
+ 1.32e+10Hz 0.00675182 -0.00165234
+ 1.33e+10Hz 0.00676574 -0.00168367
+ 1.34e+10Hz 0.00677945 -0.0017152
+ 1.35e+10Hz 0.00679294 -0.00174692
+ 1.36e+10Hz 0.00680621 -0.00177882
+ 1.37e+10Hz 0.00681926 -0.00181089
+ 1.38e+10Hz 0.00683208 -0.00184314
+ 1.39e+10Hz 0.00684468 -0.00187555
+ 1.4e+10Hz 0.00685706 -0.00190813
+ 1.41e+10Hz 0.00686921 -0.00194087
+ 1.42e+10Hz 0.00688113 -0.00197377
+ 1.43e+10Hz 0.00689282 -0.00200681
+ 1.44e+10Hz 0.00690427 -0.00204001
+ 1.45e+10Hz 0.0069155 -0.00207334
+ 1.46e+10Hz 0.00692649 -0.00210681
+ 1.47e+10Hz 0.00693724 -0.00214041
+ 1.48e+10Hz 0.00694776 -0.00217414
+ 1.49e+10Hz 0.00695804 -0.00220799
+ 1.5e+10Hz 0.00696809 -0.00224196
+ 1.51e+10Hz 0.0069779 -0.00227604
+ 1.52e+10Hz 0.00698746 -0.00231024
+ 1.53e+10Hz 0.00699679 -0.00234454
+ 1.54e+10Hz 0.00700588 -0.00237894
+ 1.55e+10Hz 0.00701474 -0.00241344
+ 1.56e+10Hz 0.00702335 -0.00244802
+ 1.57e+10Hz 0.00703172 -0.0024827
+ 1.58e+10Hz 0.00703985 -0.00251746
+ 1.59e+10Hz 0.00704774 -0.0025523
+ 1.6e+10Hz 0.0070554 -0.00258721
+ 1.61e+10Hz 0.00706281 -0.00262219
+ 1.62e+10Hz 0.00706999 -0.00265724
+ 1.63e+10Hz 0.00707693 -0.00269235
+ 1.64e+10Hz 0.00708363 -0.00272752
+ 1.65e+10Hz 0.00709009 -0.00276274
+ 1.66e+10Hz 0.00709632 -0.00279801
+ 1.67e+10Hz 0.00710231 -0.00283332
+ 1.68e+10Hz 0.00710806 -0.00286868
+ 1.69e+10Hz 0.00711359 -0.00290407
+ 1.7e+10Hz 0.00711888 -0.0029395
+ 1.71e+10Hz 0.00712393 -0.00297496
+ 1.72e+10Hz 0.00712876 -0.00301044
+ 1.73e+10Hz 0.00713336 -0.00304594
+ 1.74e+10Hz 0.00713773 -0.00308147
+ 1.75e+10Hz 0.00714187 -0.003117
+ 1.76e+10Hz 0.00714579 -0.00315255
+ 1.77e+10Hz 0.00714948 -0.0031881
+ 1.78e+10Hz 0.00715295 -0.00322366
+ 1.79e+10Hz 0.00715621 -0.00325922
+ 1.8e+10Hz 0.00715924 -0.00329477
+ 1.81e+10Hz 0.00716205 -0.00333032
+ 1.82e+10Hz 0.00716465 -0.00336586
+ 1.83e+10Hz 0.00716703 -0.00340138
+ 1.84e+10Hz 0.00716921 -0.00343689
+ 1.85e+10Hz 0.00717117 -0.00347238
+ 1.86e+10Hz 0.00717293 -0.00350784
+ 1.87e+10Hz 0.00717447 -0.00354328
+ 1.88e+10Hz 0.00717582 -0.00357869
+ 1.89e+10Hz 0.00717696 -0.00361407
+ 1.9e+10Hz 0.00717791 -0.00364941
+ 1.91e+10Hz 0.00717866 -0.00368472
+ 1.92e+10Hz 0.00717921 -0.00371999
+ 1.93e+10Hz 0.00717957 -0.00375522
+ 1.94e+10Hz 0.00717974 -0.0037904
+ 1.95e+10Hz 0.00717972 -0.00382553
+ 1.96e+10Hz 0.00717951 -0.00386061
+ 1.97e+10Hz 0.00717912 -0.00389564
+ 1.98e+10Hz 0.00717856 -0.00393062
+ 1.99e+10Hz 0.00717781 -0.00396554
+ 2e+10Hz 0.00717689 -0.0040004
+ 2.01e+10Hz 0.00717579 -0.0040352
+ 2.02e+10Hz 0.00717453 -0.00406994
+ 2.03e+10Hz 0.00717309 -0.00410461
+ 2.04e+10Hz 0.00717149 -0.00413921
+ 2.05e+10Hz 0.00716973 -0.00417375
+ 2.06e+10Hz 0.00716781 -0.00420822
+ 2.07e+10Hz 0.00716573 -0.00424261
+ 2.08e+10Hz 0.0071635 -0.00427693
+ 2.09e+10Hz 0.00716111 -0.00431118
+ 2.1e+10Hz 0.00715858 -0.00434535
+ 2.11e+10Hz 0.0071559 -0.00437944
+ 2.12e+10Hz 0.00715308 -0.00441345
+ 2.13e+10Hz 0.00715011 -0.00444738
+ 2.14e+10Hz 0.00714701 -0.00448123
+ 2.15e+10Hz 0.00714377 -0.004515
+ 2.16e+10Hz 0.0071404 -0.00454868
+ 2.17e+10Hz 0.0071369 -0.00458228
+ 2.18e+10Hz 0.00713327 -0.0046158
+ 2.19e+10Hz 0.00712952 -0.00464922
+ 2.2e+10Hz 0.00712565 -0.00468256
+ 2.21e+10Hz 0.00712165 -0.00471582
+ 2.22e+10Hz 0.00711755 -0.00474898
+ 2.23e+10Hz 0.00711332 -0.00478206
+ 2.24e+10Hz 0.00710899 -0.00481504
+ 2.25e+10Hz 0.00710455 -0.00484794
+ 2.26e+10Hz 0.00710001 -0.00488074
+ 2.27e+10Hz 0.00709536 -0.00491346
+ 2.28e+10Hz 0.00709061 -0.00494608
+ 2.29e+10Hz 0.00708577 -0.00497862
+ 2.3e+10Hz 0.00708083 -0.00501106
+ 2.31e+10Hz 0.00707579 -0.00504341
+ 2.32e+10Hz 0.00707067 -0.00507567
+ 2.33e+10Hz 0.00706546 -0.00510784
+ 2.34e+10Hz 0.00706017 -0.00513992
+ 2.35e+10Hz 0.0070548 -0.00517191
+ 2.36e+10Hz 0.00704934 -0.00520381
+ 2.37e+10Hz 0.00704381 -0.00523561
+ 2.38e+10Hz 0.00703821 -0.00526733
+ 2.39e+10Hz 0.00703253 -0.00529896
+ 2.4e+10Hz 0.00702678 -0.0053305
+ 2.41e+10Hz 0.00702097 -0.00536195
+ 2.42e+10Hz 0.00701509 -0.00539332
+ 2.43e+10Hz 0.00700915 -0.00542459
+ 2.44e+10Hz 0.00700315 -0.00545578
+ 2.45e+10Hz 0.00699709 -0.00548688
+ 2.46e+10Hz 0.00699097 -0.0055179
+ 2.47e+10Hz 0.0069848 -0.00554884
+ 2.48e+10Hz 0.00697857 -0.00557969
+ 2.49e+10Hz 0.0069723 -0.00561046
+ 2.5e+10Hz 0.00696598 -0.00564114
+ 2.51e+10Hz 0.00695961 -0.00567175
+ 2.52e+10Hz 0.0069532 -0.00570228
+ 2.53e+10Hz 0.00694675 -0.00573272
+ 2.54e+10Hz 0.00694026 -0.00576309
+ 2.55e+10Hz 0.00693372 -0.00579339
+ 2.56e+10Hz 0.00692716 -0.00582361
+ 2.57e+10Hz 0.00692055 -0.00585375
+ 2.58e+10Hz 0.00691392 -0.00588382
+ 2.59e+10Hz 0.00690725 -0.00591382
+ 2.6e+10Hz 0.00690055 -0.00594375
+ 2.61e+10Hz 0.00689382 -0.00597361
+ 2.62e+10Hz 0.00688707 -0.0060034
+ 2.63e+10Hz 0.00688029 -0.00603313
+ 2.64e+10Hz 0.00687348 -0.00606279
+ 2.65e+10Hz 0.00686665 -0.00609239
+ 2.66e+10Hz 0.0068598 -0.00612192
+ 2.67e+10Hz 0.00685293 -0.00615139
+ 2.68e+10Hz 0.00684605 -0.00618081
+ 2.69e+10Hz 0.00683914 -0.00621016
+ 2.7e+10Hz 0.00683221 -0.00623947
+ 2.71e+10Hz 0.00682527 -0.00626871
+ 2.72e+10Hz 0.00681832 -0.0062979
+ 2.73e+10Hz 0.00681135 -0.00632704
+ 2.74e+10Hz 0.00680436 -0.00635613
+ 2.75e+10Hz 0.00679737 -0.00638517
+ 2.76e+10Hz 0.00679036 -0.00641417
+ 2.77e+10Hz 0.00678335 -0.00644311
+ 2.78e+10Hz 0.00677632 -0.00647202
+ 2.79e+10Hz 0.00676928 -0.00650088
+ 2.8e+10Hz 0.00676224 -0.0065297
+ 2.81e+10Hz 0.00675518 -0.00655848
+ 2.82e+10Hz 0.00674812 -0.00658722
+ 2.83e+10Hz 0.00674105 -0.00661593
+ 2.84e+10Hz 0.00673398 -0.0066446
+ 2.85e+10Hz 0.00672689 -0.00667324
+ 2.86e+10Hz 0.0067198 -0.00670184
+ 2.87e+10Hz 0.00671271 -0.00673042
+ 2.88e+10Hz 0.00670561 -0.00675897
+ 2.89e+10Hz 0.00669851 -0.00678749
+ 2.9e+10Hz 0.00669139 -0.00681599
+ 2.91e+10Hz 0.00668428 -0.00684446
+ 2.92e+10Hz 0.00667716 -0.00687291
+ 2.93e+10Hz 0.00667003 -0.00690134
+ 2.94e+10Hz 0.0066629 -0.00692975
+ 2.95e+10Hz 0.00665576 -0.00695814
+ 2.96e+10Hz 0.00664862 -0.00698652
+ 2.97e+10Hz 0.00664148 -0.00701488
+ 2.98e+10Hz 0.00663432 -0.00704322
+ 2.99e+10Hz 0.00662716 -0.00707156
+ 3e+10Hz 0.00662 -0.00709988
+ 3.01e+10Hz 0.00661283 -0.0071282
+ 3.02e+10Hz 0.00660565 -0.00715651
+ 3.03e+10Hz 0.00659846 -0.00718481
+ 3.04e+10Hz 0.00659127 -0.0072131
+ 3.05e+10Hz 0.00658407 -0.00724139
+ 3.06e+10Hz 0.00657686 -0.00726968
+ 3.07e+10Hz 0.00656964 -0.00729797
+ 3.08e+10Hz 0.00656241 -0.00732626
+ 3.09e+10Hz 0.00655517 -0.00735454
+ 3.1e+10Hz 0.00654792 -0.00738283
+ 3.11e+10Hz 0.00654066 -0.00741113
+ 3.12e+10Hz 0.00653339 -0.00743943
+ 3.13e+10Hz 0.0065261 -0.00746773
+ 3.14e+10Hz 0.0065188 -0.00749604
+ 3.15e+10Hz 0.00651149 -0.00752436
+ 3.16e+10Hz 0.00650416 -0.00755268
+ 3.17e+10Hz 0.00649682 -0.00758102
+ 3.18e+10Hz 0.00648946 -0.00760937
+ 3.19e+10Hz 0.00648208 -0.00763772
+ 3.2e+10Hz 0.00647468 -0.00766609
+ 3.21e+10Hz 0.00646726 -0.00769448
+ 3.22e+10Hz 0.00645983 -0.00772288
+ 3.23e+10Hz 0.00645237 -0.00775129
+ 3.24e+10Hz 0.00644489 -0.00777972
+ 3.25e+10Hz 0.00643738 -0.00780816
+ 3.26e+10Hz 0.00642986 -0.00783662
+ 3.27e+10Hz 0.0064223 -0.0078651
+ 3.28e+10Hz 0.00641473 -0.0078936
+ 3.29e+10Hz 0.00640712 -0.00792212
+ 3.3e+10Hz 0.00639949 -0.00795065
+ 3.31e+10Hz 0.00639182 -0.00797921
+ 3.32e+10Hz 0.00638413 -0.00800779
+ 3.33e+10Hz 0.00637641 -0.00803639
+ 3.34e+10Hz 0.00636865 -0.008065
+ 3.35e+10Hz 0.00636086 -0.00809365
+ 3.36e+10Hz 0.00635303 -0.00812231
+ 3.37e+10Hz 0.00634517 -0.008151
+ 3.38e+10Hz 0.00633728 -0.0081797
+ 3.39e+10Hz 0.00632934 -0.00820844
+ 3.4e+10Hz 0.00632137 -0.00823719
+ 3.41e+10Hz 0.00631335 -0.00826597
+ 3.42e+10Hz 0.0063053 -0.00829477
+ 3.43e+10Hz 0.0062972 -0.0083236
+ 3.44e+10Hz 0.00628906 -0.00835245
+ 3.45e+10Hz 0.00628087 -0.00838133
+ 3.46e+10Hz 0.00627264 -0.00841022
+ 3.47e+10Hz 0.00626436 -0.00843915
+ 3.48e+10Hz 0.00625603 -0.00846809
+ 3.49e+10Hz 0.00624766 -0.00849706
+ 3.5e+10Hz 0.00623923 -0.00852606
+ 3.51e+10Hz 0.00623075 -0.00855508
+ 3.52e+10Hz 0.00622222 -0.00858412
+ 3.53e+10Hz 0.00621364 -0.00861318
+ 3.54e+10Hz 0.006205 -0.00864227
+ 3.55e+10Hz 0.00619631 -0.00867138
+ 3.56e+10Hz 0.00618756 -0.00870052
+ 3.57e+10Hz 0.00617875 -0.00872968
+ 3.58e+10Hz 0.00616989 -0.00875885
+ 3.59e+10Hz 0.00616096 -0.00878805
+ 3.6e+10Hz 0.00615198 -0.00881728
+ 3.61e+10Hz 0.00614293 -0.00884652
+ 3.62e+10Hz 0.00613382 -0.00887578
+ 3.63e+10Hz 0.00612464 -0.00890507
+ 3.64e+10Hz 0.00611541 -0.00893437
+ 3.65e+10Hz 0.0061061 -0.00896369
+ 3.66e+10Hz 0.00609673 -0.00899303
+ 3.67e+10Hz 0.00608729 -0.00902239
+ 3.68e+10Hz 0.00607778 -0.00905177
+ 3.69e+10Hz 0.00606821 -0.00908116
+ 3.7e+10Hz 0.00605856 -0.00911057
+ 3.71e+10Hz 0.00604885 -0.00913999
+ 3.72e+10Hz 0.00603906 -0.00916943
+ 3.73e+10Hz 0.0060292 -0.00919888
+ 3.74e+10Hz 0.00601926 -0.00922835
+ 3.75e+10Hz 0.00600926 -0.00925783
+ 3.76e+10Hz 0.00599917 -0.00928732
+ 3.77e+10Hz 0.00598901 -0.00931682
+ 3.78e+10Hz 0.00597878 -0.00934633
+ 3.79e+10Hz 0.00596847 -0.00937585
+ 3.8e+10Hz 0.00595808 -0.00940538
+ 3.81e+10Hz 0.00594761 -0.00943492
+ 3.82e+10Hz 0.00593707 -0.00946447
+ 3.83e+10Hz 0.00592644 -0.00949402
+ 3.84e+10Hz 0.00591574 -0.00952358
+ 3.85e+10Hz 0.00590495 -0.00955314
+ 3.86e+10Hz 0.00589408 -0.0095827
+ 3.87e+10Hz 0.00588314 -0.00961227
+ 3.88e+10Hz 0.00587211 -0.00964184
+ 3.89e+10Hz 0.00586099 -0.00967141
+ 3.9e+10Hz 0.0058498 -0.00970098
+ 3.91e+10Hz 0.00583852 -0.00973055
+ 3.92e+10Hz 0.00582716 -0.00976011
+ 3.93e+10Hz 0.00581571 -0.00978968
+ 3.94e+10Hz 0.00580418 -0.00981924
+ 3.95e+10Hz 0.00579257 -0.00984879
+ 3.96e+10Hz 0.00578087 -0.00987834
+ 3.97e+10Hz 0.00576908 -0.00990788
+ 3.98e+10Hz 0.00575722 -0.00993741
+ 3.99e+10Hz 0.00574526 -0.00996694
+ 4e+10Hz 0.00573322 -0.00999645
+ 4.01e+10Hz 0.00572109 -0.010026
+ 4.02e+10Hz 0.00570888 -0.0100554
+ 4.03e+10Hz 0.00569658 -0.0100849
+ 4.04e+10Hz 0.00568419 -0.0101144
+ 4.05e+10Hz 0.00567172 -0.0101438
+ 4.06e+10Hz 0.00565916 -0.0101733
+ 4.07e+10Hz 0.00564652 -0.0102027
+ 4.08e+10Hz 0.00563379 -0.0102321
+ 4.09e+10Hz 0.00562097 -0.0102615
+ 4.1e+10Hz 0.00560807 -0.0102908
+ 4.11e+10Hz 0.00559508 -0.0103202
+ 4.12e+10Hz 0.00558201 -0.0103495
+ 4.13e+10Hz 0.00556884 -0.0103788
+ 4.14e+10Hz 0.0055556 -0.010408
+ 4.15e+10Hz 0.00554227 -0.0104373
+ 4.16e+10Hz 0.00552885 -0.0104665
+ 4.17e+10Hz 0.00551534 -0.0104957
+ 4.18e+10Hz 0.00550176 -0.0105248
+ 4.19e+10Hz 0.00548809 -0.010554
+ 4.2e+10Hz 0.00547433 -0.0105831
+ 4.21e+10Hz 0.00546049 -0.0106121
+ 4.22e+10Hz 0.00544656 -0.0106412
+ 4.23e+10Hz 0.00543256 -0.0106702
+ 4.24e+10Hz 0.00541846 -0.0106992
+ 4.25e+10Hz 0.00540429 -0.0107281
+ 4.26e+10Hz 0.00539004 -0.010757
+ 4.27e+10Hz 0.0053757 -0.0107859
+ 4.28e+10Hz 0.00536128 -0.0108147
+ 4.29e+10Hz 0.00534678 -0.0108435
+ 4.3e+10Hz 0.0053322 -0.0108723
+ 4.31e+10Hz 0.00531754 -0.010901
+ 4.32e+10Hz 0.0053028 -0.0109297
+ 4.33e+10Hz 0.00528798 -0.0109583
+ 4.34e+10Hz 0.00527308 -0.0109869
+ 4.35e+10Hz 0.00525811 -0.0110154
+ 4.36e+10Hz 0.00524306 -0.0110439
+ 4.37e+10Hz 0.00522793 -0.0110724
+ 4.38e+10Hz 0.00521272 -0.0111008
+ 4.39e+10Hz 0.00519744 -0.0111292
+ 4.4e+10Hz 0.00518209 -0.0111575
+ 4.41e+10Hz 0.00516666 -0.0111858
+ 4.42e+10Hz 0.00515116 -0.011214
+ 4.43e+10Hz 0.00513558 -0.0112422
+ 4.44e+10Hz 0.00511993 -0.0112703
+ 4.45e+10Hz 0.00510421 -0.0112984
+ 4.46e+10Hz 0.00508842 -0.0113265
+ 4.47e+10Hz 0.00507256 -0.0113545
+ 4.48e+10Hz 0.00505663 -0.0113824
+ 4.49e+10Hz 0.00504063 -0.0114103
+ 4.5e+10Hz 0.00502457 -0.0114381
+ 4.51e+10Hz 0.00500843 -0.0114659
+ 4.52e+10Hz 0.00499223 -0.0114936
+ 4.53e+10Hz 0.00497597 -0.0115213
+ 4.54e+10Hz 0.00495964 -0.0115489
+ 4.55e+10Hz 0.00494324 -0.0115765
+ 4.56e+10Hz 0.00492678 -0.011604
+ 4.57e+10Hz 0.00491026 -0.0116314
+ 4.58e+10Hz 0.00489368 -0.0116588
+ 4.59e+10Hz 0.00487703 -0.0116862
+ 4.6e+10Hz 0.00486033 -0.0117135
+ 4.61e+10Hz 0.00484356 -0.0117407
+ 4.62e+10Hz 0.00482674 -0.0117679
+ 4.63e+10Hz 0.00480986 -0.011795
+ 4.64e+10Hz 0.00479292 -0.011822
+ 4.65e+10Hz 0.00477592 -0.011849
+ 4.66e+10Hz 0.00475887 -0.011876
+ 4.67e+10Hz 0.00474177 -0.0119029
+ 4.68e+10Hz 0.00472461 -0.0119297
+ 4.69e+10Hz 0.0047074 -0.0119565
+ 4.7e+10Hz 0.00469013 -0.0119832
+ 4.71e+10Hz 0.00467281 -0.0120098
+ 4.72e+10Hz 0.00465544 -0.0120364
+ 4.73e+10Hz 0.00463803 -0.012063
+ 4.74e+10Hz 0.00462056 -0.0120895
+ 4.75e+10Hz 0.00460304 -0.0121159
+ 4.76e+10Hz 0.00458548 -0.0121422
+ 4.77e+10Hz 0.00456787 -0.0121685
+ 4.78e+10Hz 0.00455021 -0.0121948
+ 4.79e+10Hz 0.00453251 -0.012221
+ 4.8e+10Hz 0.00451476 -0.0122471
+ 4.81e+10Hz 0.00449697 -0.0122732
+ 4.82e+10Hz 0.00447914 -0.0122992
+ 4.83e+10Hz 0.00446126 -0.0123251
+ 4.84e+10Hz 0.00444334 -0.012351
+ 4.85e+10Hz 0.00442538 -0.0123769
+ 4.86e+10Hz 0.00440738 -0.0124027
+ 4.87e+10Hz 0.00438934 -0.0124284
+ 4.88e+10Hz 0.00437126 -0.0124541
+ 4.89e+10Hz 0.00435314 -0.0124797
+ 4.9e+10Hz 0.00433498 -0.0125052
+ 4.91e+10Hz 0.00431679 -0.0125307
+ 4.92e+10Hz 0.00429856 -0.0125561
+ 4.93e+10Hz 0.0042803 -0.0125815
+ 4.94e+10Hz 0.004262 -0.0126068
+ 4.95e+10Hz 0.00424366 -0.0126321
+ 4.96e+10Hz 0.00422529 -0.0126573
+ 4.97e+10Hz 0.00420689 -0.0126825
+ 4.98e+10Hz 0.00418846 -0.0127076
+ 4.99e+10Hz 0.00416999 -0.0127326
+ 5e+10Hz 0.00415149 -0.0127576
+ 5.01e+10Hz 0.00413296 -0.0127826
+ 5.02e+10Hz 0.0041144 -0.0128074
+ 5.03e+10Hz 0.00409581 -0.0128323
+ 5.04e+10Hz 0.00407719 -0.0128571
+ 5.05e+10Hz 0.00405854 -0.0128818
+ 5.06e+10Hz 0.00403987 -0.0129065
+ 5.07e+10Hz 0.00402116 -0.0129311
+ 5.08e+10Hz 0.00400243 -0.0129556
+ 5.09e+10Hz 0.00398367 -0.0129802
+ 5.1e+10Hz 0.00396488 -0.0130046
+ 5.11e+10Hz 0.00394607 -0.013029
+ 5.12e+10Hz 0.00392723 -0.0130534
+ 5.13e+10Hz 0.00390836 -0.0130777
+ 5.14e+10Hz 0.00388947 -0.013102
+ 5.15e+10Hz 0.00387056 -0.0131262
+ 5.16e+10Hz 0.00385162 -0.0131504
+ 5.17e+10Hz 0.00383265 -0.0131745
+ 5.18e+10Hz 0.00381367 -0.0131986
+ 5.19e+10Hz 0.00379466 -0.0132226
+ 5.2e+10Hz 0.00377562 -0.0132466
+ 5.21e+10Hz 0.00375656 -0.0132705
+ 5.22e+10Hz 0.00373748 -0.0132944
+ 5.23e+10Hz 0.00371838 -0.0133183
+ 5.24e+10Hz 0.00369925 -0.0133421
+ 5.25e+10Hz 0.00368011 -0.0133658
+ 5.26e+10Hz 0.00366094 -0.0133896
+ 5.27e+10Hz 0.00364175 -0.0134132
+ 5.28e+10Hz 0.00362253 -0.0134369
+ 5.29e+10Hz 0.0036033 -0.0134604
+ 5.3e+10Hz 0.00358404 -0.013484
+ 5.31e+10Hz 0.00356477 -0.0135075
+ 5.32e+10Hz 0.00354547 -0.013531
+ 5.33e+10Hz 0.00352615 -0.0135544
+ 5.34e+10Hz 0.00350681 -0.0135778
+ 5.35e+10Hz 0.00348745 -0.0136011
+ 5.36e+10Hz 0.00346807 -0.0136244
+ 5.37e+10Hz 0.00344867 -0.0136477
+ 5.38e+10Hz 0.00342925 -0.0136709
+ 5.39e+10Hz 0.0034098 -0.0136941
+ 5.4e+10Hz 0.00339034 -0.0137172
+ 5.41e+10Hz 0.00337085 -0.0137403
+ 5.42e+10Hz 0.00335135 -0.0137634
+ 5.43e+10Hz 0.00333182 -0.0137865
+ 5.44e+10Hz 0.00331228 -0.0138095
+ 5.45e+10Hz 0.00329271 -0.0138324
+ 5.46e+10Hz 0.00327312 -0.0138554
+ 5.47e+10Hz 0.00325351 -0.0138783
+ 5.48e+10Hz 0.00323388 -0.0139011
+ 5.49e+10Hz 0.00321423 -0.013924
+ 5.5e+10Hz 0.00319455 -0.0139468
+ 5.51e+10Hz 0.00317486 -0.0139695
+ 5.52e+10Hz 0.00315514 -0.0139923
+ 5.53e+10Hz 0.0031354 -0.014015
+ 5.54e+10Hz 0.00311564 -0.0140376
+ 5.55e+10Hz 0.00309586 -0.0140603
+ 5.56e+10Hz 0.00307606 -0.0140829
+ 5.57e+10Hz 0.00305623 -0.0141055
+ 5.58e+10Hz 0.00303638 -0.014128
+ 5.59e+10Hz 0.00301651 -0.0141505
+ 5.6e+10Hz 0.00299662 -0.014173
+ 5.61e+10Hz 0.0029767 -0.0141955
+ 5.62e+10Hz 0.00295676 -0.0142179
+ 5.63e+10Hz 0.00293679 -0.0142403
+ 5.64e+10Hz 0.0029168 -0.0142626
+ 5.65e+10Hz 0.00289679 -0.014285
+ 5.66e+10Hz 0.00287675 -0.0143073
+ 5.67e+10Hz 0.00285669 -0.0143296
+ 5.68e+10Hz 0.0028366 -0.0143518
+ 5.69e+10Hz 0.00281649 -0.014374
+ 5.7e+10Hz 0.00279635 -0.0143962
+ 5.71e+10Hz 0.00277619 -0.0144184
+ 5.72e+10Hz 0.002756 -0.0144406
+ 5.73e+10Hz 0.00273579 -0.0144627
+ 5.74e+10Hz 0.00271554 -0.0144848
+ 5.75e+10Hz 0.00269527 -0.0145068
+ 5.76e+10Hz 0.00267498 -0.0145288
+ 5.77e+10Hz 0.00265465 -0.0145509
+ 5.78e+10Hz 0.0026343 -0.0145728
+ 5.79e+10Hz 0.00261392 -0.0145948
+ 5.8e+10Hz 0.00259351 -0.0146167
+ 5.81e+10Hz 0.00257308 -0.0146386
+ 5.82e+10Hz 0.00255261 -0.0146605
+ 5.83e+10Hz 0.00253212 -0.0146823
+ 5.84e+10Hz 0.00251159 -0.0147042
+ 5.85e+10Hz 0.00249104 -0.014726
+ 5.86e+10Hz 0.00247045 -0.0147477
+ 5.87e+10Hz 0.00244984 -0.0147695
+ 5.88e+10Hz 0.00242919 -0.0147912
+ 5.89e+10Hz 0.00240851 -0.0148129
+ 5.9e+10Hz 0.00238781 -0.0148345
+ 5.91e+10Hz 0.00236707 -0.0148562
+ 5.92e+10Hz 0.00234629 -0.0148778
+ 5.93e+10Hz 0.00232549 -0.0148994
+ 5.94e+10Hz 0.00230465 -0.0149209
+ 5.95e+10Hz 0.00228378 -0.0149425
+ 5.96e+10Hz 0.00226287 -0.014964
+ 5.97e+10Hz 0.00224194 -0.0149854
+ 5.98e+10Hz 0.00222096 -0.0150069
+ 5.99e+10Hz 0.00219996 -0.0150283
+ 6e+10Hz 0.00217892 -0.0150497
+ 6.01e+10Hz 0.00215784 -0.0150711
+ 6.02e+10Hz 0.00213673 -0.0150924
+ 6.03e+10Hz 0.00211559 -0.0151137
+ 6.04e+10Hz 0.00209441 -0.015135
+ 6.05e+10Hz 0.00207319 -0.0151563
+ 6.06e+10Hz 0.00205194 -0.0151775
+ 6.07e+10Hz 0.00203065 -0.0151987
+ 6.08e+10Hz 0.00200932 -0.0152199
+ 6.09e+10Hz 0.00198796 -0.015241
+ 6.1e+10Hz 0.00196656 -0.0152621
+ 6.11e+10Hz 0.00194512 -0.0152832
+ 6.12e+10Hz 0.00192364 -0.0153043
+ 6.13e+10Hz 0.00190213 -0.0153253
+ 6.14e+10Hz 0.00188058 -0.0153463
+ 6.15e+10Hz 0.00185899 -0.0153672
+ 6.16e+10Hz 0.00183736 -0.0153882
+ 6.17e+10Hz 0.0018157 -0.0154091
+ 6.18e+10Hz 0.00179399 -0.0154299
+ 6.19e+10Hz 0.00177225 -0.0154508
+ 6.2e+10Hz 0.00175047 -0.0154716
+ 6.21e+10Hz 0.00172865 -0.0154924
+ 6.22e+10Hz 0.00170678 -0.0155131
+ 6.23e+10Hz 0.00168488 -0.0155338
+ 6.24e+10Hz 0.00166294 -0.0155545
+ 6.25e+10Hz 0.00164096 -0.0155751
+ 6.26e+10Hz 0.00161894 -0.0155957
+ 6.27e+10Hz 0.00159688 -0.0156163
+ 6.28e+10Hz 0.00157478 -0.0156368
+ 6.29e+10Hz 0.00155264 -0.0156574
+ 6.3e+10Hz 0.00153046 -0.0156778
+ 6.31e+10Hz 0.00150824 -0.0156983
+ 6.32e+10Hz 0.00148597 -0.0157187
+ 6.33e+10Hz 0.00146367 -0.015739
+ 6.34e+10Hz 0.00144133 -0.0157593
+ 6.35e+10Hz 0.00141894 -0.0157796
+ 6.36e+10Hz 0.00139652 -0.0157999
+ 6.37e+10Hz 0.00137405 -0.0158201
+ 6.38e+10Hz 0.00135155 -0.0158403
+ 6.39e+10Hz 0.001329 -0.0158604
+ 6.4e+10Hz 0.00130641 -0.0158805
+ 6.41e+10Hz 0.00128378 -0.0159006
+ 6.42e+10Hz 0.00126111 -0.0159206
+ 6.43e+10Hz 0.00123841 -0.0159406
+ 6.44e+10Hz 0.00121566 -0.0159605
+ 6.45e+10Hz 0.00119286 -0.0159804
+ 6.46e+10Hz 0.00117003 -0.0160003
+ 6.47e+10Hz 0.00114716 -0.0160201
+ 6.48e+10Hz 0.00112425 -0.0160399
+ 6.49e+10Hz 0.0011013 -0.0160596
+ 6.5e+10Hz 0.0010783 -0.0160793
+ 6.51e+10Hz 0.00105527 -0.0160989
+ 6.52e+10Hz 0.0010322 -0.0161185
+ 6.53e+10Hz 0.00100909 -0.0161381
+ 6.54e+10Hz 0.000985935 -0.0161576
+ 6.55e+10Hz 0.000962743 -0.0161771
+ 6.56e+10Hz 0.000939512 -0.0161965
+ 6.57e+10Hz 0.000916242 -0.0162159
+ 6.58e+10Hz 0.000892933 -0.0162352
+ 6.59e+10Hz 0.000869584 -0.0162545
+ 6.6e+10Hz 0.000846197 -0.0162737
+ 6.61e+10Hz 0.000822772 -0.0162929
+ 6.62e+10Hz 0.000799308 -0.0163121
+ 6.63e+10Hz 0.000775805 -0.0163312
+ 6.64e+10Hz 0.000752265 -0.0163502
+ 6.65e+10Hz 0.000728688 -0.0163693
+ 6.66e+10Hz 0.000705072 -0.0163882
+ 6.67e+10Hz 0.00068142 -0.0164071
+ 6.68e+10Hz 0.00065773 -0.016426
+ 6.69e+10Hz 0.000634004 -0.0164448
+ 6.7e+10Hz 0.000610241 -0.0164636
+ 6.71e+10Hz 0.000586442 -0.0164823
+ 6.72e+10Hz 0.000562607 -0.0165009
+ 6.73e+10Hz 0.000538736 -0.0165195
+ 6.74e+10Hz 0.00051483 -0.0165381
+ 6.75e+10Hz 0.000490889 -0.0165566
+ 6.76e+10Hz 0.000466913 -0.0165751
+ 6.77e+10Hz 0.000442902 -0.0165935
+ 6.78e+10Hz 0.000418857 -0.0166118
+ 6.79e+10Hz 0.000394778 -0.0166301
+ 6.8e+10Hz 0.000370666 -0.0166484
+ 6.81e+10Hz 0.00034652 -0.0166666
+ 6.82e+10Hz 0.000322341 -0.0166847
+ 6.83e+10Hz 0.00029813 -0.0167028
+ 6.84e+10Hz 0.000273886 -0.0167209
+ 6.85e+10Hz 0.000249611 -0.0167388
+ 6.86e+10Hz 0.000225304 -0.0167568
+ 6.87e+10Hz 0.000200965 -0.0167747
+ 6.88e+10Hz 0.000176596 -0.0167925
+ 6.89e+10Hz 0.000152196 -0.0168102
+ 6.9e+10Hz 0.000127766 -0.016828
+ 6.91e+10Hz 0.000103306 -0.0168456
+ 6.92e+10Hz 7.88161e-05 -0.0168632
+ 6.93e+10Hz 5.42975e-05 -0.0168808
+ 6.94e+10Hz 2.97502e-05 -0.0168983
+ 6.95e+10Hz 5.17445e-06 -0.0169157
+ 6.96e+10Hz -1.94293e-05 -0.0169331
+ 6.97e+10Hz -4.40606e-05 -0.0169504
+ 6.98e+10Hz -6.87192e-05 -0.0169677
+ 6.99e+10Hz -9.34047e-05 -0.0169849
+ 7e+10Hz -0.000118117 -0.0170021
+ 7.01e+10Hz -0.000142855 -0.0170192
+ 7.02e+10Hz -0.000167619 -0.0170362
+ 7.03e+10Hz -0.000192408 -0.0170532
+ 7.04e+10Hz -0.000217222 -0.0170701
+ 7.05e+10Hz -0.00024206 -0.017087
+ 7.06e+10Hz -0.000266923 -0.0171039
+ 7.07e+10Hz -0.00029181 -0.0171206
+ 7.08e+10Hz -0.00031672 -0.0171373
+ 7.09e+10Hz -0.000341654 -0.017154
+ 7.1e+10Hz -0.000366609 -0.0171706
+ 7.11e+10Hz -0.000391588 -0.0171871
+ 7.12e+10Hz -0.000416588 -0.0172036
+ 7.13e+10Hz -0.000441609 -0.01722
+ 7.14e+10Hz -0.000466652 -0.0172364
+ 7.15e+10Hz -0.000491716 -0.0172527
+ 7.16e+10Hz -0.0005168 -0.017269
+ 7.17e+10Hz -0.000541904 -0.0172852
+ 7.18e+10Hz -0.000567028 -0.0173013
+ 7.19e+10Hz -0.000592171 -0.0173174
+ 7.2e+10Hz -0.000617333 -0.0173335
+ 7.21e+10Hz -0.000642514 -0.0173494
+ 7.22e+10Hz -0.000667713 -0.0173654
+ 7.23e+10Hz -0.000692929 -0.0173812
+ 7.24e+10Hz -0.000718164 -0.017397
+ 7.25e+10Hz -0.000743415 -0.0174128
+ 7.26e+10Hz -0.000768684 -0.0174285
+ 7.27e+10Hz -0.000793969 -0.0174441
+ 7.28e+10Hz -0.00081927 -0.0174597
+ 7.29e+10Hz -0.000844587 -0.0174752
+ 7.3e+10Hz -0.000869919 -0.0174907
+ 7.31e+10Hz -0.000895267 -0.0175061
+ 7.32e+10Hz -0.000920629 -0.0175215
+ 7.33e+10Hz -0.000946006 -0.0175368
+ 7.34e+10Hz -0.000971398 -0.017552
+ 7.35e+10Hz -0.000996803 -0.0175672
+ 7.36e+10Hz -0.00102222 -0.0175824
+ 7.37e+10Hz -0.00104765 -0.0175975
+ 7.38e+10Hz -0.0010731 -0.0176125
+ 7.39e+10Hz -0.00109856 -0.0176275
+ 7.4e+10Hz -0.00112403 -0.0176424
+ 7.41e+10Hz -0.00114951 -0.0176573
+ 7.42e+10Hz -0.00117501 -0.0176721
+ 7.43e+10Hz -0.00120051 -0.0176869
+ 7.44e+10Hz -0.00122603 -0.0177016
+ 7.45e+10Hz -0.00125156 -0.0177162
+ 7.46e+10Hz -0.0012771 -0.0177308
+ 7.47e+10Hz -0.00130265 -0.0177454
+ 7.48e+10Hz -0.00132821 -0.0177599
+ 7.49e+10Hz -0.00135379 -0.0177743
+ 7.5e+10Hz -0.00137937 -0.0177887
+ 7.51e+10Hz -0.00140496 -0.0178031
+ 7.52e+10Hz -0.00143056 -0.0178174
+ 7.53e+10Hz -0.00145617 -0.0178316
+ 7.54e+10Hz -0.00148179 -0.0178458
+ 7.55e+10Hz -0.00150742 -0.0178599
+ 7.56e+10Hz -0.00153306 -0.017874
+ 7.57e+10Hz -0.00155871 -0.0178881
+ 7.58e+10Hz -0.00158436 -0.0179021
+ 7.59e+10Hz -0.00161003 -0.017916
+ 7.6e+10Hz -0.0016357 -0.0179299
+ 7.61e+10Hz -0.00166138 -0.0179437
+ 7.62e+10Hz -0.00168707 -0.0179575
+ 7.63e+10Hz -0.00171277 -0.0179712
+ 7.64e+10Hz -0.00173847 -0.0179849
+ 7.65e+10Hz -0.00176418 -0.0179986
+ 7.66e+10Hz -0.0017899 -0.0180121
+ 7.67e+10Hz -0.00181563 -0.0180257
+ 7.68e+10Hz -0.00184136 -0.0180392
+ 7.69e+10Hz -0.0018671 -0.0180526
+ 7.7e+10Hz -0.00189285 -0.018066
+ 7.71e+10Hz -0.00191861 -0.0180794
+ 7.72e+10Hz -0.00194437 -0.0180927
+ 7.73e+10Hz -0.00197014 -0.0181059
+ 7.74e+10Hz -0.00199592 -0.0181191
+ 7.75e+10Hz -0.0020217 -0.0181323
+ 7.76e+10Hz -0.00204749 -0.0181454
+ 7.77e+10Hz -0.00207328 -0.0181585
+ 7.78e+10Hz -0.00209909 -0.0181715
+ 7.79e+10Hz -0.0021249 -0.0181845
+ 7.8e+10Hz -0.00215071 -0.0181974
+ 7.81e+10Hz -0.00217654 -0.0182103
+ 7.82e+10Hz -0.00220237 -0.0182231
+ 7.83e+10Hz -0.0022282 -0.0182359
+ 7.84e+10Hz -0.00225405 -0.0182487
+ 7.85e+10Hz -0.0022799 -0.0182614
+ 7.86e+10Hz -0.00230575 -0.018274
+ 7.87e+10Hz -0.00233162 -0.0182867
+ 7.88e+10Hz -0.00235749 -0.0182992
+ 7.89e+10Hz -0.00238336 -0.0183118
+ 7.9e+10Hz -0.00240925 -0.0183242
+ 7.91e+10Hz -0.00243514 -0.0183367
+ 7.92e+10Hz -0.00246103 -0.0183491
+ 7.93e+10Hz -0.00248694 -0.0183614
+ 7.94e+10Hz -0.00251285 -0.0183737
+ 7.95e+10Hz -0.00253876 -0.018386
+ 7.96e+10Hz -0.00256469 -0.0183982
+ 7.97e+10Hz -0.00259062 -0.0184104
+ 7.98e+10Hz -0.00261656 -0.0184226
+ 7.99e+10Hz -0.00264251 -0.0184347
+ 8e+10Hz -0.00266846 -0.0184467
+ 8.01e+10Hz -0.00269442 -0.0184587
+ 8.02e+10Hz -0.00272039 -0.0184707
+ 8.03e+10Hz -0.00274637 -0.0184826
+ 8.04e+10Hz -0.00277235 -0.0184945
+ 8.05e+10Hz -0.00279834 -0.0185064
+ 8.06e+10Hz -0.00282434 -0.0185182
+ 8.07e+10Hz -0.00285035 -0.0185299
+ 8.08e+10Hz -0.00287637 -0.0185417
+ 8.09e+10Hz -0.00290239 -0.0185534
+ 8.1e+10Hz -0.00292842 -0.018565
+ 8.11e+10Hz -0.00295446 -0.0185766
+ 8.12e+10Hz -0.00298051 -0.0185882
+ 8.13e+10Hz -0.00300657 -0.0185997
+ 8.14e+10Hz -0.00303264 -0.0186111
+ 8.15e+10Hz -0.00305872 -0.0186226
+ 8.16e+10Hz -0.0030848 -0.018634
+ 8.17e+10Hz -0.00311089 -0.0186453
+ 8.18e+10Hz -0.003137 -0.0186567
+ 8.19e+10Hz -0.00316311 -0.0186679
+ 8.2e+10Hz -0.00318923 -0.0186792
+ 8.21e+10Hz -0.00321537 -0.0186904
+ 8.22e+10Hz -0.00324151 -0.0187015
+ 8.23e+10Hz -0.00326766 -0.0187126
+ 8.24e+10Hz -0.00329382 -0.0187237
+ 8.25e+10Hz -0.00332 -0.0187347
+ 8.26e+10Hz -0.00334618 -0.0187457
+ 8.27e+10Hz -0.00337237 -0.0187567
+ 8.28e+10Hz -0.00339858 -0.0187676
+ 8.29e+10Hz -0.00342479 -0.0187784
+ 8.3e+10Hz -0.00345102 -0.0187893
+ 8.31e+10Hz -0.00347725 -0.0188001
+ 8.32e+10Hz -0.0035035 -0.0188108
+ 8.33e+10Hz -0.00352976 -0.0188215
+ 8.34e+10Hz -0.00355603 -0.0188322
+ 8.35e+10Hz -0.00358231 -0.0188428
+ 8.36e+10Hz -0.00360861 -0.0188534
+ 8.37e+10Hz -0.00363491 -0.0188639
+ 8.38e+10Hz -0.00366123 -0.0188744
+ 8.39e+10Hz -0.00368756 -0.0188849
+ 8.4e+10Hz -0.0037139 -0.0188953
+ 8.41e+10Hz -0.00374026 -0.0189057
+ 8.42e+10Hz -0.00376662 -0.018916
+ 8.43e+10Hz -0.003793 -0.0189263
+ 8.44e+10Hz -0.00381939 -0.0189366
+ 8.45e+10Hz -0.0038458 -0.0189468
+ 8.46e+10Hz -0.00387221 -0.018957
+ 8.47e+10Hz -0.00389864 -0.0189671
+ 8.48e+10Hz -0.00392508 -0.0189772
+ 8.49e+10Hz -0.00395154 -0.0189872
+ 8.5e+10Hz -0.00397801 -0.0189972
+ 8.51e+10Hz -0.00400449 -0.0190072
+ 8.52e+10Hz -0.00403099 -0.0190171
+ 8.53e+10Hz -0.00405749 -0.019027
+ 8.54e+10Hz -0.00408402 -0.0190368
+ 8.55e+10Hz -0.00411055 -0.0190466
+ 8.56e+10Hz -0.0041371 -0.0190563
+ 8.57e+10Hz -0.00416367 -0.019066
+ 8.58e+10Hz -0.00419024 -0.0190757
+ 8.59e+10Hz -0.00421683 -0.0190853
+ 8.6e+10Hz -0.00424344 -0.0190948
+ 8.61e+10Hz -0.00427006 -0.0191044
+ 8.62e+10Hz -0.00429669 -0.0191138
+ 8.63e+10Hz -0.00432333 -0.0191233
+ 8.64e+10Hz -0.00435 -0.0191327
+ 8.65e+10Hz -0.00437667 -0.019142
+ 8.66e+10Hz -0.00440336 -0.0191513
+ 8.67e+10Hz -0.00443006 -0.0191606
+ 8.68e+10Hz -0.00445678 -0.0191698
+ 8.69e+10Hz -0.00448351 -0.0191789
+ 8.7e+10Hz -0.00451025 -0.0191881
+ 8.71e+10Hz -0.00453701 -0.0191971
+ 8.72e+10Hz -0.00456379 -0.0192062
+ 8.73e+10Hz -0.00459057 -0.0192151
+ 8.74e+10Hz -0.00461738 -0.0192241
+ 8.75e+10Hz -0.00464419 -0.0192329
+ 8.76e+10Hz -0.00467102 -0.0192418
+ 8.77e+10Hz -0.00469786 -0.0192506
+ 8.78e+10Hz -0.00472472 -0.0192593
+ 8.79e+10Hz -0.00475159 -0.019268
+ 8.8e+10Hz -0.00477848 -0.0192766
+ 8.81e+10Hz -0.00480538 -0.0192852
+ 8.82e+10Hz -0.00483229 -0.0192938
+ 8.83e+10Hz -0.00485922 -0.0193023
+ 8.84e+10Hz -0.00488616 -0.0193107
+ 8.85e+10Hz -0.00491311 -0.0193191
+ 8.86e+10Hz -0.00494008 -0.0193275
+ 8.87e+10Hz -0.00496706 -0.0193358
+ 8.88e+10Hz -0.00499405 -0.019344
+ 8.89e+10Hz -0.00502106 -0.0193522
+ 8.9e+10Hz -0.00504808 -0.0193604
+ 8.91e+10Hz -0.00507512 -0.0193685
+ 8.92e+10Hz -0.00510216 -0.0193765
+ 8.93e+10Hz -0.00512922 -0.0193845
+ 8.94e+10Hz -0.00515629 -0.0193925
+ 8.95e+10Hz -0.00518338 -0.0194004
+ 8.96e+10Hz -0.00521047 -0.0194082
+ 8.97e+10Hz -0.00523758 -0.019416
+ 8.98e+10Hz -0.0052647 -0.0194237
+ 8.99e+10Hz -0.00529184 -0.0194314
+ 9e+10Hz -0.00531898 -0.019439
+ 9.01e+10Hz -0.00534614 -0.0194466
+ 9.02e+10Hz -0.0053733 -0.0194541
+ 9.03e+10Hz -0.00540048 -0.0194616
+ 9.04e+10Hz -0.00542767 -0.019469
+ 9.05e+10Hz -0.00545487 -0.0194764
+ 9.06e+10Hz -0.00548208 -0.0194837
+ 9.07e+10Hz -0.00550931 -0.0194909
+ 9.08e+10Hz -0.00553654 -0.0194981
+ 9.09e+10Hz -0.00556378 -0.0195053
+ 9.1e+10Hz -0.00559103 -0.0195124
+ 9.11e+10Hz -0.00561829 -0.0195194
+ 9.12e+10Hz -0.00564557 -0.0195264
+ 9.13e+10Hz -0.00567285 -0.0195333
+ 9.14e+10Hz -0.00570014 -0.0195402
+ 9.15e+10Hz -0.00572743 -0.019547
+ 9.16e+10Hz -0.00575474 -0.0195537
+ 9.17e+10Hz -0.00578206 -0.0195604
+ 9.18e+10Hz -0.00580938 -0.0195671
+ 9.19e+10Hz -0.00583671 -0.0195737
+ 9.2e+10Hz -0.00586405 -0.0195802
+ 9.21e+10Hz -0.0058914 -0.0195867
+ 9.22e+10Hz -0.00591875 -0.0195931
+ 9.23e+10Hz -0.00594611 -0.0195994
+ 9.24e+10Hz -0.00597347 -0.0196057
+ 9.25e+10Hz -0.00600085 -0.019612
+ 9.26e+10Hz -0.00602823 -0.0196182
+ 9.27e+10Hz -0.00605561 -0.0196243
+ 9.28e+10Hz -0.006083 -0.0196304
+ 9.29e+10Hz -0.00611039 -0.0196364
+ 9.3e+10Hz -0.00613779 -0.0196423
+ 9.31e+10Hz -0.0061652 -0.0196482
+ 9.32e+10Hz -0.00619261 -0.019654
+ 9.33e+10Hz -0.00622002 -0.0196598
+ 9.34e+10Hz -0.00624744 -0.0196655
+ 9.35e+10Hz -0.00627485 -0.0196712
+ 9.36e+10Hz -0.00630228 -0.0196768
+ 9.37e+10Hz -0.0063297 -0.0196823
+ 9.38e+10Hz -0.00635713 -0.0196878
+ 9.39e+10Hz -0.00638456 -0.0196932
+ 9.4e+10Hz -0.00641199 -0.0196986
+ 9.41e+10Hz -0.00643943 -0.0197039
+ 9.42e+10Hz -0.00646686 -0.0197091
+ 9.43e+10Hz -0.0064943 -0.0197143
+ 9.44e+10Hz -0.00652173 -0.0197194
+ 9.45e+10Hz -0.00654917 -0.0197245
+ 9.46e+10Hz -0.0065766 -0.0197295
+ 9.47e+10Hz -0.00660404 -0.0197344
+ 9.48e+10Hz -0.00663148 -0.0197393
+ 9.49e+10Hz -0.00665891 -0.0197441
+ 9.5e+10Hz -0.00668634 -0.0197489
+ 9.51e+10Hz -0.00671377 -0.0197536
+ 9.52e+10Hz -0.0067412 -0.0197582
+ 9.53e+10Hz -0.00676863 -0.0197628
+ 9.54e+10Hz -0.00679605 -0.0197673
+ 9.55e+10Hz -0.00682347 -0.0197718
+ 9.56e+10Hz -0.00685089 -0.0197762
+ 9.57e+10Hz -0.00687831 -0.0197805
+ 9.58e+10Hz -0.00690572 -0.0197848
+ 9.59e+10Hz -0.00693312 -0.019789
+ 9.6e+10Hz -0.00696052 -0.0197932
+ 9.61e+10Hz -0.00698792 -0.0197973
+ 9.62e+10Hz -0.00701531 -0.0198014
+ 9.63e+10Hz -0.0070427 -0.0198053
+ 9.64e+10Hz -0.00707008 -0.0198093
+ 9.65e+10Hz -0.00709745 -0.0198131
+ 9.66e+10Hz -0.00712482 -0.0198169
+ 9.67e+10Hz -0.00715218 -0.0198207
+ 9.68e+10Hz -0.00717953 -0.0198243
+ 9.69e+10Hz -0.00720688 -0.019828
+ 9.7e+10Hz -0.00723421 -0.0198315
+ 9.71e+10Hz -0.00726154 -0.019835
+ 9.72e+10Hz -0.00728887 -0.0198385
+ 9.73e+10Hz -0.00731618 -0.0198418
+ 9.74e+10Hz -0.00734348 -0.0198452
+ 9.75e+10Hz -0.00737078 -0.0198484
+ 9.76e+10Hz -0.00739806 -0.0198516
+ 9.77e+10Hz -0.00742533 -0.0198548
+ 9.78e+10Hz -0.0074526 -0.0198579
+ 9.79e+10Hz -0.00747985 -0.0198609
+ 9.8e+10Hz -0.0075071 -0.0198639
+ 9.81e+10Hz -0.00753433 -0.0198668
+ 9.82e+10Hz -0.00756155 -0.0198696
+ 9.83e+10Hz -0.00758876 -0.0198724
+ 9.84e+10Hz -0.00761595 -0.0198752
+ 9.85e+10Hz -0.00764314 -0.0198778
+ 9.86e+10Hz -0.00767031 -0.0198805
+ 9.87e+10Hz -0.00769747 -0.019883
+ 9.88e+10Hz -0.00772461 -0.0198855
+ 9.89e+10Hz -0.00775175 -0.019888
+ 9.9e+10Hz -0.00777887 -0.0198904
+ 9.91e+10Hz -0.00780597 -0.0198927
+ 9.92e+10Hz -0.00783306 -0.019895
+ 9.93e+10Hz -0.00786014 -0.0198972
+ 9.94e+10Hz -0.0078872 -0.0198993
+ 9.95e+10Hz -0.00791425 -0.0199014
+ 9.96e+10Hz -0.00794128 -0.0199035
+ 9.97e+10Hz -0.00796829 -0.0199055
+ 9.98e+10Hz -0.0079953 -0.0199074
+ 9.99e+10Hz -0.00802228 -0.0199093
+ 1e+11Hz -0.00804925 -0.0199111
+ 1.001e+11Hz -0.0080762 -0.0199129
+ 1.002e+11Hz -0.00810314 -0.0199146
+ 1.003e+11Hz -0.00813006 -0.0199162
+ 1.004e+11Hz -0.00815696 -0.0199178
+ 1.005e+11Hz -0.00818384 -0.0199194
+ 1.006e+11Hz -0.00821071 -0.0199209
+ 1.007e+11Hz -0.00823756 -0.0199223
+ 1.008e+11Hz -0.00826439 -0.0199237
+ 1.009e+11Hz -0.00829121 -0.019925
+ 1.01e+11Hz -0.008318 -0.0199263
+ 1.011e+11Hz -0.00834478 -0.0199275
+ 1.012e+11Hz -0.00837154 -0.0199287
+ 1.013e+11Hz -0.00839828 -0.0199298
+ 1.014e+11Hz -0.008425 -0.0199309
+ 1.015e+11Hz -0.0084517 -0.0199319
+ 1.016e+11Hz -0.00847838 -0.0199328
+ 1.017e+11Hz -0.00850504 -0.0199337
+ 1.018e+11Hz -0.00853169 -0.0199346
+ 1.019e+11Hz -0.00855831 -0.0199354
+ 1.02e+11Hz -0.00858491 -0.0199361
+ 1.021e+11Hz -0.0086115 -0.0199368
+ 1.022e+11Hz -0.00863806 -0.0199374
+ 1.023e+11Hz -0.0086646 -0.019938
+ 1.024e+11Hz -0.00869113 -0.0199386
+ 1.025e+11Hz -0.00871763 -0.019939
+ 1.026e+11Hz -0.00874411 -0.0199395
+ 1.027e+11Hz -0.00877057 -0.0199399
+ 1.028e+11Hz -0.00879701 -0.0199402
+ 1.029e+11Hz -0.00882343 -0.0199405
+ 1.03e+11Hz -0.00884982 -0.0199407
+ 1.031e+11Hz -0.0088762 -0.0199409
+ 1.032e+11Hz -0.00890255 -0.019941
+ 1.033e+11Hz -0.00892888 -0.0199411
+ 1.034e+11Hz -0.00895519 -0.0199412
+ 1.035e+11Hz -0.00898148 -0.0199412
+ 1.036e+11Hz -0.00900775 -0.0199411
+ 1.037e+11Hz -0.00903399 -0.019941
+ 1.038e+11Hz -0.00906022 -0.0199408
+ 1.039e+11Hz -0.00908642 -0.0199406
+ 1.04e+11Hz -0.0091126 -0.0199404
+ 1.041e+11Hz -0.00913875 -0.0199401
+ 1.042e+11Hz -0.00916489 -0.0199397
+ 1.043e+11Hz -0.009191 -0.0199393
+ 1.044e+11Hz -0.00921709 -0.0199389
+ 1.045e+11Hz -0.00924315 -0.0199384
+ 1.046e+11Hz -0.0092692 -0.0199378
+ 1.047e+11Hz -0.00929522 -0.0199373
+ 1.048e+11Hz -0.00932122 -0.0199366
+ 1.049e+11Hz -0.00934719 -0.0199359
+ 1.05e+11Hz -0.00937315 -0.0199352
+ 1.051e+11Hz -0.00939908 -0.0199345
+ 1.052e+11Hz -0.00942498 -0.0199336
+ 1.053e+11Hz -0.00945087 -0.0199328
+ 1.054e+11Hz -0.00947673 -0.0199319
+ 1.055e+11Hz -0.00950257 -0.0199309
+ 1.056e+11Hz -0.00952838 -0.0199299
+ 1.057e+11Hz -0.00955417 -0.0199289
+ 1.058e+11Hz -0.00957994 -0.0199278
+ 1.059e+11Hz -0.00960569 -0.0199267
+ 1.06e+11Hz -0.00963141 -0.0199255
+ 1.061e+11Hz -0.00965711 -0.0199243
+ 1.062e+11Hz -0.00968279 -0.019923
+ 1.063e+11Hz -0.00970844 -0.0199217
+ 1.064e+11Hz -0.00973407 -0.0199203
+ 1.065e+11Hz -0.00975968 -0.0199189
+ 1.066e+11Hz -0.00978526 -0.0199175
+ 1.067e+11Hz -0.00981082 -0.019916
+ 1.068e+11Hz -0.00983636 -0.0199145
+ 1.069e+11Hz -0.00986187 -0.0199129
+ 1.07e+11Hz -0.00988736 -0.0199113
+ 1.071e+11Hz -0.00991283 -0.0199096
+ 1.072e+11Hz -0.00993828 -0.019908
+ 1.073e+11Hz -0.0099637 -0.0199062
+ 1.074e+11Hz -0.00998909 -0.0199044
+ 1.075e+11Hz -0.0100145 -0.0199026
+ 1.076e+11Hz -0.0100398 -0.0199007
+ 1.077e+11Hz -0.0100651 -0.0198988
+ 1.078e+11Hz -0.0100905 -0.0198969
+ 1.079e+11Hz -0.0101157 -0.0198949
+ 1.08e+11Hz -0.010141 -0.0198928
+ 1.081e+11Hz -0.0101662 -0.0198908
+ 1.082e+11Hz -0.0101914 -0.0198886
+ 1.083e+11Hz -0.0102166 -0.0198865
+ 1.084e+11Hz -0.0102418 -0.0198843
+ 1.085e+11Hz -0.0102669 -0.019882
+ 1.086e+11Hz -0.0102921 -0.0198797
+ 1.087e+11Hz -0.0103172 -0.0198774
+ 1.088e+11Hz -0.0103422 -0.019875
+ 1.089e+11Hz -0.0103673 -0.0198726
+ 1.09e+11Hz -0.0103923 -0.0198702
+ 1.091e+11Hz -0.0104173 -0.0198677
+ 1.092e+11Hz -0.0104423 -0.0198652
+ 1.093e+11Hz -0.0104672 -0.0198626
+ 1.094e+11Hz -0.0104922 -0.01986
+ 1.095e+11Hz -0.0105171 -0.0198573
+ 1.096e+11Hz -0.010542 -0.0198546
+ 1.097e+11Hz -0.0105668 -0.0198519
+ 1.098e+11Hz -0.0105917 -0.0198491
+ 1.099e+11Hz -0.0106165 -0.0198463
+ 1.1e+11Hz -0.0106413 -0.0198434
+ 1.101e+11Hz -0.0106661 -0.0198405
+ 1.102e+11Hz -0.0106908 -0.0198376
+ 1.103e+11Hz -0.0107155 -0.0198346
+ 1.104e+11Hz -0.0107403 -0.0198316
+ 1.105e+11Hz -0.0107649 -0.0198285
+ 1.106e+11Hz -0.0107896 -0.0198254
+ 1.107e+11Hz -0.0108142 -0.0198223
+ 1.108e+11Hz -0.0108388 -0.0198191
+ 1.109e+11Hz -0.0108634 -0.0198159
+ 1.11e+11Hz -0.010888 -0.0198126
+ 1.111e+11Hz -0.0109125 -0.0198093
+ 1.112e+11Hz -0.010937 -0.019806
+ 1.113e+11Hz -0.0109615 -0.0198026
+ 1.114e+11Hz -0.010986 -0.0197992
+ 1.115e+11Hz -0.0110105 -0.0197957
+ 1.116e+11Hz -0.0110349 -0.0197922
+ 1.117e+11Hz -0.0110593 -0.0197887
+ 1.118e+11Hz -0.0110837 -0.0197851
+ 1.119e+11Hz -0.011108 -0.0197815
+ 1.12e+11Hz -0.0111324 -0.0197778
+ 1.121e+11Hz -0.0111567 -0.0197741
+ 1.122e+11Hz -0.011181 -0.0197704
+ 1.123e+11Hz -0.0112052 -0.0197666
+ 1.124e+11Hz -0.0112295 -0.0197628
+ 1.125e+11Hz -0.0112537 -0.0197589
+ 1.126e+11Hz -0.0112779 -0.019755
+ 1.127e+11Hz -0.011302 -0.0197511
+ 1.128e+11Hz -0.0113262 -0.0197471
+ 1.129e+11Hz -0.0113503 -0.0197431
+ 1.13e+11Hz -0.0113744 -0.019739
+ 1.131e+11Hz -0.0113985 -0.0197349
+ 1.132e+11Hz -0.0114225 -0.0197308
+ 1.133e+11Hz -0.0114466 -0.0197266
+ 1.134e+11Hz -0.0114706 -0.0197224
+ 1.135e+11Hz -0.0114945 -0.0197181
+ 1.136e+11Hz -0.0115185 -0.0197138
+ 1.137e+11Hz -0.0115424 -0.0197095
+ 1.138e+11Hz -0.0115663 -0.0197051
+ 1.139e+11Hz -0.0115902 -0.0197007
+ 1.14e+11Hz -0.0116141 -0.0196962
+ 1.141e+11Hz -0.0116379 -0.0196917
+ 1.142e+11Hz -0.0116617 -0.0196872
+ 1.143e+11Hz -0.0116855 -0.0196826
+ 1.144e+11Hz -0.0117093 -0.019678
+ 1.145e+11Hz -0.011733 -0.0196733
+ 1.146e+11Hz -0.0117567 -0.0196686
+ 1.147e+11Hz -0.0117804 -0.0196638
+ 1.148e+11Hz -0.0118041 -0.0196591
+ 1.149e+11Hz -0.0118277 -0.0196542
+ 1.15e+11Hz -0.0118513 -0.0196494
+ 1.151e+11Hz -0.0118749 -0.0196445
+ 1.152e+11Hz -0.0118985 -0.0196395
+ 1.153e+11Hz -0.011922 -0.0196345
+ 1.154e+11Hz -0.0119455 -0.0196295
+ 1.155e+11Hz -0.011969 -0.0196245
+ 1.156e+11Hz -0.0119925 -0.0196194
+ 1.157e+11Hz -0.0120159 -0.0196142
+ 1.158e+11Hz -0.0120393 -0.019609
+ 1.159e+11Hz -0.0120627 -0.0196038
+ 1.16e+11Hz -0.012086 -0.0195985
+ 1.161e+11Hz -0.0121094 -0.0195932
+ 1.162e+11Hz -0.0121327 -0.0195879
+ 1.163e+11Hz -0.0121559 -0.0195825
+ 1.164e+11Hz -0.0121792 -0.019577
+ 1.165e+11Hz -0.0122024 -0.0195716
+ 1.166e+11Hz -0.0122256 -0.0195661
+ 1.167e+11Hz -0.0122488 -0.0195605
+ 1.168e+11Hz -0.0122719 -0.0195549
+ 1.169e+11Hz -0.012295 -0.0195493
+ 1.17e+11Hz -0.0123181 -0.0195436
+ 1.171e+11Hz -0.0123412 -0.0195379
+ 1.172e+11Hz -0.0123642 -0.0195322
+ 1.173e+11Hz -0.0123872 -0.0195264
+ 1.174e+11Hz -0.0124102 -0.0195205
+ 1.175e+11Hz -0.0124331 -0.0195147
+ 1.176e+11Hz -0.012456 -0.0195087
+ 1.177e+11Hz -0.0124789 -0.0195028
+ 1.178e+11Hz -0.0125018 -0.0194968
+ 1.179e+11Hz -0.0125246 -0.0194908
+ 1.18e+11Hz -0.0125474 -0.0194847
+ 1.181e+11Hz -0.0125702 -0.0194786
+ 1.182e+11Hz -0.0125929 -0.0194724
+ 1.183e+11Hz -0.0126157 -0.0194662
+ 1.184e+11Hz -0.0126383 -0.01946
+ 1.185e+11Hz -0.012661 -0.0194537
+ 1.186e+11Hz -0.0126836 -0.0194474
+ 1.187e+11Hz -0.0127062 -0.019441
+ 1.188e+11Hz -0.0127288 -0.0194346
+ 1.189e+11Hz -0.0127513 -0.0194282
+ 1.19e+11Hz -0.0127738 -0.0194217
+ 1.191e+11Hz -0.0127963 -0.0194152
+ 1.192e+11Hz -0.0128187 -0.0194086
+ 1.193e+11Hz -0.0128411 -0.019402
+ 1.194e+11Hz -0.0128635 -0.0193954
+ 1.195e+11Hz -0.0128859 -0.0193887
+ 1.196e+11Hz -0.0129082 -0.019382
+ 1.197e+11Hz -0.0129304 -0.0193752
+ 1.198e+11Hz -0.0129527 -0.0193684
+ 1.199e+11Hz -0.0129749 -0.0193616
+ 1.2e+11Hz -0.0129971 -0.0193547
+ 1.201e+11Hz -0.0130192 -0.0193478
+ 1.202e+11Hz -0.0130414 -0.0193409
+ 1.203e+11Hz -0.0130635 -0.0193339
+ 1.204e+11Hz -0.0130855 -0.0193268
+ 1.205e+11Hz -0.0131075 -0.0193198
+ 1.206e+11Hz -0.0131295 -0.0193126
+ 1.207e+11Hz -0.0131515 -0.0193055
+ 1.208e+11Hz -0.0131734 -0.0192983
+ 1.209e+11Hz -0.0131953 -0.0192911
+ 1.21e+11Hz -0.0132171 -0.0192838
+ 1.211e+11Hz -0.0132389 -0.0192765
+ 1.212e+11Hz -0.0132607 -0.0192692
+ 1.213e+11Hz -0.0132824 -0.0192618
+ 1.214e+11Hz -0.0133041 -0.0192544
+ 1.215e+11Hz -0.0133258 -0.0192469
+ 1.216e+11Hz -0.0133475 -0.0192394
+ 1.217e+11Hz -0.0133691 -0.0192319
+ 1.218e+11Hz -0.0133906 -0.0192243
+ 1.219e+11Hz -0.0134122 -0.0192167
+ 1.22e+11Hz -0.0134336 -0.019209
+ 1.221e+11Hz -0.0134551 -0.0192013
+ 1.222e+11Hz -0.0134765 -0.0191936
+ 1.223e+11Hz -0.0134979 -0.0191859
+ 1.224e+11Hz -0.0135192 -0.0191781
+ 1.225e+11Hz -0.0135405 -0.0191702
+ 1.226e+11Hz -0.0135618 -0.0191624
+ 1.227e+11Hz -0.013583 -0.0191544
+ 1.228e+11Hz -0.0136042 -0.0191465
+ 1.229e+11Hz -0.0136254 -0.0191385
+ 1.23e+11Hz -0.0136465 -0.0191305
+ 1.231e+11Hz -0.0136676 -0.0191225
+ 1.232e+11Hz -0.0136886 -0.0191144
+ 1.233e+11Hz -0.0137096 -0.0191062
+ 1.234e+11Hz -0.0137306 -0.0190981
+ 1.235e+11Hz -0.0137515 -0.0190899
+ 1.236e+11Hz -0.0137724 -0.0190816
+ 1.237e+11Hz -0.0137932 -0.0190734
+ 1.238e+11Hz -0.013814 -0.0190651
+ 1.239e+11Hz -0.0138348 -0.0190567
+ 1.24e+11Hz -0.0138555 -0.0190484
+ 1.241e+11Hz -0.0138762 -0.01904
+ 1.242e+11Hz -0.0138969 -0.0190315
+ 1.243e+11Hz -0.0139175 -0.019023
+ 1.244e+11Hz -0.013938 -0.0190145
+ 1.245e+11Hz -0.0139585 -0.019006
+ 1.246e+11Hz -0.013979 -0.0189974
+ 1.247e+11Hz -0.0139995 -0.0189888
+ 1.248e+11Hz -0.0140199 -0.0189802
+ 1.249e+11Hz -0.0140402 -0.0189715
+ 1.25e+11Hz -0.0140605 -0.0189628
+ 1.251e+11Hz -0.0140808 -0.018954
+ 1.252e+11Hz -0.014101 -0.0189452
+ 1.253e+11Hz -0.0141212 -0.0189364
+ 1.254e+11Hz -0.0141414 -0.0189276
+ 1.255e+11Hz -0.0141615 -0.0189187
+ 1.256e+11Hz -0.0141815 -0.0189098
+ 1.257e+11Hz -0.0142015 -0.0189009
+ 1.258e+11Hz -0.0142215 -0.0188919
+ 1.259e+11Hz -0.0142414 -0.0188829
+ 1.26e+11Hz -0.0142613 -0.0188739
+ 1.261e+11Hz -0.0142812 -0.0188648
+ 1.262e+11Hz -0.014301 -0.0188557
+ 1.263e+11Hz -0.0143207 -0.0188466
+ 1.264e+11Hz -0.0143404 -0.0188375
+ 1.265e+11Hz -0.0143601 -0.0188283
+ 1.266e+11Hz -0.0143797 -0.0188191
+ 1.267e+11Hz -0.0143993 -0.0188098
+ 1.268e+11Hz -0.0144188 -0.0188006
+ 1.269e+11Hz -0.0144383 -0.0187913
+ 1.27e+11Hz -0.0144578 -0.018782
+ 1.271e+11Hz -0.0144772 -0.0187726
+ 1.272e+11Hz -0.0144965 -0.0187632
+ 1.273e+11Hz -0.0145159 -0.0187538
+ 1.274e+11Hz -0.0145351 -0.0187444
+ 1.275e+11Hz -0.0145543 -0.0187349
+ 1.276e+11Hz -0.0145735 -0.0187254
+ 1.277e+11Hz -0.0145926 -0.0187159
+ 1.278e+11Hz -0.0146117 -0.0187063
+ 1.279e+11Hz -0.0146308 -0.0186968
+ 1.28e+11Hz -0.0146498 -0.0186872
+ 1.281e+11Hz -0.0146687 -0.0186775
+ 1.282e+11Hz -0.0146876 -0.0186679
+ 1.283e+11Hz -0.0147065 -0.0186582
+ 1.284e+11Hz -0.0147253 -0.0186485
+ 1.285e+11Hz -0.0147441 -0.0186388
+ 1.286e+11Hz -0.0147628 -0.018629
+ 1.287e+11Hz -0.0147814 -0.0186192
+ 1.288e+11Hz -0.0148001 -0.0186094
+ 1.289e+11Hz -0.0148186 -0.0185996
+ 1.29e+11Hz -0.0148372 -0.0185897
+ 1.291e+11Hz -0.0148557 -0.0185799
+ 1.292e+11Hz -0.0148741 -0.01857
+ 1.293e+11Hz -0.0148925 -0.01856
+ 1.294e+11Hz -0.0149108 -0.0185501
+ 1.295e+11Hz -0.0149291 -0.0185401
+ 1.296e+11Hz -0.0149474 -0.0185301
+ 1.297e+11Hz -0.0149656 -0.0185201
+ 1.298e+11Hz -0.0149838 -0.0185101
+ 1.299e+11Hz -0.0150019 -0.0185
+ 1.3e+11Hz -0.0150199 -0.0184899
+ 1.301e+11Hz -0.0150379 -0.0184798
+ 1.302e+11Hz -0.0150559 -0.0184697
+ 1.303e+11Hz -0.0150738 -0.0184595
+ 1.304e+11Hz -0.0150917 -0.0184494
+ 1.305e+11Hz -0.0151095 -0.0184392
+ 1.306e+11Hz -0.0151273 -0.018429
+ 1.307e+11Hz -0.015145 -0.0184187
+ 1.308e+11Hz -0.0151627 -0.0184085
+ 1.309e+11Hz -0.0151804 -0.0183982
+ 1.31e+11Hz -0.0151979 -0.0183879
+ 1.311e+11Hz -0.0152155 -0.0183776
+ 1.312e+11Hz -0.015233 -0.0183673
+ 1.313e+11Hz -0.0152504 -0.018357
+ 1.314e+11Hz -0.0152678 -0.0183466
+ 1.315e+11Hz -0.0152852 -0.0183362
+ 1.316e+11Hz -0.0153025 -0.0183258
+ 1.317e+11Hz -0.0153197 -0.0183154
+ 1.318e+11Hz -0.0153369 -0.018305
+ 1.319e+11Hz -0.0153541 -0.0182945
+ 1.32e+11Hz -0.0153712 -0.018284
+ 1.321e+11Hz -0.0153883 -0.0182735
+ 1.322e+11Hz -0.0154053 -0.018263
+ 1.323e+11Hz -0.0154222 -0.0182525
+ 1.324e+11Hz -0.0154392 -0.018242
+ 1.325e+11Hz -0.015456 -0.0182314
+ 1.326e+11Hz -0.0154729 -0.0182209
+ 1.327e+11Hz -0.0154896 -0.0182103
+ 1.328e+11Hz -0.0155064 -0.0181997
+ 1.329e+11Hz -0.015523 -0.0181891
+ 1.33e+11Hz -0.0155397 -0.0181784
+ 1.331e+11Hz -0.0155562 -0.0181678
+ 1.332e+11Hz -0.0155728 -0.0181571
+ 1.333e+11Hz -0.0155893 -0.0181464
+ 1.334e+11Hz -0.0156057 -0.0181358
+ 1.335e+11Hz -0.0156221 -0.0181251
+ 1.336e+11Hz -0.0156384 -0.0181143
+ 1.337e+11Hz -0.0156547 -0.0181036
+ 1.338e+11Hz -0.015671 -0.0180929
+ 1.339e+11Hz -0.0156872 -0.0180821
+ 1.34e+11Hz -0.0157033 -0.0180714
+ 1.341e+11Hz -0.0157194 -0.0180606
+ 1.342e+11Hz -0.0157355 -0.0180498
+ 1.343e+11Hz -0.0157515 -0.018039
+ 1.344e+11Hz -0.0157674 -0.0180282
+ 1.345e+11Hz -0.0157833 -0.0180173
+ 1.346e+11Hz -0.0157992 -0.0180065
+ 1.347e+11Hz -0.015815 -0.0179956
+ 1.348e+11Hz -0.0158308 -0.0179848
+ 1.349e+11Hz -0.0158465 -0.0179739
+ 1.35e+11Hz -0.0158622 -0.017963
+ 1.351e+11Hz -0.0158778 -0.0179521
+ 1.352e+11Hz -0.0158933 -0.0179412
+ 1.353e+11Hz -0.0159089 -0.0179303
+ 1.354e+11Hz -0.0159243 -0.0179194
+ 1.355e+11Hz -0.0159398 -0.0179084
+ 1.356e+11Hz -0.0159552 -0.0178975
+ 1.357e+11Hz -0.0159705 -0.0178865
+ 1.358e+11Hz -0.0159858 -0.0178756
+ 1.359e+11Hz -0.016001 -0.0178646
+ 1.36e+11Hz -0.0160162 -0.0178536
+ 1.361e+11Hz -0.0160313 -0.0178426
+ 1.362e+11Hz -0.0160464 -0.0178316
+ 1.363e+11Hz -0.0160615 -0.0178206
+ 1.364e+11Hz -0.0160765 -0.0178096
+ 1.365e+11Hz -0.0160914 -0.0177986
+ 1.366e+11Hz -0.0161063 -0.0177876
+ 1.367e+11Hz -0.0161212 -0.0177765
+ 1.368e+11Hz -0.016136 -0.0177655
+ 1.369e+11Hz -0.0161507 -0.0177544
+ 1.37e+11Hz -0.0161654 -0.0177434
+ 1.371e+11Hz -0.0161801 -0.0177323
+ 1.372e+11Hz -0.0161947 -0.0177212
+ 1.373e+11Hz -0.0162093 -0.0177101
+ 1.374e+11Hz -0.0162238 -0.0176991
+ 1.375e+11Hz -0.0162383 -0.017688
+ 1.376e+11Hz -0.0162527 -0.0176769
+ 1.377e+11Hz -0.0162671 -0.0176658
+ 1.378e+11Hz -0.0162814 -0.0176547
+ 1.379e+11Hz -0.0162957 -0.0176436
+ 1.38e+11Hz -0.0163099 -0.0176324
+ 1.381e+11Hz -0.0163241 -0.0176213
+ 1.382e+11Hz -0.0163382 -0.0176102
+ 1.383e+11Hz -0.0163523 -0.0175991
+ 1.384e+11Hz -0.0163663 -0.0175879
+ 1.385e+11Hz -0.0163803 -0.0175768
+ 1.386e+11Hz -0.0163943 -0.0175656
+ 1.387e+11Hz -0.0164082 -0.0175545
+ 1.388e+11Hz -0.016422 -0.0175433
+ 1.389e+11Hz -0.0164358 -0.0175322
+ 1.39e+11Hz -0.0164495 -0.017521
+ 1.391e+11Hz -0.0164633 -0.0175099
+ 1.392e+11Hz -0.0164769 -0.0174987
+ 1.393e+11Hz -0.0164905 -0.0174875
+ 1.394e+11Hz -0.0165041 -0.0174764
+ 1.395e+11Hz -0.0165176 -0.0174652
+ 1.396e+11Hz -0.016531 -0.017454
+ 1.397e+11Hz -0.0165445 -0.0174429
+ 1.398e+11Hz -0.0165578 -0.0174317
+ 1.399e+11Hz -0.0165711 -0.0174205
+ 1.4e+11Hz -0.0165844 -0.0174093
+ 1.401e+11Hz -0.0165976 -0.0173981
+ 1.402e+11Hz -0.0166108 -0.017387
+ 1.403e+11Hz -0.0166239 -0.0173758
+ 1.404e+11Hz -0.016637 -0.0173646
+ 1.405e+11Hz -0.0166501 -0.0173534
+ 1.406e+11Hz -0.016663 -0.0173422
+ 1.407e+11Hz -0.016676 -0.017331
+ 1.408e+11Hz -0.0166889 -0.0173199
+ 1.409e+11Hz -0.0167017 -0.0173087
+ 1.41e+11Hz -0.0167145 -0.0172975
+ 1.411e+11Hz -0.0167272 -0.0172863
+ 1.412e+11Hz -0.0167399 -0.0172751
+ 1.413e+11Hz -0.0167526 -0.017264
+ 1.414e+11Hz -0.0167652 -0.0172528
+ 1.415e+11Hz -0.0167777 -0.0172416
+ 1.416e+11Hz -0.0167902 -0.0172304
+ 1.417e+11Hz -0.0168027 -0.0172193
+ 1.418e+11Hz -0.0168151 -0.0172081
+ 1.419e+11Hz -0.0168274 -0.0171969
+ 1.42e+11Hz -0.0168398 -0.0171858
+ 1.421e+11Hz -0.016852 -0.0171746
+ 1.422e+11Hz -0.0168642 -0.0171634
+ 1.423e+11Hz -0.0168764 -0.0171523
+ 1.424e+11Hz -0.0168885 -0.0171411
+ 1.425e+11Hz -0.0169006 -0.01713
+ 1.426e+11Hz -0.0169126 -0.0171189
+ 1.427e+11Hz -0.0169246 -0.0171077
+ 1.428e+11Hz -0.0169365 -0.0170966
+ 1.429e+11Hz -0.0169484 -0.0170855
+ 1.43e+11Hz -0.0169602 -0.0170743
+ 1.431e+11Hz -0.016972 -0.0170632
+ 1.432e+11Hz -0.0169837 -0.0170521
+ 1.433e+11Hz -0.0169954 -0.017041
+ 1.434e+11Hz -0.017007 -0.0170299
+ 1.435e+11Hz -0.0170186 -0.0170188
+ 1.436e+11Hz -0.0170301 -0.0170077
+ 1.437e+11Hz -0.0170416 -0.0169966
+ 1.438e+11Hz -0.017053 -0.0169856
+ 1.439e+11Hz -0.0170644 -0.0169745
+ 1.44e+11Hz -0.0170757 -0.0169634
+ 1.441e+11Hz -0.017087 -0.0169524
+ 1.442e+11Hz -0.0170983 -0.0169413
+ 1.443e+11Hz -0.0171094 -0.0169303
+ 1.444e+11Hz -0.0171206 -0.0169193
+ 1.445e+11Hz -0.0171317 -0.0169083
+ 1.446e+11Hz -0.0171427 -0.0168973
+ 1.447e+11Hz -0.0171537 -0.0168863
+ 1.448e+11Hz -0.0171646 -0.0168753
+ 1.449e+11Hz -0.0171755 -0.0168643
+ 1.45e+11Hz -0.0171864 -0.0168533
+ 1.451e+11Hz -0.0171972 -0.0168424
+ 1.452e+11Hz -0.0172079 -0.0168314
+ 1.453e+11Hz -0.0172186 -0.0168205
+ 1.454e+11Hz -0.0172293 -0.0168096
+ 1.455e+11Hz -0.0172399 -0.0167987
+ 1.456e+11Hz -0.0172504 -0.0167878
+ 1.457e+11Hz -0.0172609 -0.0167769
+ 1.458e+11Hz -0.0172714 -0.016766
+ 1.459e+11Hz -0.0172818 -0.0167551
+ 1.46e+11Hz -0.0172921 -0.0167443
+ 1.461e+11Hz -0.0173024 -0.0167335
+ 1.462e+11Hz -0.0173127 -0.0167227
+ 1.463e+11Hz -0.0173229 -0.0167119
+ 1.464e+11Hz -0.017333 -0.0167011
+ 1.465e+11Hz -0.0173432 -0.0166903
+ 1.466e+11Hz -0.0173532 -0.0166795
+ 1.467e+11Hz -0.0173632 -0.0166688
+ 1.468e+11Hz -0.0173732 -0.0166581
+ 1.469e+11Hz -0.0173831 -0.0166474
+ 1.47e+11Hz -0.017393 -0.0166367
+ 1.471e+11Hz -0.0174028 -0.016626
+ 1.472e+11Hz -0.0174125 -0.0166154
+ 1.473e+11Hz -0.0174222 -0.0166047
+ 1.474e+11Hz -0.0174319 -0.0165941
+ 1.475e+11Hz -0.0174415 -0.0165835
+ 1.476e+11Hz -0.0174511 -0.0165729
+ 1.477e+11Hz -0.0174606 -0.0165624
+ 1.478e+11Hz -0.0174701 -0.0165518
+ 1.479e+11Hz -0.0174795 -0.0165413
+ 1.48e+11Hz -0.0174889 -0.0165308
+ 1.481e+11Hz -0.0174982 -0.0165203
+ 1.482e+11Hz -0.0175074 -0.0165099
+ 1.483e+11Hz -0.0175167 -0.0164994
+ 1.484e+11Hz -0.0175258 -0.016489
+ 1.485e+11Hz -0.017535 -0.0164787
+ 1.486e+11Hz -0.0175441 -0.0164683
+ 1.487e+11Hz -0.0175531 -0.0164579
+ 1.488e+11Hz -0.0175621 -0.0164476
+ 1.489e+11Hz -0.017571 -0.0164373
+ 1.49e+11Hz -0.0175799 -0.0164271
+ 1.491e+11Hz -0.0175887 -0.0164168
+ 1.492e+11Hz -0.0175975 -0.0164066
+ 1.493e+11Hz -0.0176063 -0.0163964
+ 1.494e+11Hz -0.0176149 -0.0163863
+ 1.495e+11Hz -0.0176236 -0.0163762
+ 1.496e+11Hz -0.0176322 -0.016366
+ 1.497e+11Hz -0.0176407 -0.016356
+ 1.498e+11Hz -0.0176492 -0.0163459
+ 1.499e+11Hz -0.0176577 -0.0163359
+ 1.5e+11Hz -0.0176661 -0.0163259
+ 1.501e+11Hz -0.0176745 -0.016316
+ 1.502e+11Hz -0.0176828 -0.016306
+ 1.503e+11Hz -0.0176911 -0.0162961
+ 1.504e+11Hz -0.0176993 -0.0162863
+ 1.505e+11Hz -0.0177075 -0.0162764
+ 1.506e+11Hz -0.0177156 -0.0162666
+ 1.507e+11Hz -0.0177237 -0.0162569
+ 1.508e+11Hz -0.0177317 -0.0162471
+ 1.509e+11Hz -0.0177397 -0.0162374
+ 1.51e+11Hz -0.0177477 -0.0162278
+ 1.511e+11Hz -0.0177556 -0.0162181
+ 1.512e+11Hz -0.0177634 -0.0162085
+ 1.513e+11Hz -0.0177713 -0.016199
+ 1.514e+11Hz -0.017779 -0.0161895
+ 1.515e+11Hz -0.0177868 -0.01618
+ 1.516e+11Hz -0.0177944 -0.0161705
+ 1.517e+11Hz -0.0178021 -0.0161611
+ 1.518e+11Hz -0.0178097 -0.0161518
+ 1.519e+11Hz -0.0178172 -0.0161424
+ 1.52e+11Hz -0.0178247 -0.0161331
+ 1.521e+11Hz -0.0178322 -0.0161239
+ 1.522e+11Hz -0.0178396 -0.0161147
+ 1.523e+11Hz -0.017847 -0.0161055
+ 1.524e+11Hz -0.0178544 -0.0160964
+ 1.525e+11Hz -0.0178617 -0.0160873
+ 1.526e+11Hz -0.0178689 -0.0160782
+ 1.527e+11Hz -0.0178762 -0.0160692
+ 1.528e+11Hz -0.0178833 -0.0160603
+ 1.529e+11Hz -0.0178905 -0.0160513
+ 1.53e+11Hz -0.0178976 -0.0160425
+ 1.531e+11Hz -0.0179046 -0.0160336
+ 1.532e+11Hz -0.0179117 -0.0160249
+ 1.533e+11Hz -0.0179187 -0.0160161
+ 1.534e+11Hz -0.0179256 -0.0160074
+ 1.535e+11Hz -0.0179325 -0.0159988
+ 1.536e+11Hz -0.0179394 -0.0159902
+ 1.537e+11Hz -0.0179462 -0.0159817
+ 1.538e+11Hz -0.017953 -0.0159732
+ 1.539e+11Hz -0.0179598 -0.0159647
+ 1.54e+11Hz -0.0179665 -0.0159563
+ 1.541e+11Hz -0.0179732 -0.015948
+ 1.542e+11Hz -0.0179799 -0.0159397
+ 1.543e+11Hz -0.0179865 -0.0159314
+ 1.544e+11Hz -0.0179931 -0.0159232
+ 1.545e+11Hz -0.0179996 -0.0159151
+ 1.546e+11Hz -0.0180062 -0.015907
+ 1.547e+11Hz -0.0180126 -0.0158989
+ 1.548e+11Hz -0.0180191 -0.0158909
+ 1.549e+11Hz -0.0180255 -0.015883
+ 1.55e+11Hz -0.0180319 -0.0158751
+ 1.551e+11Hz -0.0180383 -0.0158673
+ 1.552e+11Hz -0.0180446 -0.0158595
+ 1.553e+11Hz -0.0180509 -0.0158518
+ 1.554e+11Hz -0.0180572 -0.0158442
+ 1.555e+11Hz -0.0180635 -0.0158366
+ 1.556e+11Hz -0.0180697 -0.015829
+ 1.557e+11Hz -0.0180759 -0.0158215
+ 1.558e+11Hz -0.0180821 -0.0158141
+ 1.559e+11Hz -0.0180882 -0.0158067
+ 1.56e+11Hz -0.0180943 -0.0157994
+ 1.561e+11Hz -0.0181004 -0.0157922
+ 1.562e+11Hz -0.0181065 -0.015785
+ 1.563e+11Hz -0.0181126 -0.0157779
+ 1.564e+11Hz -0.0181186 -0.0157708
+ 1.565e+11Hz -0.0181246 -0.0157638
+ 1.566e+11Hz -0.0181306 -0.0157568
+ 1.567e+11Hz -0.0181365 -0.0157499
+ 1.568e+11Hz -0.0181425 -0.0157431
+ 1.569e+11Hz -0.0181484 -0.0157364
+ 1.57e+11Hz -0.0181543 -0.0157297
+ 1.571e+11Hz -0.0181602 -0.015723
+ 1.572e+11Hz -0.0181661 -0.0157164
+ 1.573e+11Hz -0.0181719 -0.0157099
+ 1.574e+11Hz -0.0181778 -0.0157035
+ 1.575e+11Hz -0.0181836 -0.0156971
+ 1.576e+11Hz -0.0181894 -0.0156908
+ 1.577e+11Hz -0.0181952 -0.0156845
+ 1.578e+11Hz -0.018201 -0.0156784
+ 1.579e+11Hz -0.0182068 -0.0156722
+ 1.58e+11Hz -0.0182125 -0.0156662
+ 1.581e+11Hz -0.0182183 -0.0156602
+ 1.582e+11Hz -0.018224 -0.0156543
+ 1.583e+11Hz -0.0182298 -0.0156484
+ 1.584e+11Hz -0.0182355 -0.0156427
+ 1.585e+11Hz -0.0182412 -0.0156369
+ 1.586e+11Hz -0.0182469 -0.0156313
+ 1.587e+11Hz -0.0182526 -0.0156257
+ 1.588e+11Hz -0.0182583 -0.0156202
+ 1.589e+11Hz -0.018264 -0.0156148
+ 1.59e+11Hz -0.0182697 -0.0156094
+ 1.591e+11Hz -0.0182754 -0.0156041
+ 1.592e+11Hz -0.0182811 -0.0155988
+ 1.593e+11Hz -0.0182868 -0.0155937
+ 1.594e+11Hz -0.0182925 -0.0155886
+ 1.595e+11Hz -0.0182982 -0.0155835
+ 1.596e+11Hz -0.0183039 -0.0155786
+ 1.597e+11Hz -0.0183096 -0.0155737
+ 1.598e+11Hz -0.0183153 -0.0155689
+ 1.599e+11Hz -0.018321 -0.0155641
+ 1.6e+11Hz -0.0183267 -0.0155595
+ 1.601e+11Hz -0.0183325 -0.0155549
+ 1.602e+11Hz -0.0183382 -0.0155503
+ 1.603e+11Hz -0.0183439 -0.0155459
+ 1.604e+11Hz -0.0183497 -0.0155415
+ 1.605e+11Hz -0.0183555 -0.0155371
+ 1.606e+11Hz -0.0183612 -0.0155329
+ 1.607e+11Hz -0.018367 -0.0155287
+ 1.608e+11Hz -0.0183728 -0.0155246
+ 1.609e+11Hz -0.0183786 -0.0155206
+ 1.61e+11Hz -0.0183845 -0.0155166
+ 1.611e+11Hz -0.0183903 -0.0155127
+ 1.612e+11Hz -0.0183962 -0.0155089
+ 1.613e+11Hz -0.0184021 -0.0155051
+ 1.614e+11Hz -0.018408 -0.0155014
+ 1.615e+11Hz -0.0184139 -0.0154978
+ 1.616e+11Hz -0.0184199 -0.0154943
+ 1.617e+11Hz -0.0184258 -0.0154908
+ 1.618e+11Hz -0.0184318 -0.0154874
+ 1.619e+11Hz -0.0184378 -0.0154841
+ 1.62e+11Hz -0.0184439 -0.0154808
+ 1.621e+11Hz -0.0184499 -0.0154776
+ 1.622e+11Hz -0.018456 -0.0154745
+ 1.623e+11Hz -0.0184622 -0.0154714
+ 1.624e+11Hz -0.0184683 -0.0154684
+ 1.625e+11Hz -0.0184745 -0.0154655
+ 1.626e+11Hz -0.0184807 -0.0154627
+ 1.627e+11Hz -0.018487 -0.0154599
+ 1.628e+11Hz -0.0184933 -0.0154572
+ 1.629e+11Hz -0.0184996 -0.0154546
+ 1.63e+11Hz -0.0185059 -0.015452
+ 1.631e+11Hz -0.0185123 -0.0154495
+ 1.632e+11Hz -0.0185187 -0.0154471
+ 1.633e+11Hz -0.0185252 -0.0154447
+ 1.634e+11Hz -0.0185317 -0.0154424
+ 1.635e+11Hz -0.0185383 -0.0154402
+ 1.636e+11Hz -0.0185448 -0.015438
+ 1.637e+11Hz -0.0185515 -0.0154359
+ 1.638e+11Hz -0.0185582 -0.0154339
+ 1.639e+11Hz -0.0185649 -0.0154319
+ 1.64e+11Hz -0.0185716 -0.01543
+ 1.641e+11Hz -0.0185785 -0.0154281
+ 1.642e+11Hz -0.0185853 -0.0154264
+ 1.643e+11Hz -0.0185922 -0.0154247
+ 1.644e+11Hz -0.0185992 -0.015423
+ 1.645e+11Hz -0.0186062 -0.0154214
+ 1.646e+11Hz -0.0186132 -0.0154199
+ 1.647e+11Hz -0.0186204 -0.0154184
+ 1.648e+11Hz -0.0186275 -0.015417
+ 1.649e+11Hz -0.0186347 -0.0154157
+ 1.65e+11Hz -0.018642 -0.0154144
+ 1.651e+11Hz -0.0186494 -0.0154132
+ 1.652e+11Hz -0.0186567 -0.015412
+ 1.653e+11Hz -0.0186642 -0.0154109
+ 1.654e+11Hz -0.0186717 -0.0154098
+ 1.655e+11Hz -0.0186793 -0.0154088
+ 1.656e+11Hz -0.0186869 -0.0154079
+ 1.657e+11Hz -0.0186946 -0.015407
+ 1.658e+11Hz -0.0187023 -0.0154062
+ 1.659e+11Hz -0.0187102 -0.0154054
+ 1.66e+11Hz -0.0187181 -0.0154047
+ 1.661e+11Hz -0.018726 -0.015404
+ 1.662e+11Hz -0.018734 -0.0154034
+ 1.663e+11Hz -0.0187421 -0.0154028
+ 1.664e+11Hz -0.0187503 -0.0154023
+ 1.665e+11Hz -0.0187585 -0.0154018
+ 1.666e+11Hz -0.0187668 -0.0154014
+ 1.667e+11Hz -0.0187751 -0.0154011
+ 1.668e+11Hz -0.0187836 -0.0154007
+ 1.669e+11Hz -0.0187921 -0.0154005
+ 1.67e+11Hz -0.0188007 -0.0154002
+ 1.671e+11Hz -0.0188093 -0.0154
+ 1.672e+11Hz -0.0188181 -0.0153999
+ 1.673e+11Hz -0.0188269 -0.0153998
+ 1.674e+11Hz -0.0188358 -0.0153997
+ 1.675e+11Hz -0.0188447 -0.0153997
+ 1.676e+11Hz -0.0188538 -0.0153997
+ 1.677e+11Hz -0.0188629 -0.0153998
+ 1.678e+11Hz -0.0188721 -0.0153999
+ 1.679e+11Hz -0.0188814 -0.0154
+ 1.68e+11Hz -0.0188908 -0.0154002
+ 1.681e+11Hz -0.0189002 -0.0154004
+ 1.682e+11Hz -0.0189097 -0.0154007
+ 1.683e+11Hz -0.0189194 -0.015401
+ 1.684e+11Hz -0.0189291 -0.0154013
+ 1.685e+11Hz -0.0189388 -0.0154016
+ 1.686e+11Hz -0.0189487 -0.015402
+ 1.687e+11Hz -0.0189587 -0.0154024
+ 1.688e+11Hz -0.0189687 -0.0154028
+ 1.689e+11Hz -0.0189789 -0.0154033
+ 1.69e+11Hz -0.0189891 -0.0154037
+ 1.691e+11Hz -0.0189994 -0.0154043
+ 1.692e+11Hz -0.0190098 -0.0154048
+ 1.693e+11Hz -0.0190203 -0.0154053
+ 1.694e+11Hz -0.0190309 -0.0154059
+ 1.695e+11Hz -0.0190415 -0.0154065
+ 1.696e+11Hz -0.0190523 -0.0154071
+ 1.697e+11Hz -0.0190632 -0.0154078
+ 1.698e+11Hz -0.0190741 -0.0154084
+ 1.699e+11Hz -0.0190852 -0.0154091
+ 1.7e+11Hz -0.0190963 -0.0154098
+ 1.701e+11Hz -0.0191075 -0.0154105
+ 1.702e+11Hz -0.0191189 -0.0154112
+ 1.703e+11Hz -0.0191303 -0.0154119
+ 1.704e+11Hz -0.0191418 -0.0154126
+ 1.705e+11Hz -0.0191534 -0.0154133
+ 1.706e+11Hz -0.0191651 -0.0154141
+ 1.707e+11Hz -0.0191769 -0.0154148
+ 1.708e+11Hz -0.0191889 -0.0154156
+ 1.709e+11Hz -0.0192009 -0.0154163
+ 1.71e+11Hz -0.019213 -0.0154171
+ 1.711e+11Hz -0.0192252 -0.0154179
+ 1.712e+11Hz -0.0192375 -0.0154186
+ 1.713e+11Hz -0.0192499 -0.0154194
+ 1.714e+11Hz -0.0192623 -0.0154201
+ 1.715e+11Hz -0.0192749 -0.0154209
+ 1.716e+11Hz -0.0192876 -0.0154216
+ 1.717e+11Hz -0.0193004 -0.0154224
+ 1.718e+11Hz -0.0193133 -0.0154231
+ 1.719e+11Hz -0.0193263 -0.0154238
+ 1.72e+11Hz -0.0193394 -0.0154246
+ 1.721e+11Hz -0.0193526 -0.0154253
+ 1.722e+11Hz -0.0193659 -0.015426
+ 1.723e+11Hz -0.0193793 -0.0154266
+ 1.724e+11Hz -0.0193928 -0.0154273
+ 1.725e+11Hz -0.0194064 -0.0154279
+ 1.726e+11Hz -0.0194201 -0.0154285
+ 1.727e+11Hz -0.0194339 -0.0154292
+ 1.728e+11Hz -0.0194478 -0.0154297
+ 1.729e+11Hz -0.0194618 -0.0154303
+ 1.73e+11Hz -0.0194759 -0.0154308
+ 1.731e+11Hz -0.0194901 -0.0154313
+ 1.732e+11Hz -0.0195044 -0.0154318
+ 1.733e+11Hz -0.0195188 -0.0154323
+ 1.734e+11Hz -0.0195334 -0.0154327
+ 1.735e+11Hz -0.019548 -0.0154331
+ 1.736e+11Hz -0.0195627 -0.0154335
+ 1.737e+11Hz -0.0195775 -0.0154338
+ 1.738e+11Hz -0.0195924 -0.0154341
+ 1.739e+11Hz -0.0196074 -0.0154343
+ 1.74e+11Hz -0.0196225 -0.0154346
+ 1.741e+11Hz -0.0196377 -0.0154348
+ 1.742e+11Hz -0.019653 -0.0154349
+ 1.743e+11Hz -0.0196684 -0.015435
+ 1.744e+11Hz -0.0196839 -0.0154351
+ 1.745e+11Hz -0.0196995 -0.0154351
+ 1.746e+11Hz -0.0197153 -0.015435
+ 1.747e+11Hz -0.0197311 -0.015435
+ 1.748e+11Hz -0.019747 -0.0154348
+ 1.749e+11Hz -0.019763 -0.0154347
+ 1.75e+11Hz -0.019779 -0.0154344
+ 1.751e+11Hz -0.0197952 -0.0154342
+ 1.752e+11Hz -0.0198115 -0.0154338
+ 1.753e+11Hz -0.0198279 -0.0154335
+ 1.754e+11Hz -0.0198444 -0.015433
+ 1.755e+11Hz -0.019861 -0.0154325
+ 1.756e+11Hz -0.0198776 -0.015432
+ 1.757e+11Hz -0.0198944 -0.0154313
+ 1.758e+11Hz -0.0199112 -0.0154307
+ 1.759e+11Hz -0.0199282 -0.0154299
+ 1.76e+11Hz -0.0199452 -0.0154291
+ 1.761e+11Hz -0.0199624 -0.0154283
+ 1.762e+11Hz -0.0199796 -0.0154273
+ 1.763e+11Hz -0.0199969 -0.0154263
+ 1.764e+11Hz -0.0200143 -0.0154252
+ 1.765e+11Hz -0.0200318 -0.0154241
+ 1.766e+11Hz -0.0200494 -0.0154229
+ 1.767e+11Hz -0.020067 -0.0154216
+ 1.768e+11Hz -0.0200848 -0.0154202
+ 1.769e+11Hz -0.0201026 -0.0154188
+ 1.77e+11Hz -0.0201206 -0.0154173
+ 1.771e+11Hz -0.0201386 -0.0154157
+ 1.772e+11Hz -0.0201567 -0.015414
+ 1.773e+11Hz -0.0201749 -0.0154123
+ 1.774e+11Hz -0.0201931 -0.0154105
+ 1.775e+11Hz -0.0202115 -0.0154086
+ 1.776e+11Hz -0.0202299 -0.0154066
+ 1.777e+11Hz -0.0202484 -0.0154045
+ 1.778e+11Hz -0.020267 -0.0154023
+ 1.779e+11Hz -0.0202857 -0.0154001
+ 1.78e+11Hz -0.0203044 -0.0153977
+ 1.781e+11Hz -0.0203232 -0.0153953
+ 1.782e+11Hz -0.0203421 -0.0153928
+ 1.783e+11Hz -0.0203611 -0.0153902
+ 1.784e+11Hz -0.0203801 -0.0153875
+ 1.785e+11Hz -0.0203993 -0.0153847
+ 1.786e+11Hz -0.0204184 -0.0153818
+ 1.787e+11Hz -0.0204377 -0.0153788
+ 1.788e+11Hz -0.020457 -0.0153757
+ 1.789e+11Hz -0.0204764 -0.0153726
+ 1.79e+11Hz -0.0204959 -0.0153693
+ 1.791e+11Hz -0.0205154 -0.0153659
+ 1.792e+11Hz -0.020535 -0.0153624
+ 1.793e+11Hz -0.0205547 -0.0153589
+ 1.794e+11Hz -0.0205744 -0.0153552
+ 1.795e+11Hz -0.0205942 -0.0153514
+ 1.796e+11Hz -0.0206141 -0.0153475
+ 1.797e+11Hz -0.020634 -0.0153435
+ 1.798e+11Hz -0.020654 -0.0153394
+ 1.799e+11Hz -0.020674 -0.0153352
+ 1.8e+11Hz -0.0206941 -0.0153309
+ 1.801e+11Hz -0.0207143 -0.0153265
+ 1.802e+11Hz -0.0207345 -0.015322
+ 1.803e+11Hz -0.0207547 -0.0153174
+ 1.804e+11Hz -0.020775 -0.0153126
+ 1.805e+11Hz -0.0207954 -0.0153078
+ 1.806e+11Hz -0.0208158 -0.0153028
+ 1.807e+11Hz -0.0208363 -0.0152977
+ 1.808e+11Hz -0.0208568 -0.0152925
+ 1.809e+11Hz -0.0208773 -0.0152872
+ 1.81e+11Hz -0.0208979 -0.0152818
+ 1.811e+11Hz -0.0209186 -0.0152762
+ 1.812e+11Hz -0.0209392 -0.0152706
+ 1.813e+11Hz -0.02096 -0.0152648
+ 1.814e+11Hz -0.0209807 -0.0152589
+ 1.815e+11Hz -0.0210015 -0.0152529
+ 1.816e+11Hz -0.0210224 -0.0152467
+ 1.817e+11Hz -0.0210433 -0.0152405
+ 1.818e+11Hz -0.0210642 -0.0152341
+ 1.819e+11Hz -0.0210851 -0.0152276
+ 1.82e+11Hz -0.0211061 -0.015221
+ 1.821e+11Hz -0.0211271 -0.0152143
+ 1.822e+11Hz -0.0211481 -0.0152074
+ 1.823e+11Hz -0.0211692 -0.0152004
+ 1.824e+11Hz -0.0211903 -0.0151933
+ 1.825e+11Hz -0.0212114 -0.0151861
+ 1.826e+11Hz -0.0212325 -0.0151787
+ 1.827e+11Hz -0.0212537 -0.0151712
+ 1.828e+11Hz -0.0212749 -0.0151636
+ 1.829e+11Hz -0.0212961 -0.0151559
+ 1.83e+11Hz -0.0213173 -0.015148
+ 1.831e+11Hz -0.0213385 -0.0151401
+ 1.832e+11Hz -0.0213598 -0.015132
+ 1.833e+11Hz -0.021381 -0.0151237
+ 1.834e+11Hz -0.0214023 -0.0151154
+ 1.835e+11Hz -0.0214236 -0.0151069
+ 1.836e+11Hz -0.0214449 -0.0150982
+ 1.837e+11Hz -0.0214662 -0.0150895
+ 1.838e+11Hz -0.0214875 -0.0150806
+ 1.839e+11Hz -0.0215088 -0.0150716
+ 1.84e+11Hz -0.0215301 -0.0150625
+ 1.841e+11Hz -0.0215515 -0.0150532
+ 1.842e+11Hz -0.0215728 -0.0150438
+ 1.843e+11Hz -0.0215941 -0.0150343
+ 1.844e+11Hz -0.0216154 -0.0150247
+ 1.845e+11Hz -0.0216367 -0.0150149
+ 1.846e+11Hz -0.021658 -0.015005
+ 1.847e+11Hz -0.0216793 -0.014995
+ 1.848e+11Hz -0.0217006 -0.0149848
+ 1.849e+11Hz -0.0217219 -0.0149745
+ 1.85e+11Hz -0.0217432 -0.0149641
+ 1.851e+11Hz -0.0217644 -0.0149536
+ 1.852e+11Hz -0.0217857 -0.0149429
+ 1.853e+11Hz -0.0218069 -0.0149321
+ 1.854e+11Hz -0.0218281 -0.0149212
+ 1.855e+11Hz -0.0218493 -0.0149101
+ 1.856e+11Hz -0.0218705 -0.0148989
+ 1.857e+11Hz -0.0218916 -0.0148876
+ 1.858e+11Hz -0.0219128 -0.0148761
+ 1.859e+11Hz -0.0219339 -0.0148646
+ 1.86e+11Hz -0.0219549 -0.0148529
+ 1.861e+11Hz -0.021976 -0.014841
+ 1.862e+11Hz -0.021997 -0.0148291
+ 1.863e+11Hz -0.022018 -0.014817
+ 1.864e+11Hz -0.022039 -0.0148048
+ 1.865e+11Hz -0.0220599 -0.0147925
+ 1.866e+11Hz -0.0220808 -0.01478
+ 1.867e+11Hz -0.0221016 -0.0147674
+ 1.868e+11Hz -0.0221224 -0.0147547
+ 1.869e+11Hz -0.0221432 -0.0147419
+ 1.87e+11Hz -0.0221639 -0.0147289
+ 1.871e+11Hz -0.0221846 -0.0147158
+ 1.872e+11Hz -0.0222053 -0.0147026
+ 1.873e+11Hz -0.0222259 -0.0146893
+ 1.874e+11Hz -0.0222464 -0.0146758
+ 1.875e+11Hz -0.0222669 -0.0146623
+ 1.876e+11Hz -0.0222874 -0.0146486
+ 1.877e+11Hz -0.0223078 -0.0146348
+ 1.878e+11Hz -0.0223282 -0.0146208
+ 1.879e+11Hz -0.0223485 -0.0146068
+ 1.88e+11Hz -0.0223687 -0.0145926
+ 1.881e+11Hz -0.0223889 -0.0145783
+ 1.882e+11Hz -0.022409 -0.0145639
+ 1.883e+11Hz -0.0224291 -0.0145494
+ 1.884e+11Hz -0.0224491 -0.0145347
+ 1.885e+11Hz -0.0224691 -0.01452
+ 1.886e+11Hz -0.022489 -0.0145051
+ 1.887e+11Hz -0.0225088 -0.0144901
+ 1.888e+11Hz -0.0225286 -0.014475
+ 1.889e+11Hz -0.0225482 -0.0144598
+ 1.89e+11Hz -0.0225679 -0.0144445
+ 1.891e+11Hz -0.0225874 -0.0144291
+ 1.892e+11Hz -0.0226069 -0.0144135
+ 1.893e+11Hz -0.0226263 -0.0143979
+ 1.894e+11Hz -0.0226457 -0.0143821
+ 1.895e+11Hz -0.0226649 -0.0143663
+ 1.896e+11Hz -0.0226841 -0.0143503
+ 1.897e+11Hz -0.0227032 -0.0143342
+ 1.898e+11Hz -0.0227223 -0.014318
+ 1.899e+11Hz -0.0227412 -0.0143017
+ 1.9e+11Hz -0.0227601 -0.0142854
+ 1.901e+11Hz -0.0227789 -0.0142689
+ 1.902e+11Hz -0.0227976 -0.0142523
+ 1.903e+11Hz -0.0228162 -0.0142356
+ 1.904e+11Hz -0.0228348 -0.0142188
+ 1.905e+11Hz -0.0228532 -0.0142019
+ 1.906e+11Hz -0.0228716 -0.014185
+ 1.907e+11Hz -0.0228899 -0.0141679
+ 1.908e+11Hz -0.0229081 -0.0141507
+ 1.909e+11Hz -0.0229262 -0.0141335
+ 1.91e+11Hz -0.0229442 -0.0141161
+ 1.911e+11Hz -0.0229621 -0.0140987
+ 1.912e+11Hz -0.0229799 -0.0140812
+ 1.913e+11Hz -0.0229976 -0.0140635
+ 1.914e+11Hz -0.0230153 -0.0140458
+ 1.915e+11Hz -0.0230328 -0.014028
+ 1.916e+11Hz -0.0230503 -0.0140102
+ 1.917e+11Hz -0.0230676 -0.0139922
+ 1.918e+11Hz -0.0230848 -0.0139742
+ 1.919e+11Hz -0.023102 -0.0139561
+ 1.92e+11Hz -0.023119 -0.0139379
+ 1.921e+11Hz -0.023136 -0.0139196
+ 1.922e+11Hz -0.0231528 -0.0139013
+ 1.923e+11Hz -0.0231695 -0.0138828
+ 1.924e+11Hz -0.0231862 -0.0138644
+ 1.925e+11Hz -0.0232027 -0.0138458
+ 1.926e+11Hz -0.0232191 -0.0138271
+ 1.927e+11Hz -0.0232354 -0.0138084
+ 1.928e+11Hz -0.0232516 -0.0137897
+ 1.929e+11Hz -0.0232677 -0.0137708
+ 1.93e+11Hz -0.0232837 -0.0137519
+ 1.931e+11Hz -0.0232996 -0.013733
+ 1.932e+11Hz -0.0233154 -0.0137139
+ 1.933e+11Hz -0.0233311 -0.0136948
+ 1.934e+11Hz -0.0233466 -0.0136757
+ 1.935e+11Hz -0.0233621 -0.0136565
+ 1.936e+11Hz -0.0233774 -0.0136372
+ 1.937e+11Hz -0.0233926 -0.0136179
+ 1.938e+11Hz -0.0234077 -0.0135985
+ 1.939e+11Hz -0.0234227 -0.0135791
+ 1.94e+11Hz -0.0234376 -0.0135596
+ 1.941e+11Hz -0.0234523 -0.0135401
+ 1.942e+11Hz -0.023467 -0.0135206
+ 1.943e+11Hz -0.0234815 -0.0135009
+ 1.944e+11Hz -0.0234959 -0.0134813
+ 1.945e+11Hz -0.0235102 -0.0134616
+ 1.946e+11Hz -0.0235244 -0.0134419
+ 1.947e+11Hz -0.0235385 -0.0134221
+ 1.948e+11Hz -0.0235525 -0.0134023
+ 1.949e+11Hz -0.0235663 -0.0133824
+ 1.95e+11Hz -0.02358 -0.0133625
+ 1.951e+11Hz -0.0235936 -0.0133426
+ 1.952e+11Hz -0.0236071 -0.0133227
+ 1.953e+11Hz -0.0236205 -0.0133027
+ 1.954e+11Hz -0.0236337 -0.0132827
+ 1.955e+11Hz -0.0236469 -0.0132627
+ 1.956e+11Hz -0.0236599 -0.0132426
+ 1.957e+11Hz -0.0236728 -0.0132226
+ 1.958e+11Hz -0.0236856 -0.0132025
+ 1.959e+11Hz -0.0236982 -0.0131824
+ 1.96e+11Hz -0.0237108 -0.0131622
+ 1.961e+11Hz -0.0237232 -0.0131421
+ 1.962e+11Hz -0.0237355 -0.0131219
+ 1.963e+11Hz -0.0237477 -0.0131018
+ 1.964e+11Hz -0.0237598 -0.0130816
+ 1.965e+11Hz -0.0237718 -0.0130614
+ 1.966e+11Hz -0.0237836 -0.0130412
+ 1.967e+11Hz -0.0237953 -0.013021
+ 1.968e+11Hz -0.0238069 -0.0130008
+ 1.969e+11Hz -0.0238184 -0.0129806
+ 1.97e+11Hz -0.0238298 -0.0129604
+ 1.971e+11Hz -0.0238411 -0.0129402
+ 1.972e+11Hz -0.0238522 -0.01292
+ 1.973e+11Hz -0.0238633 -0.0128998
+ 1.974e+11Hz -0.0238742 -0.0128796
+ 1.975e+11Hz -0.023885 -0.0128594
+ 1.976e+11Hz -0.0238957 -0.0128392
+ 1.977e+11Hz -0.0239063 -0.012819
+ 1.978e+11Hz -0.0239168 -0.0127989
+ 1.979e+11Hz -0.0239271 -0.0127787
+ 1.98e+11Hz -0.0239374 -0.0127586
+ 1.981e+11Hz -0.0239475 -0.0127385
+ 1.982e+11Hz -0.0239575 -0.0127184
+ 1.983e+11Hz -0.0239675 -0.0126984
+ 1.984e+11Hz -0.0239773 -0.0126783
+ 1.985e+11Hz -0.023987 -0.0126583
+ 1.986e+11Hz -0.0239966 -0.0126383
+ 1.987e+11Hz -0.0240061 -0.0126183
+ 1.988e+11Hz -0.0240155 -0.0125984
+ 1.989e+11Hz -0.0240247 -0.0125785
+ 1.99e+11Hz -0.0240339 -0.0125586
+ 1.991e+11Hz -0.024043 -0.0125388
+ 1.992e+11Hz -0.024052 -0.012519
+ 1.993e+11Hz -0.0240608 -0.0124992
+ 1.994e+11Hz -0.0240696 -0.0124795
+ 1.995e+11Hz -0.0240783 -0.0124598
+ 1.996e+11Hz -0.0240869 -0.0124401
+ 1.997e+11Hz -0.0240954 -0.0124205
+ 1.998e+11Hz -0.0241037 -0.0124009
+ 1.999e+11Hz -0.024112 -0.0123814
+ 2e+11Hz -0.0241202 -0.0123619
+ 2.001e+11Hz -0.0241283 -0.0123425
+ 2.002e+11Hz -0.0241364 -0.0123231
+ 2.003e+11Hz -0.0241443 -0.0123038
+ 2.004e+11Hz -0.0241521 -0.0122845
+ 2.005e+11Hz -0.0241599 -0.0122653
+ 2.006e+11Hz -0.0241675 -0.0122461
+ 2.007e+11Hz -0.0241751 -0.012227
+ 2.008e+11Hz -0.0241826 -0.0122079
+ 2.009e+11Hz -0.02419 -0.0121889
+ 2.01e+11Hz -0.0241974 -0.01217
+ 2.011e+11Hz -0.0242046 -0.0121511
+ 2.012e+11Hz -0.0242118 -0.0121323
+ 2.013e+11Hz -0.0242189 -0.0121136
+ 2.014e+11Hz -0.024226 -0.0120949
+ 2.015e+11Hz -0.0242329 -0.0120762
+ 2.016e+11Hz -0.0242398 -0.0120577
+ 2.017e+11Hz -0.0242466 -0.0120392
+ 2.018e+11Hz -0.0242534 -0.0120208
+ 2.019e+11Hz -0.0242601 -0.0120024
+ 2.02e+11Hz -0.0242667 -0.0119841
+ 2.021e+11Hz -0.0242732 -0.0119659
+ 2.022e+11Hz -0.0242797 -0.0119478
+ 2.023e+11Hz -0.0242861 -0.0119297
+ 2.024e+11Hz -0.0242925 -0.0119118
+ 2.025e+11Hz -0.0242988 -0.0118938
+ 2.026e+11Hz -0.0243051 -0.011876
+ 2.027e+11Hz -0.0243113 -0.0118582
+ 2.028e+11Hz -0.0243175 -0.0118406
+ 2.029e+11Hz -0.0243236 -0.011823
+ 2.03e+11Hz -0.0243296 -0.0118054
+ 2.031e+11Hz -0.0243357 -0.011788
+ 2.032e+11Hz -0.0243416 -0.0117706
+ 2.033e+11Hz -0.0243476 -0.0117533
+ 2.034e+11Hz -0.0243535 -0.0117361
+ 2.035e+11Hz -0.0243593 -0.011719
+ 2.036e+11Hz -0.0243651 -0.011702
+ 2.037e+11Hz -0.0243709 -0.011685
+ 2.038e+11Hz -0.0243767 -0.0116682
+ 2.039e+11Hz -0.0243824 -0.0116514
+ 2.04e+11Hz -0.0243881 -0.0116347
+ 2.041e+11Hz -0.0243938 -0.0116181
+ 2.042e+11Hz -0.0243994 -0.0116016
+ 2.043e+11Hz -0.024405 -0.0115851
+ 2.044e+11Hz -0.0244106 -0.0115688
+ 2.045e+11Hz -0.0244162 -0.0115525
+ 2.046e+11Hz -0.0244218 -0.0115363
+ 2.047e+11Hz -0.0244273 -0.0115202
+ 2.048e+11Hz -0.0244329 -0.0115042
+ 2.049e+11Hz -0.0244384 -0.0114883
+ 2.05e+11Hz -0.0244439 -0.0114724
+ 2.051e+11Hz -0.0244495 -0.0114567
+ 2.052e+11Hz -0.024455 -0.011441
+ 2.053e+11Hz -0.0244605 -0.0114254
+ 2.054e+11Hz -0.024466 -0.0114099
+ 2.055e+11Hz -0.0244715 -0.0113945
+ 2.056e+11Hz -0.0244771 -0.0113792
+ 2.057e+11Hz -0.0244826 -0.011364
+ 2.058e+11Hz -0.0244881 -0.0113489
+ 2.059e+11Hz -0.0244937 -0.0113338
+ 2.06e+11Hz -0.0244993 -0.0113188
+ 2.061e+11Hz -0.0245049 -0.0113039
+ 2.062e+11Hz -0.0245105 -0.0112891
+ 2.063e+11Hz -0.0245161 -0.0112744
+ 2.064e+11Hz -0.0245217 -0.0112598
+ 2.065e+11Hz -0.0245274 -0.0112452
+ 2.066e+11Hz -0.0245331 -0.0112307
+ 2.067e+11Hz -0.0245389 -0.0112163
+ 2.068e+11Hz -0.0245446 -0.011202
+ 2.069e+11Hz -0.0245504 -0.0111878
+ 2.07e+11Hz -0.0245563 -0.0111737
+ 2.071e+11Hz -0.0245621 -0.0111596
+ 2.072e+11Hz -0.024568 -0.0111456
+ 2.073e+11Hz -0.024574 -0.0111317
+ 2.074e+11Hz -0.02458 -0.0111178
+ 2.075e+11Hz -0.0245861 -0.0111041
+ 2.076e+11Hz -0.0245921 -0.0110904
+ 2.077e+11Hz -0.0245983 -0.0110768
+ 2.078e+11Hz -0.0246045 -0.0110632
+ 2.079e+11Hz -0.0246107 -0.0110497
+ 2.08e+11Hz -0.0246171 -0.0110363
+ 2.081e+11Hz -0.0246234 -0.011023
+ 2.082e+11Hz -0.0246299 -0.0110097
+ 2.083e+11Hz -0.0246364 -0.0109965
+ 2.084e+11Hz -0.0246429 -0.0109834
+ 2.085e+11Hz -0.0246496 -0.0109703
+ 2.086e+11Hz -0.0246563 -0.0109573
+ 2.087e+11Hz -0.024663 -0.0109444
+ 2.088e+11Hz -0.0246699 -0.0109315
+ 2.089e+11Hz -0.0246768 -0.0109186
+ 2.09e+11Hz -0.0246838 -0.0109058
+ 2.091e+11Hz -0.0246909 -0.0108931
+ 2.092e+11Hz -0.024698 -0.0108804
+ 2.093e+11Hz -0.0247053 -0.0108678
+ 2.094e+11Hz -0.0247126 -0.0108553
+ 2.095e+11Hz -0.02472 -0.0108427
+ 2.096e+11Hz -0.0247275 -0.0108302
+ 2.097e+11Hz -0.0247351 -0.0108178
+ 2.098e+11Hz -0.0247428 -0.0108054
+ 2.099e+11Hz -0.0247505 -0.0107931
+ 2.1e+11Hz -0.0247584 -0.0107807
+ 2.101e+11Hz -0.0247664 -0.0107685
+ 2.102e+11Hz -0.0247744 -0.0107562
+ 2.103e+11Hz -0.0247826 -0.010744
+ 2.104e+11Hz -0.0247909 -0.0107318
+ 2.105e+11Hz -0.0247992 -0.0107197
+ 2.106e+11Hz -0.0248077 -0.0107075
+ 2.107e+11Hz -0.0248163 -0.0106954
+ 2.108e+11Hz -0.024825 -0.0106833
+ 2.109e+11Hz -0.0248338 -0.0106712
+ 2.11e+11Hz -0.0248427 -0.0106592
+ 2.111e+11Hz -0.0248517 -0.0106472
+ 2.112e+11Hz -0.0248608 -0.0106351
+ 2.113e+11Hz -0.02487 -0.0106231
+ 2.114e+11Hz -0.0248794 -0.0106111
+ 2.115e+11Hz -0.0248889 -0.0105991
+ 2.116e+11Hz -0.0248985 -0.0105871
+ 2.117e+11Hz -0.0249082 -0.0105751
+ 2.118e+11Hz -0.024918 -0.010563
+ 2.119e+11Hz -0.024928 -0.010551
+ 2.12e+11Hz -0.024938 -0.010539
+ 2.121e+11Hz -0.0249482 -0.0105269
+ 2.122e+11Hz -0.0249586 -0.0105149
+ 2.123e+11Hz -0.024969 -0.0105028
+ 2.124e+11Hz -0.0249796 -0.0104907
+ 2.125e+11Hz -0.0249903 -0.0104786
+ 2.126e+11Hz -0.0250011 -0.0104665
+ 2.127e+11Hz -0.025012 -0.0104543
+ 2.128e+11Hz -0.0250231 -0.0104421
+ 2.129e+11Hz -0.0250343 -0.0104299
+ 2.13e+11Hz -0.0250456 -0.0104176
+ 2.131e+11Hz -0.0250571 -0.0104053
+ 2.132e+11Hz -0.0250687 -0.0103929
+ 2.133e+11Hz -0.0250804 -0.0103805
+ 2.134e+11Hz -0.0250923 -0.0103681
+ 2.135e+11Hz -0.0251043 -0.0103556
+ 2.136e+11Hz -0.0251164 -0.010343
+ 2.137e+11Hz -0.0251286 -0.0103304
+ 2.138e+11Hz -0.025141 -0.0103177
+ 2.139e+11Hz -0.0251535 -0.010305
+ 2.14e+11Hz -0.0251661 -0.0102922
+ 2.141e+11Hz -0.0251789 -0.0102793
+ 2.142e+11Hz -0.0251918 -0.0102663
+ 2.143e+11Hz -0.0252048 -0.0102533
+ 2.144e+11Hz -0.025218 -0.0102402
+ 2.145e+11Hz -0.0252313 -0.010227
+ 2.146e+11Hz -0.0252447 -0.0102137
+ 2.147e+11Hz -0.0252583 -0.0102004
+ 2.148e+11Hz -0.0252719 -0.0101869
+ 2.149e+11Hz -0.0252857 -0.0101733
+ 2.15e+11Hz -0.0252997 -0.0101597
+ 2.151e+11Hz -0.0253137 -0.0101459
+ 2.152e+11Hz -0.0253279 -0.0101321
+ 2.153e+11Hz -0.0253422 -0.0101181
+ 2.154e+11Hz -0.0253567 -0.010104
+ 2.155e+11Hz -0.0253713 -0.0100898
+ 2.156e+11Hz -0.0253859 -0.0100755
+ 2.157e+11Hz -0.0254008 -0.0100611
+ 2.158e+11Hz -0.0254157 -0.0100466
+ 2.159e+11Hz -0.0254307 -0.0100319
+ 2.16e+11Hz -0.0254459 -0.0100171
+ 2.161e+11Hz -0.0254612 -0.0100021
+ 2.162e+11Hz -0.0254766 -0.00998704
+ 2.163e+11Hz -0.0254921 -0.00997182
+ 2.164e+11Hz -0.0255078 -0.00995646
+ 2.165e+11Hz -0.0255235 -0.00994096
+ 2.166e+11Hz -0.0255394 -0.0099253
+ 2.167e+11Hz -0.0255553 -0.00990949
+ 2.168e+11Hz -0.0255714 -0.00989353
+ 2.169e+11Hz -0.0255876 -0.00987741
+ 2.17e+11Hz -0.0256039 -0.00986113
+ 2.171e+11Hz -0.0256203 -0.00984469
+ 2.172e+11Hz -0.0256368 -0.00982807
+ 2.173e+11Hz -0.0256533 -0.00981129
+ 2.174e+11Hz -0.02567 -0.00979434
+ 2.175e+11Hz -0.0256868 -0.00977721
+ 2.176e+11Hz -0.0257037 -0.0097599
+ 2.177e+11Hz -0.0257206 -0.00974241
+ 2.178e+11Hz -0.0257377 -0.00972474
+ 2.179e+11Hz -0.0257548 -0.00970688
+ 2.18e+11Hz -0.025772 -0.00968883
+ 2.181e+11Hz -0.0257893 -0.00967059
+ 2.182e+11Hz -0.0258067 -0.00965215
+ 2.183e+11Hz -0.0258242 -0.00963351
+ 2.184e+11Hz -0.0258417 -0.00961468
+ 2.185e+11Hz -0.0258593 -0.00959564
+ 2.186e+11Hz -0.025877 -0.00957639
+ 2.187e+11Hz -0.0258947 -0.00955694
+ 2.188e+11Hz -0.0259125 -0.00953728
+ 2.189e+11Hz -0.0259304 -0.0095174
+ 2.19e+11Hz -0.0259483 -0.00949731
+ 2.191e+11Hz -0.0259663 -0.00947699
+ 2.192e+11Hz -0.0259843 -0.00945646
+ 2.193e+11Hz -0.0260024 -0.00943571
+ 2.194e+11Hz -0.0260205 -0.00941473
+ 2.195e+11Hz -0.0260386 -0.00939352
+ 2.196e+11Hz -0.0260568 -0.00937209
+ 2.197e+11Hz -0.0260751 -0.00935042
+ 2.198e+11Hz -0.0260933 -0.00932852
+ 2.199e+11Hz -0.0261116 -0.00930638
+ 2.2e+11Hz -0.02613 -0.00928401
+ 2.201e+11Hz -0.0261483 -0.00926139
+ 2.202e+11Hz -0.0261667 -0.00923854
+ 2.203e+11Hz -0.0261851 -0.00921544
+ 2.204e+11Hz -0.0262035 -0.00919209
+ 2.205e+11Hz -0.0262219 -0.0091685
+ 2.206e+11Hz -0.0262403 -0.00914466
+ 2.207e+11Hz -0.0262587 -0.00912057
+ 2.208e+11Hz -0.0262771 -0.00909623
+ 2.209e+11Hz -0.0262955 -0.00907164
+ 2.21e+11Hz -0.0263139 -0.00904679
+ 2.211e+11Hz -0.0263323 -0.00902169
+ 2.212e+11Hz -0.0263506 -0.00899633
+ 2.213e+11Hz -0.026369 -0.00897071
+ 2.214e+11Hz -0.0263873 -0.00894483
+ 2.215e+11Hz -0.0264056 -0.00891869
+ 2.216e+11Hz -0.0264238 -0.00889229
+ 2.217e+11Hz -0.026442 -0.00886562
+ 2.218e+11Hz -0.0264602 -0.00883869
+ 2.219e+11Hz -0.0264783 -0.0088115
+ 2.22e+11Hz -0.0264964 -0.00878404
+ 2.221e+11Hz -0.0265144 -0.00875631
+ 2.222e+11Hz -0.0265324 -0.00872832
+ 2.223e+11Hz -0.0265503 -0.00870006
+ 2.224e+11Hz -0.0265682 -0.00867153
+ 2.225e+11Hz -0.0265859 -0.00864274
+ 2.226e+11Hz -0.0266036 -0.00861367
+ 2.227e+11Hz -0.0266213 -0.00858434
+ 2.228e+11Hz -0.0266388 -0.00855473
+ 2.229e+11Hz -0.0266563 -0.00852486
+ 2.23e+11Hz -0.0266736 -0.00849471
+ 2.231e+11Hz -0.0266909 -0.0084643
+ 2.232e+11Hz -0.0267081 -0.00843362
+ 2.233e+11Hz -0.0267251 -0.00840266
+ 2.234e+11Hz -0.0267421 -0.00837144
+ 2.235e+11Hz -0.0267589 -0.00833994
+ 2.236e+11Hz -0.0267757 -0.00830818
+ 2.237e+11Hz -0.0267923 -0.00827615
+ 2.238e+11Hz -0.0268087 -0.00824385
+ 2.239e+11Hz -0.0268251 -0.00821128
+ 2.24e+11Hz -0.0268413 -0.00817845
+ 2.241e+11Hz -0.0268574 -0.00814535
+ 2.242e+11Hz -0.0268733 -0.00811198
+ 2.243e+11Hz -0.0268891 -0.00807835
+ 2.244e+11Hz -0.0269047 -0.00804445
+ 2.245e+11Hz -0.0269202 -0.00801029
+ 2.246e+11Hz -0.0269355 -0.00797587
+ 2.247e+11Hz -0.0269507 -0.00794119
+ 2.248e+11Hz -0.0269657 -0.00790625
+ 2.249e+11Hz -0.0269805 -0.00787105
+ 2.25e+11Hz -0.0269951 -0.00783559
+ 2.251e+11Hz -0.0270096 -0.00779987
+ 2.252e+11Hz -0.0270238 -0.00776391
+ 2.253e+11Hz -0.0270379 -0.00772769
+ 2.254e+11Hz -0.0270518 -0.00769121
+ 2.255e+11Hz -0.0270655 -0.00765449
+ 2.256e+11Hz -0.027079 -0.00761752
+ 2.257e+11Hz -0.0270922 -0.00758031
+ 2.258e+11Hz -0.0271053 -0.00754285
+ 2.259e+11Hz -0.0271182 -0.00750515
+ 2.26e+11Hz -0.0271308 -0.00746721
+ 2.261e+11Hz -0.0271432 -0.00742904
+ 2.262e+11Hz -0.0271554 -0.00739062
+ 2.263e+11Hz -0.0271673 -0.00735198
+ 2.264e+11Hz -0.027179 -0.0073131
+ 2.265e+11Hz -0.0271905 -0.007274
+ 2.266e+11Hz -0.0272017 -0.00723467
+ 2.267e+11Hz -0.0272127 -0.00719512
+ 2.268e+11Hz -0.0272234 -0.00715534
+ 2.269e+11Hz -0.0272339 -0.00711535
+ 2.27e+11Hz -0.0272441 -0.00707515
+ 2.271e+11Hz -0.027254 -0.00703473
+ 2.272e+11Hz -0.0272637 -0.0069941
+ 2.273e+11Hz -0.0272731 -0.00695327
+ 2.274e+11Hz -0.0272823 -0.00691223
+ 2.275e+11Hz -0.0272911 -0.00687099
+ 2.276e+11Hz -0.0272997 -0.00682956
+ 2.277e+11Hz -0.027308 -0.00678793
+ 2.278e+11Hz -0.027316 -0.00674611
+ 2.279e+11Hz -0.0273237 -0.00670411
+ 2.28e+11Hz -0.0273311 -0.00666192
+ 2.281e+11Hz -0.0273383 -0.00661955
+ 2.282e+11Hz -0.0273451 -0.00657701
+ 2.283e+11Hz -0.0273516 -0.00653429
+ 2.284e+11Hz -0.0273578 -0.0064914
+ 2.285e+11Hz -0.0273637 -0.00644835
+ 2.286e+11Hz -0.0273693 -0.00640514
+ 2.287e+11Hz -0.0273746 -0.00636176
+ 2.288e+11Hz -0.0273795 -0.00631824
+ 2.289e+11Hz -0.0273841 -0.00627456
+ 2.29e+11Hz -0.0273884 -0.00623074
+ 2.291e+11Hz -0.0273924 -0.00618678
+ 2.292e+11Hz -0.0273961 -0.00614267
+ 2.293e+11Hz -0.0273994 -0.00609844
+ 2.294e+11Hz -0.0274024 -0.00605407
+ 2.295e+11Hz -0.027405 -0.00600958
+ 2.296e+11Hz -0.0274073 -0.00596497
+ 2.297e+11Hz -0.0274092 -0.00592024
+ 2.298e+11Hz -0.0274109 -0.0058754
+ 2.299e+11Hz -0.0274121 -0.00583045
+ 2.3e+11Hz -0.027413 -0.00578539
+ 2.301e+11Hz -0.0274136 -0.00574024
+ 2.302e+11Hz -0.0274138 -0.00569499
+ 2.303e+11Hz -0.0274137 -0.00564965
+ 2.304e+11Hz -0.0274131 -0.00560423
+ 2.305e+11Hz -0.0274123 -0.00555873
+ 2.306e+11Hz -0.0274111 -0.00551315
+ 2.307e+11Hz -0.0274095 -0.0054675
+ 2.308e+11Hz -0.0274075 -0.00542178
+ 2.309e+11Hz -0.0274052 -0.005376
+ 2.31e+11Hz -0.0274025 -0.00533016
+ 2.311e+11Hz -0.0273995 -0.00528427
+ 2.312e+11Hz -0.0273961 -0.00523833
+ 2.313e+11Hz -0.0273923 -0.00519235
+ 2.314e+11Hz -0.0273881 -0.00514633
+ 2.315e+11Hz -0.0273836 -0.00510028
+ 2.316e+11Hz -0.0273787 -0.0050542
+ 2.317e+11Hz -0.0273734 -0.0050081
+ 2.318e+11Hz -0.0273678 -0.00496198
+ 2.319e+11Hz -0.0273617 -0.00491584
+ 2.32e+11Hz -0.0273553 -0.0048697
+ 2.321e+11Hz -0.0273485 -0.00482355
+ 2.322e+11Hz -0.0273414 -0.00477741
+ 2.323e+11Hz -0.0273339 -0.00473127
+ 2.324e+11Hz -0.0273259 -0.00468514
+ 2.325e+11Hz -0.0273177 -0.00463904
+ 2.326e+11Hz -0.027309 -0.00459295
+ 2.327e+11Hz -0.0272999 -0.00454689
+ 2.328e+11Hz -0.0272905 -0.00450086
+ 2.329e+11Hz -0.0272807 -0.00445486
+ 2.33e+11Hz -0.0272705 -0.00440891
+ 2.331e+11Hz -0.02726 -0.00436301
+ 2.332e+11Hz -0.027249 -0.00431716
+ 2.333e+11Hz -0.0272377 -0.00427136
+ 2.334e+11Hz -0.0272261 -0.00422563
+ 2.335e+11Hz -0.027214 -0.00417996
+ 2.336e+11Hz -0.0272016 -0.00413437
+ 2.337e+11Hz -0.0271888 -0.00408885
+ 2.338e+11Hz -0.0271756 -0.00404342
+ 2.339e+11Hz -0.027162 -0.00399807
+ 2.34e+11Hz -0.0271481 -0.00395281
+ 2.341e+11Hz -0.0271338 -0.00390765
+ 2.342e+11Hz -0.0271191 -0.00386259
+ 2.343e+11Hz -0.0271041 -0.00381764
+ 2.344e+11Hz -0.0270887 -0.00377279
+ 2.345e+11Hz -0.027073 -0.00372807
+ 2.346e+11Hz -0.0270568 -0.00368346
+ 2.347e+11Hz -0.0270404 -0.00363898
+ 2.348e+11Hz -0.0270235 -0.00359464
+ 2.349e+11Hz -0.0270063 -0.00355042
+ 2.35e+11Hz -0.0269888 -0.00350635
+ 2.351e+11Hz -0.0269709 -0.00346242
+ 2.352e+11Hz -0.0269526 -0.00341864
+ 2.353e+11Hz -0.026934 -0.00337501
+ 2.354e+11Hz -0.026915 -0.00333154
+ 2.355e+11Hz -0.0268957 -0.00328823
+ 2.356e+11Hz -0.0268761 -0.00324509
+ 2.357e+11Hz -0.0268561 -0.00320213
+ 2.358e+11Hz -0.0268357 -0.00315934
+ 2.359e+11Hz -0.0268151 -0.00311673
+ 2.36e+11Hz -0.0267941 -0.0030743
+ 2.361e+11Hz -0.0267727 -0.00303206
+ 2.362e+11Hz -0.0267511 -0.00299002
+ 2.363e+11Hz -0.0267291 -0.00294817
+ 2.364e+11Hz -0.0267068 -0.00290653
+ 2.365e+11Hz -0.0266842 -0.00286509
+ 2.366e+11Hz -0.0266612 -0.00282386
+ 2.367e+11Hz -0.026638 -0.00278284
+ 2.368e+11Hz -0.0266144 -0.00274204
+ 2.369e+11Hz -0.0265905 -0.00270146
+ 2.37e+11Hz -0.0265663 -0.00266111
+ 2.371e+11Hz -0.0265418 -0.00262099
+ 2.372e+11Hz -0.026517 -0.0025811
+ 2.373e+11Hz -0.026492 -0.00254144
+ 2.374e+11Hz -0.0264666 -0.00250203
+ 2.375e+11Hz -0.0264409 -0.00246286
+ 2.376e+11Hz -0.026415 -0.00242394
+ 2.377e+11Hz -0.0263888 -0.00238526
+ 2.378e+11Hz -0.0263623 -0.00234684
+ 2.379e+11Hz -0.0263355 -0.00230868
+ 2.38e+11Hz -0.0263084 -0.00227078
+ 2.381e+11Hz -0.0262811 -0.00223314
+ 2.382e+11Hz -0.0262535 -0.00219577
+ 2.383e+11Hz -0.0262257 -0.00215867
+ 2.384e+11Hz -0.0261976 -0.00212184
+ 2.385e+11Hz -0.0261693 -0.00208528
+ 2.386e+11Hz -0.0261407 -0.00204901
+ 2.387e+11Hz -0.0261119 -0.00201301
+ 2.388e+11Hz -0.0260828 -0.0019773
+ 2.389e+11Hz -0.0260535 -0.00194187
+ 2.39e+11Hz -0.0260239 -0.00190674
+ 2.391e+11Hz -0.0259942 -0.00187189
+ 2.392e+11Hz -0.0259642 -0.00183734
+ 2.393e+11Hz -0.025934 -0.00180309
+ 2.394e+11Hz -0.0259036 -0.00176913
+ 2.395e+11Hz -0.0258729 -0.00173548
+ 2.396e+11Hz -0.0258421 -0.00170213
+ 2.397e+11Hz -0.0258111 -0.00166908
+ 2.398e+11Hz -0.0257798 -0.00163634
+ 2.399e+11Hz -0.0257484 -0.0016039
+ 2.4e+11Hz -0.0257168 -0.00157178
+ 2.401e+11Hz -0.025685 -0.00153997
+ 2.402e+11Hz -0.025653 -0.00150848
+ 2.403e+11Hz -0.0256209 -0.0014773
+ 2.404e+11Hz -0.0255886 -0.00144644
+ 2.405e+11Hz -0.0255561 -0.00141589
+ 2.406e+11Hz -0.0255234 -0.00138567
+ 2.407e+11Hz -0.0254906 -0.00135577
+ 2.408e+11Hz -0.0254577 -0.00132619
+ 2.409e+11Hz -0.0254246 -0.00129693
+ 2.41e+11Hz -0.0253913 -0.001268
+ 2.411e+11Hz -0.0253579 -0.0012394
+ 2.412e+11Hz -0.0253244 -0.00121112
+ 2.413e+11Hz -0.0252908 -0.00118317
+ 2.414e+11Hz -0.025257 -0.00115555
+ 2.415e+11Hz -0.0252231 -0.00112826
+ 2.416e+11Hz -0.0251891 -0.00110129
+ 2.417e+11Hz -0.025155 -0.00107466
+ 2.418e+11Hz -0.0251207 -0.00104836
+ 2.419e+11Hz -0.0250864 -0.00102239
+ 2.42e+11Hz -0.025052 -0.000996754
+ 2.421e+11Hz -0.0250174 -0.000971449
+ 2.422e+11Hz -0.0249828 -0.000946475
+ 2.423e+11Hz -0.0249481 -0.000921835
+ 2.424e+11Hz -0.0249134 -0.000897527
+ 2.425e+11Hz -0.0248785 -0.000873551
+ 2.426e+11Hz -0.0248436 -0.000849908
+ 2.427e+11Hz -0.0248086 -0.000826598
+ 2.428e+11Hz -0.0247735 -0.000803619
+ 2.429e+11Hz -0.0247384 -0.000780973
+ 2.43e+11Hz -0.0247033 -0.000758658
+ 2.431e+11Hz -0.0246681 -0.000736674
+ 2.432e+11Hz -0.0246328 -0.000715021
+ 2.433e+11Hz -0.0245975 -0.000693698
+ 2.434e+11Hz -0.0245622 -0.000672704
+ 2.435e+11Hz -0.0245268 -0.000652039
+ 2.436e+11Hz -0.0244914 -0.000631703
+ 2.437e+11Hz -0.024456 -0.000611694
+ 2.438e+11Hz -0.0244206 -0.000592011
+ 2.439e+11Hz -0.0243851 -0.000572654
+ 2.44e+11Hz -0.0243497 -0.000553621
+ 2.441e+11Hz -0.0243142 -0.000534912
+ 2.442e+11Hz -0.0242788 -0.000516525
+ 2.443e+11Hz -0.0242433 -0.000498459
+ 2.444e+11Hz -0.0242078 -0.000480714
+ 2.445e+11Hz -0.0241724 -0.000463287
+ 2.446e+11Hz -0.024137 -0.000446178
+ 2.447e+11Hz -0.0241015 -0.000429384
+ 2.448e+11Hz -0.0240662 -0.000412905
+ 2.449e+11Hz -0.0240308 -0.00039674
+ 2.45e+11Hz -0.0239955 -0.000380885
+ 2.451e+11Hz -0.0239601 -0.000365341
+ 2.452e+11Hz -0.0239249 -0.000350105
+ 2.453e+11Hz -0.0238897 -0.000335176
+ 2.454e+11Hz -0.0238545 -0.000320551
+ 2.455e+11Hz -0.0238193 -0.000306229
+ 2.456e+11Hz -0.0237843 -0.000292209
+ 2.457e+11Hz -0.0237492 -0.000278487
+ 2.458e+11Hz -0.0237143 -0.000265063
+ 2.459e+11Hz -0.0236794 -0.000251935
+ 2.46e+11Hz -0.0236445 -0.000239099
+ 2.461e+11Hz -0.0236097 -0.000226555
+ 2.462e+11Hz -0.023575 -0.0002143
+ 2.463e+11Hz -0.0235404 -0.000202332
+ 2.464e+11Hz -0.0235059 -0.000190649
+ 2.465e+11Hz -0.0234714 -0.000179248
+ 2.466e+11Hz -0.023437 -0.000168128
+ 2.467e+11Hz -0.0234027 -0.000157285
+ 2.468e+11Hz -0.0233685 -0.000146718
+ 2.469e+11Hz -0.0233344 -0.000136425
+ 2.47e+11Hz -0.0233004 -0.000126402
+ 2.471e+11Hz -0.0232665 -0.000116648
+ 2.472e+11Hz -0.0232327 -0.00010716
+ 2.473e+11Hz -0.023199 -9.7935e-05
+ 2.474e+11Hz -0.0231654 -8.89712e-05
+ 2.475e+11Hz -0.023132 -8.02658e-05
+ 2.476e+11Hz -0.0230986 -7.18163e-05
+ 2.477e+11Hz -0.0230653 -6.36199e-05
+ 2.478e+11Hz -0.0230322 -5.56742e-05
+ 2.479e+11Hz -0.0229992 -4.79764e-05
+ 2.48e+11Hz -0.0229663 -4.05238e-05
+ 2.481e+11Hz -0.0229336 -3.33139e-05
+ 2.482e+11Hz -0.0229009 -2.63438e-05
+ 2.483e+11Hz -0.0228684 -1.96108e-05
+ 2.484e+11Hz -0.0228361 -1.31123e-05
+ 2.485e+11Hz -0.0228038 -6.84528e-06
+ 2.486e+11Hz -0.0227717 -8.0713e-07
+ 2.487e+11Hz -0.0227398 5.005e-06
+ 2.488e+11Hz -0.022708 1.05939e-05
+ 2.489e+11Hz -0.0226763 1.59625e-05
+ 2.49e+11Hz -0.0226448 2.11135e-05
+ 2.491e+11Hz -0.0226134 2.60498e-05
+ 2.492e+11Hz -0.0225822 3.07743e-05
+ 2.493e+11Hz -0.0225511 3.52899e-05
+ 2.494e+11Hz -0.0225202 3.95994e-05
+ 2.495e+11Hz -0.0224894 4.37058e-05
+ 2.496e+11Hz -0.0224588 4.76118e-05
+ 2.497e+11Hz -0.0224284 5.13205e-05
+ 2.498e+11Hz -0.0223981 5.48347e-05
+ 2.499e+11Hz -0.0223679 5.81574e-05
+ 2.5e+11Hz -0.022338 6.12915e-05
+ 2.501e+11Hz -0.0223082 6.42398e-05
+ 2.502e+11Hz -0.0222785 6.70053e-05
+ 2.503e+11Hz -0.022249 6.9591e-05
+ 2.504e+11Hz -0.0222197 7.19997e-05
+ 2.505e+11Hz -0.0221906 7.42343e-05
+ 2.506e+11Hz -0.0221616 7.62979e-05
+ 2.507e+11Hz -0.0221328 7.81932e-05
+ 2.508e+11Hz -0.0221042 7.99233e-05
+ 2.509e+11Hz -0.0220758 8.1491e-05
+ 2.51e+11Hz -0.0220475 8.28993e-05
+ 2.511e+11Hz -0.0220194 8.4151e-05
+ 2.512e+11Hz -0.0219915 8.52491e-05
+ 2.513e+11Hz -0.0219637 8.61964e-05
+ 2.514e+11Hz -0.0219362 8.69958e-05
+ 2.515e+11Hz -0.0219088 8.76503e-05
+ 2.516e+11Hz -0.0218816 8.81626e-05
+ 2.517e+11Hz -0.0218545 8.85356e-05
+ 2.518e+11Hz -0.0218277 8.87723e-05
+ 2.519e+11Hz -0.021801 8.88754e-05
+ 2.52e+11Hz -0.0217745 8.88478e-05
+ 2.521e+11Hz -0.0217482 8.86923e-05
+ 2.522e+11Hz -0.0217221 8.84117e-05
+ 2.523e+11Hz -0.0216962 8.80088e-05
+ 2.524e+11Hz -0.0216704 8.74864e-05
+ 2.525e+11Hz -0.0216449 8.68474e-05
+ 2.526e+11Hz -0.0216195 8.60944e-05
+ 2.527e+11Hz -0.0215943 8.52302e-05
+ 2.528e+11Hz -0.0215693 8.42576e-05
+ 2.529e+11Hz -0.0215445 8.31793e-05
+ 2.53e+11Hz -0.0215198 8.1998e-05
+ 2.531e+11Hz -0.0214954 8.07164e-05
+ 2.532e+11Hz -0.0214711 7.93372e-05
+ 2.533e+11Hz -0.0214471 7.78631e-05
+ 2.534e+11Hz -0.0214232 7.62967e-05
+ 2.535e+11Hz -0.0213995 7.46407e-05
+ 2.536e+11Hz -0.021376 7.28978e-05
+ 2.537e+11Hz -0.0213526 7.10704e-05
+ 2.538e+11Hz -0.0213295 6.91612e-05
+ 2.539e+11Hz -0.0213066 6.71729e-05
+ 2.54e+11Hz -0.0212838 6.5108e-05
+ 2.541e+11Hz -0.0212612 6.29689e-05
+ 2.542e+11Hz -0.0212389 6.07584e-05
+ 2.543e+11Hz -0.0212167 5.84788e-05
+ 2.544e+11Hz -0.0211947 5.61327e-05
+ 2.545e+11Hz -0.0211728 5.37226e-05
+ 2.546e+11Hz -0.0211512 5.1251e-05
+ 2.547e+11Hz -0.0211298 4.87203e-05
+ 2.548e+11Hz -0.0211085 4.61329e-05
+ 2.549e+11Hz -0.0210874 4.34914e-05
+ 2.55e+11Hz -0.0210665 4.0798e-05
+ 2.551e+11Hz -0.0210458 3.80552e-05
+ 2.552e+11Hz -0.0210253 3.52655e-05
+ 2.553e+11Hz -0.021005 3.2431e-05
+ 2.554e+11Hz -0.0209849 2.95543e-05
+ 2.555e+11Hz -0.0209649 2.66376e-05
+ 2.556e+11Hz -0.0209451 2.36832e-05
+ 2.557e+11Hz -0.0209255 2.06935e-05
+ 2.558e+11Hz -0.0209061 1.76707e-05
+ 2.559e+11Hz -0.0208869 1.46172e-05
+ 2.56e+11Hz -0.0208679 1.15352e-05
+ 2.561e+11Hz -0.020849 8.42689e-06
+ 2.562e+11Hz -0.0208303 5.29458e-06
+ 2.563e+11Hz -0.0208119 2.14047e-06
+ 2.564e+11Hz -0.0207935 -1.03323e-06
+ 2.565e+11Hz -0.0207754 -4.22433e-06
+ 2.566e+11Hz -0.0207575 -7.43064e-06
+ 2.567e+11Hz -0.0207397 -1.065e-05
+ 2.568e+11Hz -0.0207221 -1.38802e-05
+ 2.569e+11Hz -0.0207047 -1.71192e-05
+ 2.57e+11Hz -0.0206875 -2.03647e-05
+ 2.571e+11Hz -0.0206704 -2.36147e-05
+ 2.572e+11Hz -0.0206535 -2.68671e-05
+ 2.573e+11Hz -0.0206368 -3.01198e-05
+ 2.574e+11Hz -0.0206203 -3.33706e-05
+ 2.575e+11Hz -0.020604 -3.66174e-05
+ 2.576e+11Hz -0.0205878 -3.98583e-05
+ 2.577e+11Hz -0.0205718 -4.30911e-05
+ 2.578e+11Hz -0.020556 -4.63138e-05
+ 2.579e+11Hz -0.0205403 -4.95243e-05
+ 2.58e+11Hz -0.0205248 -5.27206e-05
+ 2.581e+11Hz -0.0205095 -5.59006e-05
+ 2.582e+11Hz -0.0204944 -5.90624e-05
+ 2.583e+11Hz -0.0204794 -6.22039e-05
+ 2.584e+11Hz -0.0204646 -6.53231e-05
+ 2.585e+11Hz -0.02045 -6.8418e-05
+ 2.586e+11Hz -0.0204355 -7.14866e-05
+ 2.587e+11Hz -0.0204212 -7.45269e-05
+ 2.588e+11Hz -0.0204071 -7.75369e-05
+ 2.589e+11Hz -0.0203931 -8.05147e-05
+ 2.59e+11Hz -0.0203793 -8.34582e-05
+ 2.591e+11Hz -0.0203657 -8.63655e-05
+ 2.592e+11Hz -0.0203522 -8.92346e-05
+ 2.593e+11Hz -0.0203389 -9.20635e-05
+ 2.594e+11Hz -0.0203258 -9.48504e-05
+ 2.595e+11Hz -0.0203128 -9.75931e-05
+ 2.596e+11Hz -0.0203 -0.00010029
+ 2.597e+11Hz -0.0202874 -0.000102939
+ 2.598e+11Hz -0.0202749 -0.000105537
+ 2.599e+11Hz -0.0202625 -0.000108084
+ 2.6e+11Hz -0.0202503 -0.000110577
+ 2.601e+11Hz -0.0202383 -0.000113014
+ 2.602e+11Hz -0.0202264 -0.000115394
+ 2.603e+11Hz -0.0202147 -0.000117713
+ 2.604e+11Hz -0.0202032 -0.000119971
+ 2.605e+11Hz -0.0201917 -0.000122166
+ 2.606e+11Hz -0.0201805 -0.000124295
+ 2.607e+11Hz -0.0201694 -0.000126356
+ 2.608e+11Hz -0.0201584 -0.000128348
+ 2.609e+11Hz -0.0201476 -0.000130269
+ 2.61e+11Hz -0.020137 -0.000132116
+ 2.611e+11Hz -0.0201265 -0.000133888
+ 2.612e+11Hz -0.0201161 -0.000135583
+ 2.613e+11Hz -0.0201059 -0.000137198
+ 2.614e+11Hz -0.0200958 -0.000138732
+ 2.615e+11Hz -0.0200859 -0.000140183
+ 2.616e+11Hz -0.0200761 -0.00014155
+ 2.617e+11Hz -0.0200664 -0.000142829
+ 2.618e+11Hz -0.0200569 -0.000144019
+ 2.619e+11Hz -0.0200476 -0.000145118
+ 2.62e+11Hz -0.0200383 -0.000146124
+ 2.621e+11Hz -0.0200292 -0.000147035
+ 2.622e+11Hz -0.0200203 -0.000147849
+ 2.623e+11Hz -0.0200115 -0.000148565
+ 2.624e+11Hz -0.0200028 -0.000149179
+ 2.625e+11Hz -0.0199942 -0.000149691
+ 2.626e+11Hz -0.0199858 -0.000150098
+ 2.627e+11Hz -0.0199775 -0.000150399
+ 2.628e+11Hz -0.0199693 -0.00015059
+ 2.629e+11Hz -0.0199613 -0.000150671
+ 2.63e+11Hz -0.0199534 -0.00015064
+ 2.631e+11Hz -0.0199456 -0.000150493
+ 2.632e+11Hz -0.0199379 -0.00015023
+ 2.633e+11Hz -0.0199303 -0.000149848
+ 2.634e+11Hz -0.0199229 -0.000149346
+ 2.635e+11Hz -0.0199156 -0.000148721
+ 2.636e+11Hz -0.0199084 -0.000147972
+ 2.637e+11Hz -0.0199013 -0.000147096
+ 2.638e+11Hz -0.0198943 -0.000146091
+ 2.639e+11Hz -0.0198875 -0.000144956
+ 2.64e+11Hz -0.0198807 -0.000143689
+ 2.641e+11Hz -0.0198741 -0.000142287
+ 2.642e+11Hz -0.0198676 -0.000140749
+ 2.643e+11Hz -0.0198611 -0.000139072
+ 2.644e+11Hz -0.0198548 -0.000137255
+ 2.645e+11Hz -0.0198486 -0.000135296
+ 2.646e+11Hz -0.0198425 -0.000133192
+ 2.647e+11Hz -0.0198364 -0.000130943
+ 2.648e+11Hz -0.0198305 -0.000128545
+ 2.649e+11Hz -0.0198247 -0.000125997
+ 2.65e+11Hz -0.0198189 -0.000123297
+ 2.651e+11Hz -0.0198133 -0.000120444
+ 2.652e+11Hz -0.0198077 -0.000117434
+ 2.653e+11Hz -0.0198022 -0.000114267
+ 2.654e+11Hz -0.0197968 -0.00011094
+ 2.655e+11Hz -0.0197915 -0.000107452
+ 2.656e+11Hz -0.0197863 -0.0001038
+ 2.657e+11Hz -0.0197811 -9.99837e-05
+ 2.658e+11Hz -0.019776 -9.59999e-05
+ 2.659e+11Hz -0.019771 -9.18472e-05
+ 2.66e+11Hz -0.0197661 -8.75239e-05
+ 2.661e+11Hz -0.0197612 -8.30281e-05
+ 2.662e+11Hz -0.0197564 -7.83581e-05
+ 2.663e+11Hz -0.0197517 -7.3512e-05
+ 2.664e+11Hz -0.019747 -6.84882e-05
+ 2.665e+11Hz -0.0197424 -6.32849e-05
+ 2.666e+11Hz -0.0197378 -5.79003e-05
+ 2.667e+11Hz -0.0197333 -5.23329e-05
+ 2.668e+11Hz -0.0197288 -4.65809e-05
+ 2.669e+11Hz -0.0197244 -4.06428e-05
+ 2.67e+11Hz -0.01972 -3.45167e-05
+ 2.671e+11Hz -0.0197157 -2.82013e-05
+ 2.672e+11Hz -0.0197114 -2.16949e-05
+ 2.673e+11Hz -0.0197072 -1.49959e-05
+ 2.674e+11Hz -0.0197029 -8.10288e-06
+ 2.675e+11Hz -0.0196988 -1.0143e-06
+ 2.676e+11Hz -0.0196946 6.27128e-06
+ 2.677e+11Hz -0.0196905 1.37553e-05
+ 2.678e+11Hz -0.0196863 2.14392e-05
+ 2.679e+11Hz -0.0196822 2.93242e-05
+ 2.68e+11Hz -0.0196782 3.74118e-05
+ 2.681e+11Hz -0.0196741 4.57032e-05
+ 2.682e+11Hz -0.01967 5.41997e-05
+ 2.683e+11Hz -0.019666 6.29025e-05
+ 2.684e+11Hz -0.0196619 7.18128e-05
+ 2.685e+11Hz -0.0196579 8.09317e-05
+ 2.686e+11Hz -0.0196538 9.02604e-05
+ 2.687e+11Hz -0.0196498 9.97999e-05
+ 2.688e+11Hz -0.0196457 0.000109551
+ 2.689e+11Hz -0.0196416 0.000119515
+ 2.69e+11Hz -0.0196375 0.000129693
+ 2.691e+11Hz -0.0196334 0.000140086
+ 2.692e+11Hz -0.0196292 0.000150694
+ 2.693e+11Hz -0.019625 0.000161518
+ 2.694e+11Hz -0.0196208 0.000172559
+ 2.695e+11Hz -0.0196166 0.000183818
+ 2.696e+11Hz -0.0196123 0.000195295
+ 2.697e+11Hz -0.019608 0.000206992
+ 2.698e+11Hz -0.0196036 0.000218907
+ 2.699e+11Hz -0.0195992 0.000231043
+ 2.7e+11Hz -0.0195947 0.000243399
+ 2.701e+11Hz -0.0195901 0.000255975
+ 2.702e+11Hz -0.0195855 0.000268773
+ 2.703e+11Hz -0.0195808 0.000281792
+ 2.704e+11Hz -0.0195761 0.000295032
+ 2.705e+11Hz -0.0195713 0.000308494
+ 2.706e+11Hz -0.0195664 0.000322178
+ 2.707e+11Hz -0.0195614 0.000336083
+ 2.708e+11Hz -0.0195563 0.00035021
+ 2.709e+11Hz -0.0195511 0.000364558
+ 2.71e+11Hz -0.0195459 0.000379128
+ 2.711e+11Hz -0.0195405 0.000393918
+ 2.712e+11Hz -0.0195351 0.00040893
+ 2.713e+11Hz -0.0195295 0.000424161
+ 2.714e+11Hz -0.0195238 0.000439612
+ 2.715e+11Hz -0.019518 0.000455283
+ 2.716e+11Hz -0.0195121 0.000471172
+ 2.717e+11Hz -0.019506 0.000487279
+ 2.718e+11Hz -0.0194999 0.000503603
+ 2.719e+11Hz -0.0194936 0.000520144
+ 2.72e+11Hz -0.0194871 0.000536899
+ 2.721e+11Hz -0.0194805 0.00055387
+ 2.722e+11Hz -0.0194738 0.000571054
+ 2.723e+11Hz -0.0194669 0.000588449
+ 2.724e+11Hz -0.0194599 0.000606056
+ 2.725e+11Hz -0.0194527 0.000623873
+ 2.726e+11Hz -0.0194453 0.000641898
+ 2.727e+11Hz -0.0194378 0.00066013
+ 2.728e+11Hz -0.01943 0.000678567
+ 2.729e+11Hz -0.0194222 0.000697208
+ 2.73e+11Hz -0.0194141 0.00071605
+ 2.731e+11Hz -0.0194058 0.000735093
+ 2.732e+11Hz -0.0193974 0.000754334
+ 2.733e+11Hz -0.0193888 0.000773772
+ 2.734e+11Hz -0.0193799 0.000793404
+ 2.735e+11Hz -0.0193709 0.000813228
+ 2.736e+11Hz -0.0193616 0.000833242
+ 2.737e+11Hz -0.0193522 0.000853444
+ 2.738e+11Hz -0.0193425 0.000873831
+ 2.739e+11Hz -0.0193326 0.000894401
+ 2.74e+11Hz -0.0193225 0.000915151
+ 2.741e+11Hz -0.0193121 0.000936079
+ 2.742e+11Hz -0.0193016 0.000957182
+ 2.743e+11Hz -0.0192907 0.000978457
+ 2.744e+11Hz -0.0192797 0.000999901
+ 2.745e+11Hz -0.0192684 0.00102151
+ 2.746e+11Hz -0.0192568 0.00104328
+ 2.747e+11Hz -0.019245 0.00106522
+ 2.748e+11Hz -0.0192329 0.00108731
+ 2.749e+11Hz -0.0192206 0.00110955
+ 2.75e+11Hz -0.019208 0.00113195
+ 2.751e+11Hz -0.0191951 0.00115449
+ 2.752e+11Hz -0.019182 0.00117717
+ 2.753e+11Hz -0.0191686 0.0012
+ 2.754e+11Hz -0.0191549 0.00122295
+ 2.755e+11Hz -0.0191409 0.00124604
+ 2.756e+11Hz -0.0191266 0.00126926
+ 2.757e+11Hz -0.0191121 0.00129261
+ 2.758e+11Hz -0.0190972 0.00131607
+ 2.759e+11Hz -0.0190821 0.00133965
+ 2.76e+11Hz -0.0190666 0.00136333
+ 2.761e+11Hz -0.0190509 0.00138713
+ 2.762e+11Hz -0.0190348 0.00141103
+ 2.763e+11Hz -0.0190184 0.00143503
+ 2.764e+11Hz -0.0190017 0.00145912
+ 2.765e+11Hz -0.0189847 0.0014833
+ 2.766e+11Hz -0.0189674 0.00150756
+ 2.767e+11Hz -0.0189497 0.00153191
+ 2.768e+11Hz -0.0189317 0.00155633
+ 2.769e+11Hz -0.0189134 0.00158082
+ 2.77e+11Hz -0.0188947 0.00160537
+ 2.771e+11Hz -0.0188757 0.00162998
+ 2.772e+11Hz -0.0188564 0.00165465
+ 2.773e+11Hz -0.0188367 0.00167937
+ 2.774e+11Hz -0.0188167 0.00170413
+ 2.775e+11Hz -0.0187964 0.00172893
+ 2.776e+11Hz -0.0187757 0.00175376
+ 2.777e+11Hz -0.0187546 0.00177862
+ 2.778e+11Hz -0.0187332 0.00180351
+ 2.779e+11Hz -0.0187114 0.00182841
+ 2.78e+11Hz -0.0186893 0.00185332
+ 2.781e+11Hz -0.0186668 0.00187824
+ 2.782e+11Hz -0.018644 0.00190316
+ 2.783e+11Hz -0.0186208 0.00192807
+ 2.784e+11Hz -0.0185972 0.00195297
+ 2.785e+11Hz -0.0185733 0.00197785
+ 2.786e+11Hz -0.018549 0.00200271
+ 2.787e+11Hz -0.0185243 0.00202753
+ 2.788e+11Hz -0.0184993 0.00205232
+ 2.789e+11Hz -0.0184739 0.00207707
+ 2.79e+11Hz -0.0184482 0.00210178
+ 2.791e+11Hz -0.018422 0.00212642
+ 2.792e+11Hz -0.0183955 0.00215101
+ 2.793e+11Hz -0.0183686 0.00217553
+ 2.794e+11Hz -0.0183414 0.00219998
+ 2.795e+11Hz -0.0183137 0.00222435
+ 2.796e+11Hz -0.0182857 0.00224863
+ 2.797e+11Hz -0.0182574 0.00227282
+ 2.798e+11Hz -0.0182286 0.00229692
+ 2.799e+11Hz -0.0181995 0.0023209
+ 2.8e+11Hz -0.01817 0.00234478
+ 2.801e+11Hz -0.0181401 0.00236854
+ 2.802e+11Hz -0.0181099 0.00239218
+ 2.803e+11Hz -0.0180793 0.00241568
+ 2.804e+11Hz -0.0180483 0.00243905
+ 2.805e+11Hz -0.018017 0.00246227
+ 2.806e+11Hz -0.0179852 0.00248535
+ 2.807e+11Hz -0.0179531 0.00250826
+ 2.808e+11Hz -0.0179207 0.00253102
+ 2.809e+11Hz -0.0178879 0.00255361
+ 2.81e+11Hz -0.0178547 0.00257602
+ 2.811e+11Hz -0.0178211 0.00259824
+ 2.812e+11Hz -0.0177872 0.00262028
+ 2.813e+11Hz -0.017753 0.00264213
+ 2.814e+11Hz -0.0177183 0.00266377
+ 2.815e+11Hz -0.0176833 0.0026852
+ 2.816e+11Hz -0.017648 0.00270642
+ 2.817e+11Hz -0.0176123 0.00272742
+ 2.818e+11Hz -0.0175763 0.00274819
+ 2.819e+11Hz -0.0175399 0.00276873
+ 2.82e+11Hz -0.0175032 0.00278903
+ 2.821e+11Hz -0.0174661 0.00280908
+ 2.822e+11Hz -0.0174287 0.00282888
+ 2.823e+11Hz -0.017391 0.00284842
+ 2.824e+11Hz -0.0173529 0.00286769
+ 2.825e+11Hz -0.0173146 0.0028867
+ 2.826e+11Hz -0.0172758 0.00290543
+ 2.827e+11Hz -0.0172368 0.00292387
+ 2.828e+11Hz -0.0171975 0.00294203
+ 2.829e+11Hz -0.0171578 0.00295989
+ 2.83e+11Hz -0.0171178 0.00297745
+ 2.831e+11Hz -0.0170775 0.00299471
+ 2.832e+11Hz -0.0170369 0.00301165
+ 2.833e+11Hz -0.0169961 0.00302828
+ 2.834e+11Hz -0.0169549 0.00304458
+ 2.835e+11Hz -0.0169134 0.00306056
+ 2.836e+11Hz -0.0168717 0.0030762
+ 2.837e+11Hz -0.0168297 0.0030915
+ 2.838e+11Hz -0.0167874 0.00310645
+ 2.839e+11Hz -0.0167448 0.00312106
+ 2.84e+11Hz -0.016702 0.00313531
+ 2.841e+11Hz -0.0166589 0.0031492
+ 2.842e+11Hz -0.0166156 0.00316272
+ 2.843e+11Hz -0.016572 0.00317587
+ 2.844e+11Hz -0.0165281 0.00318865
+ 2.845e+11Hz -0.0164841 0.00320105
+ 2.846e+11Hz -0.0164398 0.00321307
+ 2.847e+11Hz -0.0163952 0.0032247
+ 2.848e+11Hz -0.0163505 0.00323593
+ 2.849e+11Hz -0.0163055 0.00324677
+ 2.85e+11Hz -0.0162604 0.0032572
+ 2.851e+11Hz -0.016215 0.00326723
+ 2.852e+11Hz -0.0161694 0.00327685
+ 2.853e+11Hz -0.0161237 0.00328606
+ 2.854e+11Hz -0.0160777 0.00329485
+ 2.855e+11Hz -0.0160316 0.00330322
+ 2.856e+11Hz -0.0159853 0.00331116
+ 2.857e+11Hz -0.0159389 0.00331868
+ 2.858e+11Hz -0.0158923 0.00332577
+ 2.859e+11Hz -0.0158455 0.00333242
+ 2.86e+11Hz -0.0157986 0.00333863
+ 2.861e+11Hz -0.0157516 0.00334441
+ 2.862e+11Hz -0.0157044 0.00334974
+ 2.863e+11Hz -0.0156571 0.00335463
+ 2.864e+11Hz -0.0156097 0.00335906
+ 2.865e+11Hz -0.0155622 0.00336305
+ 2.866e+11Hz -0.0155146 0.00336659
+ 2.867e+11Hz -0.0154669 0.00336967
+ 2.868e+11Hz -0.0154191 0.00337229
+ 2.869e+11Hz -0.0153712 0.00337446
+ 2.87e+11Hz -0.0153233 0.00337616
+ 2.871e+11Hz -0.0152753 0.00337741
+ 2.872e+11Hz -0.0152272 0.00337819
+ 2.873e+11Hz -0.0151791 0.0033785
+ 2.874e+11Hz -0.0151309 0.00337835
+ 2.875e+11Hz -0.0150827 0.00337774
+ 2.876e+11Hz -0.0150345 0.00337665
+ 2.877e+11Hz -0.0149863 0.0033751
+ 2.878e+11Hz -0.014938 0.00337308
+ 2.879e+11Hz -0.0148898 0.00337059
+ 2.88e+11Hz -0.0148415 0.00336763
+ 2.881e+11Hz -0.0147933 0.0033642
+ 2.882e+11Hz -0.0147451 0.0033603
+ 2.883e+11Hz -0.0146969 0.00335593
+ 2.884e+11Hz -0.0146487 0.00335109
+ 2.885e+11Hz -0.0146006 0.00334578
+ 2.886e+11Hz -0.0145525 0.00334001
+ 2.887e+11Hz -0.0145045 0.00333376
+ 2.888e+11Hz -0.0144566 0.00332705
+ 2.889e+11Hz -0.0144087 0.00331988
+ 2.89e+11Hz -0.0143609 0.00331224
+ 2.891e+11Hz -0.0143132 0.00330414
+ 2.892e+11Hz -0.0142656 0.00329557
+ 2.893e+11Hz -0.0142181 0.00328655
+ 2.894e+11Hz -0.0141707 0.00327707
+ 2.895e+11Hz -0.0141234 0.00326713
+ 2.896e+11Hz -0.0140763 0.00325674
+ 2.897e+11Hz -0.0140293 0.0032459
+ 2.898e+11Hz -0.0139824 0.00323461
+ 2.899e+11Hz -0.0139357 0.00322287
+ 2.9e+11Hz -0.0138891 0.00321068
+ 2.901e+11Hz -0.0138427 0.00319805
+ 2.902e+11Hz -0.0137964 0.00318499
+ 2.903e+11Hz -0.0137504 0.00317149
+ 2.904e+11Hz -0.0137045 0.00315756
+ 2.905e+11Hz -0.0136588 0.0031432
+ 2.906e+11Hz -0.0136133 0.00312841
+ 2.907e+11Hz -0.013568 0.0031132
+ 2.908e+11Hz -0.0135229 0.00309757
+ 2.909e+11Hz -0.013478 0.00308153
+ 2.91e+11Hz -0.0134334 0.00306507
+ 2.911e+11Hz -0.013389 0.00304821
+ 2.912e+11Hz -0.0133448 0.00303095
+ 2.913e+11Hz -0.0133009 0.00301329
+ 2.914e+11Hz -0.0132572 0.00299524
+ 2.915e+11Hz -0.0132138 0.0029768
+ 2.916e+11Hz -0.0131706 0.00295797
+ 2.917e+11Hz -0.0131277 0.00293877
+ 2.918e+11Hz -0.0130851 0.00291919
+ 2.919e+11Hz -0.0130427 0.00289924
+ 2.92e+11Hz -0.0130007 0.00287893
+ 2.921e+11Hz -0.0129589 0.00285826
+ 2.922e+11Hz -0.0129174 0.00283723
+ 2.923e+11Hz -0.0128763 0.00281586
+ 2.924e+11Hz -0.0128354 0.00279415
+ 2.925e+11Hz -0.0127949 0.0027721
+ 2.926e+11Hz -0.0127546 0.00274972
+ 2.927e+11Hz -0.0127147 0.00272701
+ 2.928e+11Hz -0.0126751 0.00270398
+ 2.929e+11Hz -0.0126359 0.00268065
+ 2.93e+11Hz -0.012597 0.002657
+ 2.931e+11Hz -0.0125584 0.00263305
+ 2.932e+11Hz -0.0125202 0.00260882
+ 2.933e+11Hz -0.0124823 0.00258429
+ 2.934e+11Hz -0.0124448 0.00255948
+ 2.935e+11Hz -0.0124076 0.0025344
+ 2.936e+11Hz -0.0123708 0.00250904
+ 2.937e+11Hz -0.0123344 0.00248343
+ 2.938e+11Hz -0.0122983 0.00245756
+ 2.939e+11Hz -0.0122626 0.00243145
+ 2.94e+11Hz -0.0122273 0.00240509
+ 2.941e+11Hz -0.0121923 0.0023785
+ 2.942e+11Hz -0.0121578 0.00235168
+ 2.943e+11Hz -0.0121236 0.00232464
+ 2.944e+11Hz -0.0120898 0.00229738
+ 2.945e+11Hz -0.0120564 0.00226993
+ 2.946e+11Hz -0.0120234 0.00224227
+ 2.947e+11Hz -0.0119908 0.00221442
+ 2.948e+11Hz -0.0119585 0.00218638
+ 2.949e+11Hz -0.0119267 0.00215817
+ 2.95e+11Hz -0.0118953 0.00212979
+ 2.951e+11Hz -0.0118642 0.00210124
+ 2.952e+11Hz -0.0118336 0.00207254
+ 2.953e+11Hz -0.0118034 0.00204369
+ 2.954e+11Hz -0.0117736 0.0020147
+ 2.955e+11Hz -0.0117442 0.00198558
+ 2.956e+11Hz -0.0117152 0.00195633
+ 2.957e+11Hz -0.0116866 0.00192696
+ 2.958e+11Hz -0.0116584 0.00189747
+ 2.959e+11Hz -0.0116306 0.00186789
+ 2.96e+11Hz -0.0116033 0.0018382
+ 2.961e+11Hz -0.0115763 0.00180843
+ 2.962e+11Hz -0.0115498 0.00177858
+ 2.963e+11Hz -0.0115237 0.00174865
+ 2.964e+11Hz -0.0114979 0.00171865
+ 2.965e+11Hz -0.0114726 0.00168859
+ 2.966e+11Hz -0.0114477 0.00165848
+ 2.967e+11Hz -0.0114232 0.00162832
+ 2.968e+11Hz -0.0113991 0.00159812
+ 2.969e+11Hz -0.0113754 0.00156789
+ 2.97e+11Hz -0.0113522 0.00153764
+ 2.971e+11Hz -0.0113293 0.00150737
+ 2.972e+11Hz -0.0113068 0.00147708
+ 2.973e+11Hz -0.0112848 0.0014468
+ 2.974e+11Hz -0.0112631 0.00141651
+ 2.975e+11Hz -0.0112418 0.00138624
+ 2.976e+11Hz -0.0112209 0.00135598
+ 2.977e+11Hz -0.0112004 0.00132575
+ 2.978e+11Hz -0.0111804 0.00129555
+ 2.979e+11Hz -0.0111607 0.00126538
+ 2.98e+11Hz -0.0111413 0.00123526
+ 2.981e+11Hz -0.0111224 0.00120519
+ 2.982e+11Hz -0.0111039 0.00117517
+ 2.983e+11Hz -0.0110857 0.00114522
+ 2.984e+11Hz -0.0110679 0.00111534
+ 2.985e+11Hz -0.0110505 0.00108553
+ 2.986e+11Hz -0.0110334 0.0010558
+ 2.987e+11Hz -0.0110167 0.00102616
+ 2.988e+11Hz -0.0110004 0.000996611
+ 2.989e+11Hz -0.0109844 0.000967163
+ 2.99e+11Hz -0.0109688 0.000937819
+ 2.991e+11Hz -0.0109536 0.000908586
+ 2.992e+11Hz -0.0109387 0.000879469
+ 2.993e+11Hz -0.0109241 0.000850473
+ 2.994e+11Hz -0.0109099 0.000821604
+ 2.995e+11Hz -0.010896 0.000792867
+ 2.996e+11Hz -0.0108824 0.000764267
+ 2.997e+11Hz -0.0108692 0.00073581
+ 2.998e+11Hz -0.0108563 0.000707499
+ 2.999e+11Hz -0.0108437 0.000679341
+ 3e+11Hz -0.0108314 0.00065134
+ ]

A12 %vd(20 3) %vd(12, 3) xfer2
.model xfer2 xfer R_I=true table=[
+ 0Hz 0.995436 0
+ 1e+08Hz 0.995435 -0.000814178
+ 2e+08Hz 0.995433 -0.00162834
+ 3e+08Hz 0.99543 -0.00244247
+ 4e+08Hz 0.995425 -0.00325656
+ 5e+08Hz 0.99542 -0.00407058
+ 6e+08Hz 0.995412 -0.00488452
+ 7e+08Hz 0.995404 -0.00569837
+ 8e+08Hz 0.995394 -0.00651211
+ 9e+08Hz 0.995383 -0.00732573
+ 1e+09Hz 0.995371 -0.0081392
+ 1.1e+09Hz 0.995358 -0.00895252
+ 1.2e+09Hz 0.995343 -0.00976567
+ 1.3e+09Hz 0.995327 -0.0105786
+ 1.4e+09Hz 0.99531 -0.0113914
+ 1.5e+09Hz 0.995291 -0.012204
+ 1.6e+09Hz 0.995271 -0.0130163
+ 1.7e+09Hz 0.99525 -0.0138284
+ 1.8e+09Hz 0.995228 -0.0146402
+ 1.9e+09Hz 0.995204 -0.0154517
+ 2e+09Hz 0.99518 -0.016263
+ 2.1e+09Hz 0.995154 -0.017074
+ 2.2e+09Hz 0.995126 -0.0178846
+ 2.3e+09Hz 0.995098 -0.0186949
+ 2.4e+09Hz 0.995068 -0.0195049
+ 2.5e+09Hz 0.995038 -0.0203146
+ 2.6e+09Hz 0.995006 -0.0211238
+ 2.7e+09Hz 0.994973 -0.0219327
+ 2.8e+09Hz 0.994938 -0.0227412
+ 2.9e+09Hz 0.994903 -0.0235493
+ 3e+09Hz 0.994866 -0.024357
+ 3.1e+09Hz 0.994829 -0.0251643
+ 3.2e+09Hz 0.99479 -0.0259711
+ 3.3e+09Hz 0.99475 -0.0267775
+ 3.4e+09Hz 0.994709 -0.0275834
+ 3.5e+09Hz 0.994667 -0.0283889
+ 3.6e+09Hz 0.994624 -0.0291939
+ 3.7e+09Hz 0.994579 -0.0299984
+ 3.8e+09Hz 0.994534 -0.0308024
+ 3.9e+09Hz 0.994488 -0.031606
+ 4e+09Hz 0.994441 -0.032409
+ 4.1e+09Hz 0.994392 -0.0332114
+ 4.2e+09Hz 0.994343 -0.0340134
+ 4.3e+09Hz 0.994292 -0.0348148
+ 4.4e+09Hz 0.994241 -0.0356157
+ 4.5e+09Hz 0.994189 -0.036416
+ 4.6e+09Hz 0.994136 -0.0372158
+ 4.7e+09Hz 0.994081 -0.038015
+ 4.8e+09Hz 0.994026 -0.0388137
+ 4.9e+09Hz 0.99397 -0.0396118
+ 5e+09Hz 0.993913 -0.0404093
+ 5.1e+09Hz 0.993856 -0.0412062
+ 5.2e+09Hz 0.993797 -0.0420026
+ 5.3e+09Hz 0.993737 -0.0427983
+ 5.4e+09Hz 0.993677 -0.0435935
+ 5.5e+09Hz 0.993616 -0.044388
+ 5.6e+09Hz 0.993554 -0.045182
+ 5.7e+09Hz 0.993491 -0.0459753
+ 5.8e+09Hz 0.993427 -0.0467681
+ 5.9e+09Hz 0.993363 -0.0475602
+ 6e+09Hz 0.993298 -0.0483518
+ 6.1e+09Hz 0.993232 -0.0491427
+ 6.2e+09Hz 0.993165 -0.049933
+ 6.3e+09Hz 0.993098 -0.0507227
+ 6.4e+09Hz 0.99303 -0.0515118
+ 6.5e+09Hz 0.992961 -0.0523003
+ 6.6e+09Hz 0.992892 -0.0530882
+ 6.7e+09Hz 0.992821 -0.0538755
+ 6.8e+09Hz 0.992751 -0.0546622
+ 6.9e+09Hz 0.992679 -0.0554482
+ 7e+09Hz 0.992607 -0.0562337
+ 7.1e+09Hz 0.992535 -0.0570185
+ 7.2e+09Hz 0.992461 -0.0578028
+ 7.3e+09Hz 0.992387 -0.0585865
+ 7.4e+09Hz 0.992313 -0.0593695
+ 7.5e+09Hz 0.992238 -0.060152
+ 7.6e+09Hz 0.992162 -0.0609339
+ 7.7e+09Hz 0.992086 -0.0617152
+ 7.8e+09Hz 0.99201 -0.062496
+ 7.9e+09Hz 0.991933 -0.0632762
+ 8e+09Hz 0.991855 -0.0640558
+ 8.1e+09Hz 0.991777 -0.0648348
+ 8.2e+09Hz 0.991698 -0.0656133
+ 8.3e+09Hz 0.991619 -0.0663912
+ 8.4e+09Hz 0.99154 -0.0671686
+ 8.5e+09Hz 0.991459 -0.0679455
+ 8.6e+09Hz 0.991379 -0.0687218
+ 8.7e+09Hz 0.991298 -0.0694976
+ 8.8e+09Hz 0.991217 -0.0702728
+ 8.9e+09Hz 0.991135 -0.0710476
+ 9e+09Hz 0.991053 -0.0718218
+ 9.1e+09Hz 0.99097 -0.0725956
+ 9.2e+09Hz 0.990888 -0.0733689
+ 9.3e+09Hz 0.990804 -0.0741417
+ 9.4e+09Hz 0.990721 -0.074914
+ 9.5e+09Hz 0.990637 -0.0756858
+ 9.6e+09Hz 0.990552 -0.0764572
+ 9.7e+09Hz 0.990467 -0.0772282
+ 9.8e+09Hz 0.990382 -0.0779987
+ 9.9e+09Hz 0.990297 -0.0787687
+ 1e+10Hz 0.990211 -0.0795384
+ 1.01e+10Hz 0.990125 -0.0803076
+ 1.02e+10Hz 0.990039 -0.0810764
+ 1.03e+10Hz 0.989952 -0.0818449
+ 1.04e+10Hz 0.989865 -0.0826129
+ 1.05e+10Hz 0.989778 -0.0833806
+ 1.06e+10Hz 0.98969 -0.0841479
+ 1.07e+10Hz 0.989603 -0.0849148
+ 1.08e+10Hz 0.989514 -0.0856814
+ 1.09e+10Hz 0.989426 -0.0864477
+ 1.1e+10Hz 0.989337 -0.0872136
+ 1.11e+10Hz 0.989248 -0.0879793
+ 1.12e+10Hz 0.989159 -0.0887446
+ 1.13e+10Hz 0.98907 -0.0895096
+ 1.14e+10Hz 0.98898 -0.0902743
+ 1.15e+10Hz 0.98889 -0.0910387
+ 1.16e+10Hz 0.9888 -0.0918029
+ 1.17e+10Hz 0.988709 -0.0925668
+ 1.18e+10Hz 0.988618 -0.0933304
+ 1.19e+10Hz 0.988527 -0.0940938
+ 1.2e+10Hz 0.988436 -0.094857
+ 1.21e+10Hz 0.988344 -0.09562
+ 1.22e+10Hz 0.988253 -0.0963827
+ 1.23e+10Hz 0.988161 -0.0971453
+ 1.24e+10Hz 0.988068 -0.0979076
+ 1.25e+10Hz 0.987976 -0.0986698
+ 1.26e+10Hz 0.987883 -0.0994318
+ 1.27e+10Hz 0.98779 -0.100194
+ 1.28e+10Hz 0.987697 -0.100955
+ 1.29e+10Hz 0.987603 -0.101717
+ 1.3e+10Hz 0.987509 -0.102478
+ 1.31e+10Hz 0.987415 -0.10324
+ 1.32e+10Hz 0.987321 -0.104001
+ 1.33e+10Hz 0.987226 -0.104762
+ 1.34e+10Hz 0.987131 -0.105523
+ 1.35e+10Hz 0.987036 -0.106283
+ 1.36e+10Hz 0.986941 -0.107044
+ 1.37e+10Hz 0.986845 -0.107805
+ 1.38e+10Hz 0.986749 -0.108566
+ 1.39e+10Hz 0.986653 -0.109326
+ 1.4e+10Hz 0.986556 -0.110087
+ 1.41e+10Hz 0.986459 -0.110847
+ 1.42e+10Hz 0.986362 -0.111607
+ 1.43e+10Hz 0.986265 -0.112368
+ 1.44e+10Hz 0.986167 -0.113128
+ 1.45e+10Hz 0.986069 -0.113888
+ 1.46e+10Hz 0.985971 -0.114649
+ 1.47e+10Hz 0.985872 -0.115409
+ 1.48e+10Hz 0.985773 -0.116169
+ 1.49e+10Hz 0.985673 -0.11693
+ 1.5e+10Hz 0.985574 -0.11769
+ 1.51e+10Hz 0.985474 -0.11845
+ 1.52e+10Hz 0.985373 -0.119211
+ 1.53e+10Hz 0.985273 -0.119971
+ 1.54e+10Hz 0.985172 -0.120732
+ 1.55e+10Hz 0.98507 -0.121492
+ 1.56e+10Hz 0.984968 -0.122253
+ 1.57e+10Hz 0.984866 -0.123013
+ 1.58e+10Hz 0.984763 -0.123774
+ 1.59e+10Hz 0.98466 -0.124535
+ 1.6e+10Hz 0.984557 -0.125295
+ 1.61e+10Hz 0.984453 -0.126056
+ 1.62e+10Hz 0.984349 -0.126817
+ 1.63e+10Hz 0.984244 -0.127578
+ 1.64e+10Hz 0.984139 -0.128339
+ 1.65e+10Hz 0.984034 -0.1291
+ 1.66e+10Hz 0.983928 -0.129861
+ 1.67e+10Hz 0.983822 -0.130623
+ 1.68e+10Hz 0.983715 -0.131384
+ 1.69e+10Hz 0.983607 -0.132145
+ 1.7e+10Hz 0.9835 -0.132907
+ 1.71e+10Hz 0.983391 -0.133669
+ 1.72e+10Hz 0.983283 -0.13443
+ 1.73e+10Hz 0.983174 -0.135192
+ 1.74e+10Hz 0.983064 -0.135954
+ 1.75e+10Hz 0.982954 -0.136716
+ 1.76e+10Hz 0.982843 -0.137478
+ 1.77e+10Hz 0.982732 -0.13824
+ 1.78e+10Hz 0.98262 -0.139002
+ 1.79e+10Hz 0.982508 -0.139765
+ 1.8e+10Hz 0.982395 -0.140527
+ 1.81e+10Hz 0.982281 -0.14129
+ 1.82e+10Hz 0.982167 -0.142052
+ 1.83e+10Hz 0.982053 -0.142815
+ 1.84e+10Hz 0.981938 -0.143578
+ 1.85e+10Hz 0.981822 -0.14434
+ 1.86e+10Hz 0.981706 -0.145103
+ 1.87e+10Hz 0.981589 -0.145866
+ 1.88e+10Hz 0.981472 -0.146629
+ 1.89e+10Hz 0.981354 -0.147393
+ 1.9e+10Hz 0.981235 -0.148156
+ 1.91e+10Hz 0.981116 -0.148919
+ 1.92e+10Hz 0.980996 -0.149682
+ 1.93e+10Hz 0.980876 -0.150446
+ 1.94e+10Hz 0.980754 -0.151209
+ 1.95e+10Hz 0.980633 -0.151973
+ 1.96e+10Hz 0.98051 -0.152736
+ 1.97e+10Hz 0.980387 -0.1535
+ 1.98e+10Hz 0.980264 -0.154264
+ 1.99e+10Hz 0.980139 -0.155027
+ 2e+10Hz 0.980014 -0.155791
+ 2.01e+10Hz 0.979889 -0.156555
+ 2.02e+10Hz 0.979762 -0.157319
+ 2.03e+10Hz 0.979635 -0.158083
+ 2.04e+10Hz 0.979508 -0.158846
+ 2.05e+10Hz 0.979379 -0.15961
+ 2.06e+10Hz 0.97925 -0.160374
+ 2.07e+10Hz 0.979121 -0.161138
+ 2.08e+10Hz 0.97899 -0.161902
+ 2.09e+10Hz 0.978859 -0.162666
+ 2.1e+10Hz 0.978727 -0.16343
+ 2.11e+10Hz 0.978595 -0.164193
+ 2.12e+10Hz 0.978461 -0.164957
+ 2.13e+10Hz 0.978327 -0.165721
+ 2.14e+10Hz 0.978193 -0.166485
+ 2.15e+10Hz 0.978057 -0.167249
+ 2.16e+10Hz 0.977921 -0.168012
+ 2.17e+10Hz 0.977785 -0.168776
+ 2.18e+10Hz 0.977647 -0.169539
+ 2.19e+10Hz 0.977509 -0.170303
+ 2.2e+10Hz 0.97737 -0.171066
+ 2.21e+10Hz 0.97723 -0.17183
+ 2.22e+10Hz 0.97709 -0.172593
+ 2.23e+10Hz 0.976948 -0.173356
+ 2.24e+10Hz 0.976807 -0.174119
+ 2.25e+10Hz 0.976664 -0.174882
+ 2.26e+10Hz 0.976521 -0.175645
+ 2.27e+10Hz 0.976377 -0.176408
+ 2.28e+10Hz 0.976232 -0.17717
+ 2.29e+10Hz 0.976086 -0.177933
+ 2.3e+10Hz 0.97594 -0.178695
+ 2.31e+10Hz 0.975793 -0.179458
+ 2.32e+10Hz 0.975645 -0.18022
+ 2.33e+10Hz 0.975497 -0.180982
+ 2.34e+10Hz 0.975348 -0.181743
+ 2.35e+10Hz 0.975198 -0.182505
+ 2.36e+10Hz 0.975047 -0.183267
+ 2.37e+10Hz 0.974896 -0.184028
+ 2.38e+10Hz 0.974744 -0.184789
+ 2.39e+10Hz 0.974591 -0.18555
+ 2.4e+10Hz 0.974438 -0.186311
+ 2.41e+10Hz 0.974284 -0.187072
+ 2.42e+10Hz 0.974129 -0.187832
+ 2.43e+10Hz 0.973973 -0.188592
+ 2.44e+10Hz 0.973817 -0.189352
+ 2.45e+10Hz 0.97366 -0.190112
+ 2.46e+10Hz 0.973502 -0.190872
+ 2.47e+10Hz 0.973344 -0.191631
+ 2.48e+10Hz 0.973185 -0.19239
+ 2.49e+10Hz 0.973025 -0.193149
+ 2.5e+10Hz 0.972864 -0.193908
+ 2.51e+10Hz 0.972703 -0.194667
+ 2.52e+10Hz 0.972541 -0.195425
+ 2.53e+10Hz 0.972379 -0.196183
+ 2.54e+10Hz 0.972216 -0.196941
+ 2.55e+10Hz 0.972052 -0.197698
+ 2.56e+10Hz 0.971887 -0.198455
+ 2.57e+10Hz 0.971722 -0.199212
+ 2.58e+10Hz 0.971556 -0.199969
+ 2.59e+10Hz 0.97139 -0.200726
+ 2.6e+10Hz 0.971223 -0.201482
+ 2.61e+10Hz 0.971055 -0.202238
+ 2.62e+10Hz 0.970886 -0.202994
+ 2.63e+10Hz 0.970717 -0.203749
+ 2.64e+10Hz 0.970548 -0.204504
+ 2.65e+10Hz 0.970377 -0.205259
+ 2.66e+10Hz 0.970206 -0.206014
+ 2.67e+10Hz 0.970035 -0.206768
+ 2.68e+10Hz 0.969863 -0.207522
+ 2.69e+10Hz 0.96969 -0.208276
+ 2.7e+10Hz 0.969516 -0.209029
+ 2.71e+10Hz 0.969342 -0.209782
+ 2.72e+10Hz 0.969168 -0.210535
+ 2.73e+10Hz 0.968993 -0.211288
+ 2.74e+10Hz 0.968817 -0.21204
+ 2.75e+10Hz 0.968641 -0.212792
+ 2.76e+10Hz 0.968464 -0.213544
+ 2.77e+10Hz 0.968286 -0.214296
+ 2.78e+10Hz 0.968108 -0.215047
+ 2.79e+10Hz 0.96793 -0.215798
+ 2.8e+10Hz 0.96775 -0.216548
+ 2.81e+10Hz 0.967571 -0.217298
+ 2.82e+10Hz 0.96739 -0.218048
+ 2.83e+10Hz 0.96721 -0.218798
+ 2.84e+10Hz 0.967028 -0.219548
+ 2.85e+10Hz 0.966846 -0.220297
+ 2.86e+10Hz 0.966664 -0.221046
+ 2.87e+10Hz 0.966481 -0.221794
+ 2.88e+10Hz 0.966298 -0.222542
+ 2.89e+10Hz 0.966114 -0.22329
+ 2.9e+10Hz 0.965929 -0.224038
+ 2.91e+10Hz 0.965744 -0.224785
+ 2.92e+10Hz 0.965559 -0.225533
+ 2.93e+10Hz 0.965373 -0.22628
+ 2.94e+10Hz 0.965186 -0.227026
+ 2.95e+10Hz 0.964999 -0.227772
+ 2.96e+10Hz 0.964812 -0.228519
+ 2.97e+10Hz 0.964624 -0.229264
+ 2.98e+10Hz 0.964435 -0.23001
+ 2.99e+10Hz 0.964246 -0.230755
+ 3e+10Hz 0.964057 -0.2315
+ 3.01e+10Hz 0.963867 -0.232245
+ 3.02e+10Hz 0.963677 -0.232989
+ 3.03e+10Hz 0.963486 -0.233734
+ 3.04e+10Hz 0.963295 -0.234478
+ 3.05e+10Hz 0.963103 -0.235221
+ 3.06e+10Hz 0.962911 -0.235965
+ 3.07e+10Hz 0.962718 -0.236708
+ 3.08e+10Hz 0.962525 -0.237451
+ 3.09e+10Hz 0.962332 -0.238194
+ 3.1e+10Hz 0.962138 -0.238936
+ 3.11e+10Hz 0.961943 -0.239679
+ 3.12e+10Hz 0.961748 -0.240421
+ 3.13e+10Hz 0.961553 -0.241163
+ 3.14e+10Hz 0.961357 -0.241905
+ 3.15e+10Hz 0.961161 -0.242646
+ 3.16e+10Hz 0.960964 -0.243387
+ 3.17e+10Hz 0.960767 -0.244128
+ 3.18e+10Hz 0.96057 -0.244869
+ 3.19e+10Hz 0.960372 -0.24561
+ 3.2e+10Hz 0.960174 -0.24635
+ 3.21e+10Hz 0.959975 -0.247091
+ 3.22e+10Hz 0.959775 -0.247831
+ 3.23e+10Hz 0.959576 -0.248571
+ 3.24e+10Hz 0.959376 -0.24931
+ 3.25e+10Hz 0.959175 -0.25005
+ 3.26e+10Hz 0.958974 -0.250789
+ 3.27e+10Hz 0.958773 -0.251528
+ 3.28e+10Hz 0.958571 -0.252267
+ 3.29e+10Hz 0.958369 -0.253006
+ 3.3e+10Hz 0.958166 -0.253745
+ 3.31e+10Hz 0.957963 -0.254484
+ 3.32e+10Hz 0.95776 -0.255222
+ 3.33e+10Hz 0.957556 -0.25596
+ 3.34e+10Hz 0.957351 -0.256698
+ 3.35e+10Hz 0.957146 -0.257436
+ 3.36e+10Hz 0.956941 -0.258174
+ 3.37e+10Hz 0.956735 -0.258912
+ 3.38e+10Hz 0.956529 -0.25965
+ 3.39e+10Hz 0.956323 -0.260387
+ 3.4e+10Hz 0.956116 -0.261125
+ 3.41e+10Hz 0.955908 -0.261862
+ 3.42e+10Hz 0.9557 -0.262599
+ 3.43e+10Hz 0.955492 -0.263336
+ 3.44e+10Hz 0.955283 -0.264073
+ 3.45e+10Hz 0.955074 -0.26481
+ 3.46e+10Hz 0.954864 -0.265546
+ 3.47e+10Hz 0.954654 -0.266283
+ 3.48e+10Hz 0.954443 -0.26702
+ 3.49e+10Hz 0.954232 -0.267756
+ 3.5e+10Hz 0.954021 -0.268492
+ 3.51e+10Hz 0.953809 -0.269228
+ 3.52e+10Hz 0.953596 -0.269965
+ 3.53e+10Hz 0.953383 -0.270701
+ 3.54e+10Hz 0.95317 -0.271437
+ 3.55e+10Hz 0.952956 -0.272173
+ 3.56e+10Hz 0.952742 -0.272908
+ 3.57e+10Hz 0.952527 -0.273644
+ 3.58e+10Hz 0.952312 -0.27438
+ 3.59e+10Hz 0.952096 -0.275115
+ 3.6e+10Hz 0.951879 -0.275851
+ 3.61e+10Hz 0.951663 -0.276586
+ 3.62e+10Hz 0.951445 -0.277322
+ 3.63e+10Hz 0.951227 -0.278057
+ 3.64e+10Hz 0.951009 -0.278792
+ 3.65e+10Hz 0.95079 -0.279528
+ 3.66e+10Hz 0.950571 -0.280263
+ 3.67e+10Hz 0.950351 -0.280998
+ 3.68e+10Hz 0.950131 -0.281733
+ 3.69e+10Hz 0.94991 -0.282468
+ 3.7e+10Hz 0.949689 -0.283203
+ 3.71e+10Hz 0.949467 -0.283938
+ 3.72e+10Hz 0.949244 -0.284672
+ 3.73e+10Hz 0.949021 -0.285407
+ 3.74e+10Hz 0.948798 -0.286142
+ 3.75e+10Hz 0.948574 -0.286876
+ 3.76e+10Hz 0.948349 -0.287611
+ 3.77e+10Hz 0.948124 -0.288345
+ 3.78e+10Hz 0.947898 -0.28908
+ 3.79e+10Hz 0.947672 -0.289814
+ 3.8e+10Hz 0.947445 -0.290549
+ 3.81e+10Hz 0.947218 -0.291283
+ 3.82e+10Hz 0.94699 -0.292017
+ 3.83e+10Hz 0.946761 -0.292751
+ 3.84e+10Hz 0.946532 -0.293485
+ 3.85e+10Hz 0.946302 -0.294219
+ 3.86e+10Hz 0.946072 -0.294953
+ 3.87e+10Hz 0.945841 -0.295687
+ 3.88e+10Hz 0.94561 -0.296421
+ 3.89e+10Hz 0.945377 -0.297154
+ 3.9e+10Hz 0.945145 -0.297888
+ 3.91e+10Hz 0.944912 -0.298622
+ 3.92e+10Hz 0.944678 -0.299355
+ 3.93e+10Hz 0.944443 -0.300088
+ 3.94e+10Hz 0.944208 -0.300822
+ 3.95e+10Hz 0.943972 -0.301555
+ 3.96e+10Hz 0.943736 -0.302288
+ 3.97e+10Hz 0.943499 -0.303021
+ 3.98e+10Hz 0.943262 -0.303754
+ 3.99e+10Hz 0.943023 -0.304487
+ 4e+10Hz 0.942785 -0.30522
+ 4.01e+10Hz 0.942545 -0.305953
+ 4.02e+10Hz 0.942305 -0.306685
+ 4.03e+10Hz 0.942065 -0.307418
+ 4.04e+10Hz 0.941823 -0.30815
+ 4.05e+10Hz 0.941581 -0.308882
+ 4.06e+10Hz 0.941339 -0.309615
+ 4.07e+10Hz 0.941095 -0.310347
+ 4.08e+10Hz 0.940851 -0.311079
+ 4.09e+10Hz 0.940607 -0.31181
+ 4.1e+10Hz 0.940362 -0.312542
+ 4.11e+10Hz 0.940116 -0.313274
+ 4.12e+10Hz 0.939869 -0.314005
+ 4.13e+10Hz 0.939622 -0.314736
+ 4.14e+10Hz 0.939374 -0.315468
+ 4.15e+10Hz 0.939126 -0.316199
+ 4.16e+10Hz 0.938877 -0.316929
+ 4.17e+10Hz 0.938627 -0.31766
+ 4.18e+10Hz 0.938377 -0.318391
+ 4.19e+10Hz 0.938126 -0.319121
+ 4.2e+10Hz 0.937874 -0.319851
+ 4.21e+10Hz 0.937621 -0.320581
+ 4.22e+10Hz 0.937368 -0.321311
+ 4.23e+10Hz 0.937114 -0.322041
+ 4.24e+10Hz 0.93686 -0.322771
+ 4.25e+10Hz 0.936605 -0.3235
+ 4.26e+10Hz 0.936349 -0.324229
+ 4.27e+10Hz 0.936093 -0.324958
+ 4.28e+10Hz 0.935836 -0.325687
+ 4.29e+10Hz 0.935578 -0.326416
+ 4.3e+10Hz 0.935319 -0.327144
+ 4.31e+10Hz 0.93506 -0.327872
+ 4.32e+10Hz 0.934801 -0.328601
+ 4.33e+10Hz 0.93454 -0.329328
+ 4.34e+10Hz 0.934279 -0.330056
+ 4.35e+10Hz 0.934017 -0.330783
+ 4.36e+10Hz 0.933755 -0.331511
+ 4.37e+10Hz 0.933492 -0.332238
+ 4.38e+10Hz 0.933228 -0.332964
+ 4.39e+10Hz 0.932964 -0.333691
+ 4.4e+10Hz 0.932698 -0.334417
+ 4.41e+10Hz 0.932433 -0.335143
+ 4.42e+10Hz 0.932166 -0.335869
+ 4.43e+10Hz 0.931899 -0.336594
+ 4.44e+10Hz 0.931632 -0.33732
+ 4.45e+10Hz 0.931363 -0.338045
+ 4.46e+10Hz 0.931094 -0.338769
+ 4.47e+10Hz 0.930825 -0.339494
+ 4.48e+10Hz 0.930554 -0.340218
+ 4.49e+10Hz 0.930283 -0.340942
+ 4.5e+10Hz 0.930012 -0.341666
+ 4.51e+10Hz 0.929739 -0.342389
+ 4.52e+10Hz 0.929467 -0.343113
+ 4.53e+10Hz 0.929193 -0.343836
+ 4.54e+10Hz 0.928919 -0.344558
+ 4.55e+10Hz 0.928644 -0.345281
+ 4.56e+10Hz 0.928369 -0.346003
+ 4.57e+10Hz 0.928093 -0.346724
+ 4.58e+10Hz 0.927816 -0.347446
+ 4.59e+10Hz 0.927539 -0.348167
+ 4.6e+10Hz 0.927261 -0.348888
+ 4.61e+10Hz 0.926982 -0.349609
+ 4.62e+10Hz 0.926703 -0.350329
+ 4.63e+10Hz 0.926423 -0.351049
+ 4.64e+10Hz 0.926143 -0.351769
+ 4.65e+10Hz 0.925862 -0.352488
+ 4.66e+10Hz 0.92558 -0.353207
+ 4.67e+10Hz 0.925298 -0.353926
+ 4.68e+10Hz 0.925015 -0.354644
+ 4.69e+10Hz 0.924732 -0.355362
+ 4.7e+10Hz 0.924448 -0.35608
+ 4.71e+10Hz 0.924163 -0.356798
+ 4.72e+10Hz 0.923878 -0.357515
+ 4.73e+10Hz 0.923592 -0.358232
+ 4.74e+10Hz 0.923306 -0.358949
+ 4.75e+10Hz 0.923019 -0.359665
+ 4.76e+10Hz 0.922732 -0.360381
+ 4.77e+10Hz 0.922444 -0.361096
+ 4.78e+10Hz 0.922155 -0.361812
+ 4.79e+10Hz 0.921866 -0.362527
+ 4.8e+10Hz 0.921576 -0.363241
+ 4.81e+10Hz 0.921286 -0.363955
+ 4.82e+10Hz 0.920995 -0.364669
+ 4.83e+10Hz 0.920704 -0.365383
+ 4.84e+10Hz 0.920412 -0.366096
+ 4.85e+10Hz 0.920119 -0.366809
+ 4.86e+10Hz 0.919826 -0.367522
+ 4.87e+10Hz 0.919532 -0.368234
+ 4.88e+10Hz 0.919238 -0.368946
+ 4.89e+10Hz 0.918944 -0.369658
+ 4.9e+10Hz 0.918649 -0.37037
+ 4.91e+10Hz 0.918353 -0.371081
+ 4.92e+10Hz 0.918057 -0.371791
+ 4.93e+10Hz 0.91776 -0.372502
+ 4.94e+10Hz 0.917463 -0.373212
+ 4.95e+10Hz 0.917165 -0.373922
+ 4.96e+10Hz 0.916866 -0.374631
+ 4.97e+10Hz 0.916568 -0.37534
+ 4.98e+10Hz 0.916268 -0.376049
+ 4.99e+10Hz 0.915969 -0.376757
+ 5e+10Hz 0.915668 -0.377465
+ 5.01e+10Hz 0.915367 -0.378173
+ 5.02e+10Hz 0.915066 -0.378881
+ 5.03e+10Hz 0.914764 -0.379588
+ 5.04e+10Hz 0.914462 -0.380295
+ 5.05e+10Hz 0.914159 -0.381002
+ 5.06e+10Hz 0.913856 -0.381708
+ 5.07e+10Hz 0.913552 -0.382414
+ 5.08e+10Hz 0.913248 -0.383119
+ 5.09e+10Hz 0.912943 -0.383825
+ 5.1e+10Hz 0.912638 -0.38453
+ 5.11e+10Hz 0.912332 -0.385234
+ 5.12e+10Hz 0.912026 -0.385939
+ 5.13e+10Hz 0.91172 -0.386643
+ 5.14e+10Hz 0.911412 -0.387347
+ 5.15e+10Hz 0.911105 -0.38805
+ 5.16e+10Hz 0.910797 -0.388754
+ 5.17e+10Hz 0.910488 -0.389457
+ 5.18e+10Hz 0.910179 -0.390159
+ 5.19e+10Hz 0.90987 -0.390862
+ 5.2e+10Hz 0.90956 -0.391564
+ 5.21e+10Hz 0.90925 -0.392266
+ 5.22e+10Hz 0.908939 -0.392967
+ 5.23e+10Hz 0.908628 -0.393668
+ 5.24e+10Hz 0.908316 -0.394369
+ 5.25e+10Hz 0.908004 -0.39507
+ 5.26e+10Hz 0.907691 -0.395771
+ 5.27e+10Hz 0.907378 -0.396471
+ 5.28e+10Hz 0.907065 -0.397171
+ 5.29e+10Hz 0.906751 -0.39787
+ 5.3e+10Hz 0.906436 -0.39857
+ 5.31e+10Hz 0.906121 -0.399269
+ 5.32e+10Hz 0.905806 -0.399968
+ 5.33e+10Hz 0.90549 -0.400666
+ 5.34e+10Hz 0.905174 -0.401365
+ 5.35e+10Hz 0.904857 -0.402063
+ 5.36e+10Hz 0.90454 -0.402761
+ 5.37e+10Hz 0.904223 -0.403458
+ 5.38e+10Hz 0.903905 -0.404156
+ 5.39e+10Hz 0.903586 -0.404853
+ 5.4e+10Hz 0.903267 -0.40555
+ 5.41e+10Hz 0.902948 -0.406246
+ 5.42e+10Hz 0.902628 -0.406943
+ 5.43e+10Hz 0.902308 -0.407639
+ 5.44e+10Hz 0.901987 -0.408335
+ 5.45e+10Hz 0.901666 -0.409031
+ 5.46e+10Hz 0.901344 -0.409726
+ 5.47e+10Hz 0.901022 -0.410421
+ 5.48e+10Hz 0.9007 -0.411116
+ 5.49e+10Hz 0.900377 -0.411811
+ 5.5e+10Hz 0.900053 -0.412506
+ 5.51e+10Hz 0.899729 -0.4132
+ 5.52e+10Hz 0.899405 -0.413894
+ 5.53e+10Hz 0.89908 -0.414588
+ 5.54e+10Hz 0.898755 -0.415282
+ 5.55e+10Hz 0.898429 -0.415976
+ 5.56e+10Hz 0.898103 -0.416669
+ 5.57e+10Hz 0.897776 -0.417362
+ 5.58e+10Hz 0.897449 -0.418055
+ 5.59e+10Hz 0.897121 -0.418748
+ 5.6e+10Hz 0.896793 -0.41944
+ 5.61e+10Hz 0.896465 -0.420133
+ 5.62e+10Hz 0.896135 -0.420825
+ 5.63e+10Hz 0.895806 -0.421517
+ 5.64e+10Hz 0.895476 -0.422209
+ 5.65e+10Hz 0.895145 -0.4229
+ 5.66e+10Hz 0.894814 -0.423592
+ 5.67e+10Hz 0.894483 -0.424283
+ 5.68e+10Hz 0.894151 -0.424974
+ 5.69e+10Hz 0.893819 -0.425665
+ 5.7e+10Hz 0.893486 -0.426355
+ 5.71e+10Hz 0.893152 -0.427046
+ 5.72e+10Hz 0.892818 -0.427736
+ 5.73e+10Hz 0.892484 -0.428426
+ 5.74e+10Hz 0.892149 -0.429116
+ 5.75e+10Hz 0.891814 -0.429805
+ 5.76e+10Hz 0.891478 -0.430495
+ 5.77e+10Hz 0.891141 -0.431184
+ 5.78e+10Hz 0.890805 -0.431873
+ 5.79e+10Hz 0.890467 -0.432562
+ 5.8e+10Hz 0.890129 -0.433251
+ 5.81e+10Hz 0.889791 -0.433939
+ 5.82e+10Hz 0.889452 -0.434628
+ 5.83e+10Hz 0.889112 -0.435316
+ 5.84e+10Hz 0.888772 -0.436004
+ 5.85e+10Hz 0.888432 -0.436692
+ 5.86e+10Hz 0.888091 -0.43738
+ 5.87e+10Hz 0.887749 -0.438067
+ 5.88e+10Hz 0.887407 -0.438754
+ 5.89e+10Hz 0.887064 -0.439441
+ 5.9e+10Hz 0.886721 -0.440128
+ 5.91e+10Hz 0.886378 -0.440815
+ 5.92e+10Hz 0.886033 -0.441501
+ 5.93e+10Hz 0.885689 -0.442188
+ 5.94e+10Hz 0.885343 -0.442874
+ 5.95e+10Hz 0.884997 -0.44356
+ 5.96e+10Hz 0.884651 -0.444246
+ 5.97e+10Hz 0.884304 -0.444931
+ 5.98e+10Hz 0.883956 -0.445617
+ 5.99e+10Hz 0.883608 -0.446302
+ 6e+10Hz 0.88326 -0.446987
+ 6.01e+10Hz 0.882911 -0.447671
+ 6.02e+10Hz 0.882561 -0.448356
+ 6.03e+10Hz 0.88221 -0.44904
+ 6.04e+10Hz 0.88186 -0.449725
+ 6.05e+10Hz 0.881508 -0.450409
+ 6.06e+10Hz 0.881156 -0.451092
+ 6.07e+10Hz 0.880804 -0.451776
+ 6.08e+10Hz 0.88045 -0.452459
+ 6.09e+10Hz 0.880097 -0.453142
+ 6.1e+10Hz 0.879742 -0.453825
+ 6.11e+10Hz 0.879388 -0.454508
+ 6.12e+10Hz 0.879032 -0.45519
+ 6.13e+10Hz 0.878676 -0.455873
+ 6.14e+10Hz 0.87832 -0.456555
+ 6.15e+10Hz 0.877962 -0.457237
+ 6.16e+10Hz 0.877605 -0.457918
+ 6.17e+10Hz 0.877246 -0.458599
+ 6.18e+10Hz 0.876887 -0.459281
+ 6.19e+10Hz 0.876528 -0.459962
+ 6.2e+10Hz 0.876168 -0.460642
+ 6.21e+10Hz 0.875807 -0.461323
+ 6.22e+10Hz 0.875446 -0.462003
+ 6.23e+10Hz 0.875084 -0.462683
+ 6.24e+10Hz 0.874721 -0.463362
+ 6.25e+10Hz 0.874358 -0.464042
+ 6.26e+10Hz 0.873995 -0.464721
+ 6.27e+10Hz 0.87363 -0.4654
+ 6.28e+10Hz 0.873265 -0.466079
+ 6.29e+10Hz 0.8729 -0.466757
+ 6.3e+10Hz 0.872534 -0.467435
+ 6.31e+10Hz 0.872167 -0.468113
+ 6.32e+10Hz 0.8718 -0.468791
+ 6.33e+10Hz 0.871432 -0.469468
+ 6.34e+10Hz 0.871064 -0.470146
+ 6.35e+10Hz 0.870695 -0.470822
+ 6.36e+10Hz 0.870325 -0.471499
+ 6.37e+10Hz 0.869955 -0.472175
+ 6.38e+10Hz 0.869584 -0.472851
+ 6.39e+10Hz 0.869213 -0.473527
+ 6.4e+10Hz 0.868841 -0.474202
+ 6.41e+10Hz 0.868468 -0.474878
+ 6.42e+10Hz 0.868095 -0.475552
+ 6.43e+10Hz 0.867721 -0.476227
+ 6.44e+10Hz 0.867347 -0.476901
+ 6.45e+10Hz 0.866972 -0.477575
+ 6.46e+10Hz 0.866596 -0.478249
+ 6.47e+10Hz 0.86622 -0.478922
+ 6.48e+10Hz 0.865843 -0.479595
+ 6.49e+10Hz 0.865466 -0.480268
+ 6.5e+10Hz 0.865088 -0.480941
+ 6.51e+10Hz 0.864709 -0.481613
+ 6.52e+10Hz 0.86433 -0.482284
+ 6.53e+10Hz 0.863951 -0.482956
+ 6.54e+10Hz 0.86357 -0.483627
+ 6.55e+10Hz 0.863189 -0.484298
+ 6.56e+10Hz 0.862808 -0.484969
+ 6.57e+10Hz 0.862426 -0.485639
+ 6.58e+10Hz 0.862043 -0.486309
+ 6.59e+10Hz 0.86166 -0.486978
+ 6.6e+10Hz 0.861276 -0.487647
+ 6.61e+10Hz 0.860892 -0.488316
+ 6.62e+10Hz 0.860507 -0.488985
+ 6.63e+10Hz 0.860121 -0.489653
+ 6.64e+10Hz 0.859735 -0.490321
+ 6.65e+10Hz 0.859349 -0.490988
+ 6.66e+10Hz 0.858961 -0.491655
+ 6.67e+10Hz 0.858573 -0.492322
+ 6.68e+10Hz 0.858185 -0.492988
+ 6.69e+10Hz 0.857796 -0.493655
+ 6.7e+10Hz 0.857407 -0.49432
+ 6.71e+10Hz 0.857017 -0.494986
+ 6.72e+10Hz 0.856626 -0.495651
+ 6.73e+10Hz 0.856235 -0.496315
+ 6.74e+10Hz 0.855843 -0.49698
+ 6.75e+10Hz 0.855451 -0.497643
+ 6.76e+10Hz 0.855058 -0.498307
+ 6.77e+10Hz 0.854665 -0.49897
+ 6.78e+10Hz 0.854271 -0.499633
+ 6.79e+10Hz 0.853876 -0.500295
+ 6.8e+10Hz 0.853481 -0.500958
+ 6.81e+10Hz 0.853085 -0.501619
+ 6.82e+10Hz 0.852689 -0.502281
+ 6.83e+10Hz 0.852293 -0.502942
+ 6.84e+10Hz 0.851896 -0.503602
+ 6.85e+10Hz 0.851498 -0.504262
+ 6.86e+10Hz 0.8511 -0.504922
+ 6.87e+10Hz 0.850701 -0.505582
+ 6.88e+10Hz 0.850302 -0.506241
+ 6.89e+10Hz 0.849902 -0.506899
+ 6.9e+10Hz 0.849501 -0.507558
+ 6.91e+10Hz 0.849101 -0.508216
+ 6.92e+10Hz 0.848699 -0.508873
+ 6.93e+10Hz 0.848297 -0.509531
+ 6.94e+10Hz 0.847895 -0.510187
+ 6.95e+10Hz 0.847492 -0.510844
+ 6.96e+10Hz 0.847089 -0.5115
+ 6.97e+10Hz 0.846685 -0.512156
+ 6.98e+10Hz 0.84628 -0.512811
+ 6.99e+10Hz 0.845875 -0.513466
+ 7e+10Hz 0.84547 -0.51412
+ 7.01e+10Hz 0.845064 -0.514774
+ 7.02e+10Hz 0.844658 -0.515428
+ 7.03e+10Hz 0.844251 -0.516082
+ 7.04e+10Hz 0.843843 -0.516735
+ 7.05e+10Hz 0.843436 -0.517387
+ 7.06e+10Hz 0.843027 -0.518039
+ 7.07e+10Hz 0.842618 -0.518691
+ 7.08e+10Hz 0.842209 -0.519343
+ 7.09e+10Hz 0.841799 -0.519994
+ 7.1e+10Hz 0.841389 -0.520645
+ 7.11e+10Hz 0.840978 -0.521295
+ 7.12e+10Hz 0.840567 -0.521945
+ 7.13e+10Hz 0.840155 -0.522595
+ 7.14e+10Hz 0.839743 -0.523244
+ 7.15e+10Hz 0.839331 -0.523893
+ 7.16e+10Hz 0.838918 -0.524541
+ 7.17e+10Hz 0.838504 -0.525189
+ 7.18e+10Hz 0.83809 -0.525837
+ 7.19e+10Hz 0.837676 -0.526484
+ 7.2e+10Hz 0.837261 -0.527131
+ 7.21e+10Hz 0.836845 -0.527778
+ 7.22e+10Hz 0.836429 -0.528424
+ 7.23e+10Hz 0.836013 -0.52907
+ 7.24e+10Hz 0.835596 -0.529716
+ 7.25e+10Hz 0.835179 -0.530361
+ 7.26e+10Hz 0.834762 -0.531005
+ 7.27e+10Hz 0.834343 -0.53165
+ 7.28e+10Hz 0.833925 -0.532294
+ 7.29e+10Hz 0.833506 -0.532938
+ 7.3e+10Hz 0.833087 -0.533581
+ 7.31e+10Hz 0.832667 -0.534224
+ 7.32e+10Hz 0.832246 -0.534867
+ 7.33e+10Hz 0.831826 -0.535509
+ 7.34e+10Hz 0.831404 -0.536151
+ 7.35e+10Hz 0.830983 -0.536792
+ 7.36e+10Hz 0.830561 -0.537434
+ 7.37e+10Hz 0.830138 -0.538075
+ 7.38e+10Hz 0.829715 -0.538715
+ 7.39e+10Hz 0.829292 -0.539355
+ 7.4e+10Hz 0.828868 -0.539995
+ 7.41e+10Hz 0.828444 -0.540635
+ 7.42e+10Hz 0.828019 -0.541274
+ 7.43e+10Hz 0.827594 -0.541913
+ 7.44e+10Hz 0.827168 -0.542551
+ 7.45e+10Hz 0.826742 -0.543189
+ 7.46e+10Hz 0.826316 -0.543827
+ 7.47e+10Hz 0.825889 -0.544465
+ 7.48e+10Hz 0.825462 -0.545102
+ 7.49e+10Hz 0.825034 -0.545739
+ 7.5e+10Hz 0.824606 -0.546375
+ 7.51e+10Hz 0.824177 -0.547011
+ 7.52e+10Hz 0.823748 -0.547647
+ 7.53e+10Hz 0.823318 -0.548283
+ 7.54e+10Hz 0.822888 -0.548918
+ 7.55e+10Hz 0.822458 -0.549553
+ 7.56e+10Hz 0.822027 -0.550187
+ 7.57e+10Hz 0.821596 -0.550821
+ 7.58e+10Hz 0.821164 -0.551455
+ 7.59e+10Hz 0.820732 -0.552089
+ 7.6e+10Hz 0.8203 -0.552722
+ 7.61e+10Hz 0.819867 -0.553355
+ 7.62e+10Hz 0.819433 -0.553988
+ 7.63e+10Hz 0.819 -0.55462
+ 7.64e+10Hz 0.818565 -0.555252
+ 7.65e+10Hz 0.818131 -0.555884
+ 7.66e+10Hz 0.817695 -0.556515
+ 7.67e+10Hz 0.81726 -0.557146
+ 7.68e+10Hz 0.816824 -0.557777
+ 7.69e+10Hz 0.816387 -0.558408
+ 7.7e+10Hz 0.81595 -0.559038
+ 7.71e+10Hz 0.815513 -0.559668
+ 7.72e+10Hz 0.815075 -0.560297
+ 7.73e+10Hz 0.814637 -0.560926
+ 7.74e+10Hz 0.814198 -0.561555
+ 7.75e+10Hz 0.813759 -0.562184
+ 7.76e+10Hz 0.813319 -0.562812
+ 7.77e+10Hz 0.812879 -0.563441
+ 7.78e+10Hz 0.812439 -0.564068
+ 7.79e+10Hz 0.811998 -0.564696
+ 7.8e+10Hz 0.811556 -0.565323
+ 7.81e+10Hz 0.811114 -0.56595
+ 7.82e+10Hz 0.810672 -0.566576
+ 7.83e+10Hz 0.810229 -0.567203
+ 7.84e+10Hz 0.809786 -0.567829
+ 7.85e+10Hz 0.809342 -0.568454
+ 7.86e+10Hz 0.808898 -0.56908
+ 7.87e+10Hz 0.808453 -0.569705
+ 7.88e+10Hz 0.808008 -0.57033
+ 7.89e+10Hz 0.807563 -0.570954
+ 7.9e+10Hz 0.807117 -0.571579
+ 7.91e+10Hz 0.80667 -0.572202
+ 7.92e+10Hz 0.806223 -0.572826
+ 7.93e+10Hz 0.805776 -0.573449
+ 7.94e+10Hz 0.805328 -0.574072
+ 7.95e+10Hz 0.804879 -0.574695
+ 7.96e+10Hz 0.804431 -0.575318
+ 7.97e+10Hz 0.803981 -0.57594
+ 7.98e+10Hz 0.803531 -0.576562
+ 7.99e+10Hz 0.803081 -0.577183
+ 8e+10Hz 0.80263 -0.577805
+ 8.01e+10Hz 0.802179 -0.578426
+ 8.02e+10Hz 0.801727 -0.579046
+ 8.03e+10Hz 0.801275 -0.579667
+ 8.04e+10Hz 0.800822 -0.580287
+ 8.05e+10Hz 0.800369 -0.580907
+ 8.06e+10Hz 0.799915 -0.581526
+ 8.07e+10Hz 0.799461 -0.582145
+ 8.08e+10Hz 0.799006 -0.582764
+ 8.09e+10Hz 0.798551 -0.583383
+ 8.1e+10Hz 0.798095 -0.584001
+ 8.11e+10Hz 0.797639 -0.584619
+ 8.12e+10Hz 0.797182 -0.585237
+ 8.13e+10Hz 0.796725 -0.585854
+ 8.14e+10Hz 0.796267 -0.586471
+ 8.15e+10Hz 0.795809 -0.587088
+ 8.16e+10Hz 0.795351 -0.587704
+ 8.17e+10Hz 0.794891 -0.58832
+ 8.18e+10Hz 0.794432 -0.588936
+ 8.19e+10Hz 0.793971 -0.589552
+ 8.2e+10Hz 0.793511 -0.590167
+ 8.21e+10Hz 0.793049 -0.590782
+ 8.22e+10Hz 0.792588 -0.591396
+ 8.23e+10Hz 0.792125 -0.592011
+ 8.24e+10Hz 0.791663 -0.592625
+ 8.25e+10Hz 0.791199 -0.593238
+ 8.26e+10Hz 0.790736 -0.593852
+ 8.27e+10Hz 0.790271 -0.594464
+ 8.28e+10Hz 0.789806 -0.595077
+ 8.29e+10Hz 0.789341 -0.595689
+ 8.3e+10Hz 0.788875 -0.596301
+ 8.31e+10Hz 0.788409 -0.596913
+ 8.32e+10Hz 0.787942 -0.597524
+ 8.33e+10Hz 0.787475 -0.598135
+ 8.34e+10Hz 0.787007 -0.598746
+ 8.35e+10Hz 0.786538 -0.599356
+ 8.36e+10Hz 0.786069 -0.599966
+ 8.37e+10Hz 0.7856 -0.600576
+ 8.38e+10Hz 0.78513 -0.601185
+ 8.39e+10Hz 0.784659 -0.601794
+ 8.4e+10Hz 0.784188 -0.602403
+ 8.41e+10Hz 0.783716 -0.603011
+ 8.42e+10Hz 0.783244 -0.603619
+ 8.43e+10Hz 0.782772 -0.604226
+ 8.44e+10Hz 0.782299 -0.604833
+ 8.45e+10Hz 0.781825 -0.60544
+ 8.46e+10Hz 0.781351 -0.606047
+ 8.47e+10Hz 0.780876 -0.606653
+ 8.48e+10Hz 0.780401 -0.607259
+ 8.49e+10Hz 0.779925 -0.607864
+ 8.5e+10Hz 0.779449 -0.608469
+ 8.51e+10Hz 0.778972 -0.609074
+ 8.52e+10Hz 0.778495 -0.609678
+ 8.53e+10Hz 0.778017 -0.610282
+ 8.54e+10Hz 0.777539 -0.610885
+ 8.55e+10Hz 0.77706 -0.611488
+ 8.56e+10Hz 0.77658 -0.612091
+ 8.57e+10Hz 0.7761 -0.612693
+ 8.58e+10Hz 0.77562 -0.613295
+ 8.59e+10Hz 0.775139 -0.613897
+ 8.6e+10Hz 0.774657 -0.614498
+ 8.61e+10Hz 0.774176 -0.615099
+ 8.62e+10Hz 0.773693 -0.6157
+ 8.63e+10Hz 0.77321 -0.6163
+ 8.64e+10Hz 0.772726 -0.616899
+ 8.65e+10Hz 0.772242 -0.617499
+ 8.66e+10Hz 0.771758 -0.618098
+ 8.67e+10Hz 0.771273 -0.618696
+ 8.68e+10Hz 0.770787 -0.619294
+ 8.69e+10Hz 0.770301 -0.619892
+ 8.7e+10Hz 0.769815 -0.620489
+ 8.71e+10Hz 0.769327 -0.621086
+ 8.72e+10Hz 0.76884 -0.621682
+ 8.73e+10Hz 0.768352 -0.622278
+ 8.74e+10Hz 0.767863 -0.622874
+ 8.75e+10Hz 0.767374 -0.623469
+ 8.76e+10Hz 0.766884 -0.624064
+ 8.77e+10Hz 0.766394 -0.624659
+ 8.78e+10Hz 0.765904 -0.625253
+ 8.79e+10Hz 0.765413 -0.625846
+ 8.8e+10Hz 0.764921 -0.626439
+ 8.81e+10Hz 0.764429 -0.627032
+ 8.82e+10Hz 0.763936 -0.627624
+ 8.83e+10Hz 0.763443 -0.628216
+ 8.84e+10Hz 0.76295 -0.628808
+ 8.85e+10Hz 0.762456 -0.629399
+ 8.86e+10Hz 0.761961 -0.629989
+ 8.87e+10Hz 0.761466 -0.63058
+ 8.88e+10Hz 0.760971 -0.631169
+ 8.89e+10Hz 0.760475 -0.631759
+ 8.9e+10Hz 0.759978 -0.632348
+ 8.91e+10Hz 0.759481 -0.632936
+ 8.92e+10Hz 0.758984 -0.633524
+ 8.93e+10Hz 0.758486 -0.634112
+ 8.94e+10Hz 0.757987 -0.634699
+ 8.95e+10Hz 0.757489 -0.635286
+ 8.96e+10Hz 0.756989 -0.635872
+ 8.97e+10Hz 0.756489 -0.636458
+ 8.98e+10Hz 0.755989 -0.637043
+ 8.99e+10Hz 0.755489 -0.637628
+ 9e+10Hz 0.754987 -0.638213
+ 9.01e+10Hz 0.754486 -0.638797
+ 9.02e+10Hz 0.753984 -0.639381
+ 9.03e+10Hz 0.753481 -0.639964
+ 9.04e+10Hz 0.752978 -0.640547
+ 9.05e+10Hz 0.752475 -0.641129
+ 9.06e+10Hz 0.751971 -0.641711
+ 9.07e+10Hz 0.751466 -0.642292
+ 9.08e+10Hz 0.750961 -0.642873
+ 9.09e+10Hz 0.750456 -0.643454
+ 9.1e+10Hz 0.749951 -0.644034
+ 9.11e+10Hz 0.749444 -0.644614
+ 9.12e+10Hz 0.748938 -0.645193
+ 9.13e+10Hz 0.748431 -0.645772
+ 9.14e+10Hz 0.747923 -0.646351
+ 9.15e+10Hz 0.747415 -0.646928
+ 9.16e+10Hz 0.746907 -0.647506
+ 9.17e+10Hz 0.746398 -0.648083
+ 9.18e+10Hz 0.745889 -0.64866
+ 9.19e+10Hz 0.745379 -0.649236
+ 9.2e+10Hz 0.744869 -0.649812
+ 9.21e+10Hz 0.744359 -0.650387
+ 9.22e+10Hz 0.743848 -0.650962
+ 9.23e+10Hz 0.743337 -0.651536
+ 9.24e+10Hz 0.742825 -0.65211
+ 9.25e+10Hz 0.742313 -0.652684
+ 9.26e+10Hz 0.7418 -0.653257
+ 9.27e+10Hz 0.741287 -0.65383
+ 9.28e+10Hz 0.740774 -0.654402
+ 9.29e+10Hz 0.74026 -0.654974
+ 9.3e+10Hz 0.739745 -0.655545
+ 9.31e+10Hz 0.739231 -0.656116
+ 9.32e+10Hz 0.738716 -0.656687
+ 9.33e+10Hz 0.7382 -0.657257
+ 9.34e+10Hz 0.737684 -0.657827
+ 9.35e+10Hz 0.737168 -0.658396
+ 9.36e+10Hz 0.736651 -0.658965
+ 9.37e+10Hz 0.736134 -0.659533
+ 9.38e+10Hz 0.735617 -0.660101
+ 9.39e+10Hz 0.735099 -0.660668
+ 9.4e+10Hz 0.73458 -0.661235
+ 9.41e+10Hz 0.734062 -0.661802
+ 9.42e+10Hz 0.733542 -0.662368
+ 9.43e+10Hz 0.733023 -0.662934
+ 9.44e+10Hz 0.732503 -0.6635
+ 9.45e+10Hz 0.731983 -0.664065
+ 9.46e+10Hz 0.731462 -0.664629
+ 9.47e+10Hz 0.730941 -0.665193
+ 9.48e+10Hz 0.730419 -0.665757
+ 9.49e+10Hz 0.729897 -0.66632
+ 9.5e+10Hz 0.729375 -0.666883
+ 9.51e+10Hz 0.728852 -0.667446
+ 9.52e+10Hz 0.728329 -0.668008
+ 9.53e+10Hz 0.727806 -0.668569
+ 9.54e+10Hz 0.727282 -0.669131
+ 9.55e+10Hz 0.726758 -0.669691
+ 9.56e+10Hz 0.726233 -0.670252
+ 9.57e+10Hz 0.725708 -0.670812
+ 9.58e+10Hz 0.725182 -0.671371
+ 9.59e+10Hz 0.724657 -0.671931
+ 9.6e+10Hz 0.72413 -0.672489
+ 9.61e+10Hz 0.723604 -0.673048
+ 9.62e+10Hz 0.723077 -0.673606
+ 9.63e+10Hz 0.722549 -0.674163
+ 9.64e+10Hz 0.722022 -0.67472
+ 9.65e+10Hz 0.721493 -0.675277
+ 9.66e+10Hz 0.720965 -0.675833
+ 9.67e+10Hz 0.720436 -0.676389
+ 9.68e+10Hz 0.719906 -0.676945
+ 9.69e+10Hz 0.719377 -0.6775
+ 9.7e+10Hz 0.718847 -0.678055
+ 9.71e+10Hz 0.718316 -0.678609
+ 9.72e+10Hz 0.717785 -0.679163
+ 9.73e+10Hz 0.717254 -0.679717
+ 9.74e+10Hz 0.716722 -0.68027
+ 9.75e+10Hz 0.71619 -0.680823
+ 9.76e+10Hz 0.715658 -0.681375
+ 9.77e+10Hz 0.715125 -0.681927
+ 9.78e+10Hz 0.714591 -0.682479
+ 9.79e+10Hz 0.714058 -0.68303
+ 9.8e+10Hz 0.713524 -0.683581
+ 9.81e+10Hz 0.712989 -0.684132
+ 9.82e+10Hz 0.712454 -0.684682
+ 9.83e+10Hz 0.711919 -0.685231
+ 9.84e+10Hz 0.711383 -0.685781
+ 9.85e+10Hz 0.710847 -0.68633
+ 9.86e+10Hz 0.710311 -0.686878
+ 9.87e+10Hz 0.709774 -0.687426
+ 9.88e+10Hz 0.709237 -0.687974
+ 9.89e+10Hz 0.708699 -0.688521
+ 9.9e+10Hz 0.708161 -0.689068
+ 9.91e+10Hz 0.707623 -0.689615
+ 9.92e+10Hz 0.707084 -0.690161
+ 9.93e+10Hz 0.706545 -0.690707
+ 9.94e+10Hz 0.706005 -0.691253
+ 9.95e+10Hz 0.705465 -0.691798
+ 9.96e+10Hz 0.704924 -0.692343
+ 9.97e+10Hz 0.704383 -0.692887
+ 9.98e+10Hz 0.703842 -0.693431
+ 9.99e+10Hz 0.7033 -0.693975
+ 1e+11Hz 0.702758 -0.694518
+ 1.001e+11Hz 0.702216 -0.695061
+ 1.002e+11Hz 0.701673 -0.695603
+ 1.003e+11Hz 0.70113 -0.696145
+ 1.004e+11Hz 0.700586 -0.696687
+ 1.005e+11Hz 0.700042 -0.697228
+ 1.006e+11Hz 0.699497 -0.697769
+ 1.007e+11Hz 0.698952 -0.69831
+ 1.008e+11Hz 0.698407 -0.69885
+ 1.009e+11Hz 0.697861 -0.69939
+ 1.01e+11Hz 0.697314 -0.699929
+ 1.011e+11Hz 0.696768 -0.700468
+ 1.012e+11Hz 0.696221 -0.701007
+ 1.013e+11Hz 0.695673 -0.701545
+ 1.014e+11Hz 0.695125 -0.702083
+ 1.015e+11Hz 0.694577 -0.702621
+ 1.016e+11Hz 0.694028 -0.703158
+ 1.017e+11Hz 0.693479 -0.703694
+ 1.018e+11Hz 0.692929 -0.704231
+ 1.019e+11Hz 0.692379 -0.704767
+ 1.02e+11Hz 0.691828 -0.705302
+ 1.021e+11Hz 0.691277 -0.705838
+ 1.022e+11Hz 0.690726 -0.706373
+ 1.023e+11Hz 0.690174 -0.706907
+ 1.024e+11Hz 0.689622 -0.707441
+ 1.025e+11Hz 0.689069 -0.707975
+ 1.026e+11Hz 0.688516 -0.708508
+ 1.027e+11Hz 0.687962 -0.709041
+ 1.028e+11Hz 0.687408 -0.709573
+ 1.029e+11Hz 0.686854 -0.710106
+ 1.03e+11Hz 0.686299 -0.710637
+ 1.031e+11Hz 0.685743 -0.711169
+ 1.032e+11Hz 0.685188 -0.711699
+ 1.033e+11Hz 0.684631 -0.71223
+ 1.034e+11Hz 0.684075 -0.71276
+ 1.035e+11Hz 0.683518 -0.71329
+ 1.036e+11Hz 0.68296 -0.713819
+ 1.037e+11Hz 0.682402 -0.714348
+ 1.038e+11Hz 0.681844 -0.714877
+ 1.039e+11Hz 0.681285 -0.715405
+ 1.04e+11Hz 0.680725 -0.715932
+ 1.041e+11Hz 0.680165 -0.71646
+ 1.042e+11Hz 0.679605 -0.716987
+ 1.043e+11Hz 0.679044 -0.717513
+ 1.044e+11Hz 0.678483 -0.718039
+ 1.045e+11Hz 0.677922 -0.718565
+ 1.046e+11Hz 0.67736 -0.71909
+ 1.047e+11Hz 0.676797 -0.719615
+ 1.048e+11Hz 0.676234 -0.720139
+ 1.049e+11Hz 0.675671 -0.720663
+ 1.05e+11Hz 0.675107 -0.721187
+ 1.051e+11Hz 0.674543 -0.72171
+ 1.052e+11Hz 0.673978 -0.722233
+ 1.053e+11Hz 0.673413 -0.722755
+ 1.054e+11Hz 0.672847 -0.723277
+ 1.055e+11Hz 0.672281 -0.723799
+ 1.056e+11Hz 0.671714 -0.72432
+ 1.057e+11Hz 0.671147 -0.72484
+ 1.058e+11Hz 0.67058 -0.72536
+ 1.059e+11Hz 0.670012 -0.72588
+ 1.06e+11Hz 0.669444 -0.7264
+ 1.061e+11Hz 0.668875 -0.726918
+ 1.062e+11Hz 0.668305 -0.727437
+ 1.063e+11Hz 0.667736 -0.727955
+ 1.064e+11Hz 0.667166 -0.728472
+ 1.065e+11Hz 0.666595 -0.728989
+ 1.066e+11Hz 0.666024 -0.729506
+ 1.067e+11Hz 0.665452 -0.730022
+ 1.068e+11Hz 0.66488 -0.730538
+ 1.069e+11Hz 0.664308 -0.731053
+ 1.07e+11Hz 0.663735 -0.731568
+ 1.071e+11Hz 0.663162 -0.732083
+ 1.072e+11Hz 0.662588 -0.732597
+ 1.073e+11Hz 0.662014 -0.73311
+ 1.074e+11Hz 0.661439 -0.733623
+ 1.075e+11Hz 0.660864 -0.734136
+ 1.076e+11Hz 0.660288 -0.734648
+ 1.077e+11Hz 0.659712 -0.73516
+ 1.078e+11Hz 0.659136 -0.735671
+ 1.079e+11Hz 0.658559 -0.736182
+ 1.08e+11Hz 0.657982 -0.736692
+ 1.081e+11Hz 0.657404 -0.737202
+ 1.082e+11Hz 0.656826 -0.737711
+ 1.083e+11Hz 0.656247 -0.73822
+ 1.084e+11Hz 0.655668 -0.738728
+ 1.085e+11Hz 0.655088 -0.739236
+ 1.086e+11Hz 0.654508 -0.739744
+ 1.087e+11Hz 0.653928 -0.740251
+ 1.088e+11Hz 0.653347 -0.740757
+ 1.089e+11Hz 0.652766 -0.741263
+ 1.09e+11Hz 0.652184 -0.741769
+ 1.091e+11Hz 0.651602 -0.742274
+ 1.092e+11Hz 0.65102 -0.742778
+ 1.093e+11Hz 0.650437 -0.743282
+ 1.094e+11Hz 0.649853 -0.743786
+ 1.095e+11Hz 0.649269 -0.744289
+ 1.096e+11Hz 0.648685 -0.744792
+ 1.097e+11Hz 0.6481 -0.745294
+ 1.098e+11Hz 0.647515 -0.745796
+ 1.099e+11Hz 0.64693 -0.746297
+ 1.1e+11Hz 0.646344 -0.746797
+ 1.101e+11Hz 0.645757 -0.747298
+ 1.102e+11Hz 0.645171 -0.747797
+ 1.103e+11Hz 0.644583 -0.748297
+ 1.104e+11Hz 0.643996 -0.748795
+ 1.105e+11Hz 0.643408 -0.749293
+ 1.106e+11Hz 0.642819 -0.749791
+ 1.107e+11Hz 0.642231 -0.750288
+ 1.108e+11Hz 0.641641 -0.750785
+ 1.109e+11Hz 0.641052 -0.751281
+ 1.11e+11Hz 0.640462 -0.751777
+ 1.111e+11Hz 0.639871 -0.752272
+ 1.112e+11Hz 0.63928 -0.752767
+ 1.113e+11Hz 0.638689 -0.753261
+ 1.114e+11Hz 0.638097 -0.753755
+ 1.115e+11Hz 0.637505 -0.754248
+ 1.116e+11Hz 0.636913 -0.754741
+ 1.117e+11Hz 0.63632 -0.755233
+ 1.118e+11Hz 0.635727 -0.755725
+ 1.119e+11Hz 0.635133 -0.756216
+ 1.12e+11Hz 0.634539 -0.756707
+ 1.121e+11Hz 0.633944 -0.757197
+ 1.122e+11Hz 0.63335 -0.757687
+ 1.123e+11Hz 0.632754 -0.758176
+ 1.124e+11Hz 0.632159 -0.758665
+ 1.125e+11Hz 0.631563 -0.759153
+ 1.126e+11Hz 0.630966 -0.75964
+ 1.127e+11Hz 0.63037 -0.760128
+ 1.128e+11Hz 0.629773 -0.760614
+ 1.129e+11Hz 0.629175 -0.761101
+ 1.13e+11Hz 0.628577 -0.761586
+ 1.131e+11Hz 0.627979 -0.762071
+ 1.132e+11Hz 0.62738 -0.762556
+ 1.133e+11Hz 0.626781 -0.76304
+ 1.134e+11Hz 0.626182 -0.763524
+ 1.135e+11Hz 0.625582 -0.764007
+ 1.136e+11Hz 0.624982 -0.76449
+ 1.137e+11Hz 0.624382 -0.764972
+ 1.138e+11Hz 0.623781 -0.765453
+ 1.139e+11Hz 0.62318 -0.765935
+ 1.14e+11Hz 0.622578 -0.766415
+ 1.141e+11Hz 0.621976 -0.766895
+ 1.142e+11Hz 0.621374 -0.767375
+ 1.143e+11Hz 0.620771 -0.767854
+ 1.144e+11Hz 0.620168 -0.768333
+ 1.145e+11Hz 0.619565 -0.768811
+ 1.146e+11Hz 0.618961 -0.769288
+ 1.147e+11Hz 0.618357 -0.769766
+ 1.148e+11Hz 0.617753 -0.770242
+ 1.149e+11Hz 0.617148 -0.770718
+ 1.15e+11Hz 0.616543 -0.771194
+ 1.151e+11Hz 0.615938 -0.771669
+ 1.152e+11Hz 0.615332 -0.772144
+ 1.153e+11Hz 0.614726 -0.772618
+ 1.154e+11Hz 0.614119 -0.773091
+ 1.155e+11Hz 0.613512 -0.773565
+ 1.156e+11Hz 0.612905 -0.774037
+ 1.157e+11Hz 0.612298 -0.774509
+ 1.158e+11Hz 0.61169 -0.774981
+ 1.159e+11Hz 0.611081 -0.775452
+ 1.16e+11Hz 0.610473 -0.775923
+ 1.161e+11Hz 0.609864 -0.776393
+ 1.162e+11Hz 0.609255 -0.776863
+ 1.163e+11Hz 0.608645 -0.777332
+ 1.164e+11Hz 0.608035 -0.777801
+ 1.165e+11Hz 0.607425 -0.778269
+ 1.166e+11Hz 0.606814 -0.778737
+ 1.167e+11Hz 0.606203 -0.779204
+ 1.168e+11Hz 0.605592 -0.779671
+ 1.169e+11Hz 0.60498 -0.780137
+ 1.17e+11Hz 0.604368 -0.780603
+ 1.171e+11Hz 0.603756 -0.781068
+ 1.172e+11Hz 0.603144 -0.781533
+ 1.173e+11Hz 0.602531 -0.781997
+ 1.174e+11Hz 0.601917 -0.782461
+ 1.175e+11Hz 0.601304 -0.782925
+ 1.176e+11Hz 0.60069 -0.783388
+ 1.177e+11Hz 0.600075 -0.78385
+ 1.178e+11Hz 0.599461 -0.784312
+ 1.179e+11Hz 0.598846 -0.784774
+ 1.18e+11Hz 0.59823 -0.785235
+ 1.181e+11Hz 0.597615 -0.785695
+ 1.182e+11Hz 0.596999 -0.786155
+ 1.183e+11Hz 0.596382 -0.786615
+ 1.184e+11Hz 0.595766 -0.787074
+ 1.185e+11Hz 0.595149 -0.787533
+ 1.186e+11Hz 0.594531 -0.787991
+ 1.187e+11Hz 0.593914 -0.788448
+ 1.188e+11Hz 0.593296 -0.788906
+ 1.189e+11Hz 0.592677 -0.789362
+ 1.19e+11Hz 0.592059 -0.789819
+ 1.191e+11Hz 0.59144 -0.790274
+ 1.192e+11Hz 0.59082 -0.79073
+ 1.193e+11Hz 0.590201 -0.791185
+ 1.194e+11Hz 0.589581 -0.791639
+ 1.195e+11Hz 0.58896 -0.792093
+ 1.196e+11Hz 0.58834 -0.792547
+ 1.197e+11Hz 0.587719 -0.793
+ 1.198e+11Hz 0.587097 -0.793452
+ 1.199e+11Hz 0.586475 -0.793904
+ 1.2e+11Hz 0.585853 -0.794356
+ 1.201e+11Hz 0.585231 -0.794807
+ 1.202e+11Hz 0.584608 -0.795258
+ 1.203e+11Hz 0.583985 -0.795708
+ 1.204e+11Hz 0.583362 -0.796158
+ 1.205e+11Hz 0.582738 -0.796607
+ 1.206e+11Hz 0.582114 -0.797056
+ 1.207e+11Hz 0.58149 -0.797504
+ 1.208e+11Hz 0.580865 -0.797952
+ 1.209e+11Hz 0.58024 -0.798399
+ 1.21e+11Hz 0.579614 -0.798846
+ 1.211e+11Hz 0.578988 -0.799293
+ 1.212e+11Hz 0.578362 -0.799739
+ 1.213e+11Hz 0.577736 -0.800185
+ 1.214e+11Hz 0.577109 -0.80063
+ 1.215e+11Hz 0.576482 -0.801074
+ 1.216e+11Hz 0.575854 -0.801519
+ 1.217e+11Hz 0.575226 -0.801962
+ 1.218e+11Hz 0.574598 -0.802406
+ 1.219e+11Hz 0.573969 -0.802848
+ 1.22e+11Hz 0.57334 -0.803291
+ 1.221e+11Hz 0.572711 -0.803733
+ 1.222e+11Hz 0.572081 -0.804174
+ 1.223e+11Hz 0.571451 -0.804615
+ 1.224e+11Hz 0.570821 -0.805055
+ 1.225e+11Hz 0.57019 -0.805495
+ 1.226e+11Hz 0.569559 -0.805935
+ 1.227e+11Hz 0.568928 -0.806374
+ 1.228e+11Hz 0.568296 -0.806813
+ 1.229e+11Hz 0.567664 -0.807251
+ 1.23e+11Hz 0.567032 -0.807689
+ 1.231e+11Hz 0.566399 -0.808126
+ 1.232e+11Hz 0.565765 -0.808563
+ 1.233e+11Hz 0.565132 -0.808999
+ 1.234e+11Hz 0.564498 -0.809435
+ 1.235e+11Hz 0.563864 -0.80987
+ 1.236e+11Hz 0.563229 -0.810305
+ 1.237e+11Hz 0.562594 -0.810739
+ 1.238e+11Hz 0.561959 -0.811173
+ 1.239e+11Hz 0.561323 -0.811607
+ 1.24e+11Hz 0.560687 -0.81204
+ 1.241e+11Hz 0.56005 -0.812472
+ 1.242e+11Hz 0.559413 -0.812904
+ 1.243e+11Hz 0.558776 -0.813336
+ 1.244e+11Hz 0.558139 -0.813767
+ 1.245e+11Hz 0.557501 -0.814198
+ 1.246e+11Hz 0.556862 -0.814628
+ 1.247e+11Hz 0.556224 -0.815057
+ 1.248e+11Hz 0.555585 -0.815487
+ 1.249e+11Hz 0.554945 -0.815915
+ 1.25e+11Hz 0.554305 -0.816343
+ 1.251e+11Hz 0.553665 -0.816771
+ 1.252e+11Hz 0.553025 -0.817198
+ 1.253e+11Hz 0.552384 -0.817625
+ 1.254e+11Hz 0.551743 -0.818051
+ 1.255e+11Hz 0.551101 -0.818477
+ 1.256e+11Hz 0.550459 -0.818902
+ 1.257e+11Hz 0.549817 -0.819327
+ 1.258e+11Hz 0.549174 -0.819752
+ 1.259e+11Hz 0.548531 -0.820175
+ 1.26e+11Hz 0.547887 -0.820599
+ 1.261e+11Hz 0.547243 -0.821021
+ 1.262e+11Hz 0.546599 -0.821444
+ 1.263e+11Hz 0.545954 -0.821866
+ 1.264e+11Hz 0.54531 -0.822287
+ 1.265e+11Hz 0.544664 -0.822708
+ 1.266e+11Hz 0.544018 -0.823128
+ 1.267e+11Hz 0.543372 -0.823548
+ 1.268e+11Hz 0.542726 -0.823967
+ 1.269e+11Hz 0.542079 -0.824386
+ 1.27e+11Hz 0.541432 -0.824804
+ 1.271e+11Hz 0.540784 -0.825222
+ 1.272e+11Hz 0.540136 -0.825639
+ 1.273e+11Hz 0.539488 -0.826056
+ 1.274e+11Hz 0.538839 -0.826472
+ 1.275e+11Hz 0.53819 -0.826888
+ 1.276e+11Hz 0.537541 -0.827303
+ 1.277e+11Hz 0.536891 -0.827718
+ 1.278e+11Hz 0.536241 -0.828132
+ 1.279e+11Hz 0.53559 -0.828546
+ 1.28e+11Hz 0.534939 -0.828959
+ 1.281e+11Hz 0.534288 -0.829372
+ 1.282e+11Hz 0.533636 -0.829784
+ 1.283e+11Hz 0.532984 -0.830195
+ 1.284e+11Hz 0.532332 -0.830606
+ 1.285e+11Hz 0.531679 -0.831017
+ 1.286e+11Hz 0.531026 -0.831427
+ 1.287e+11Hz 0.530373 -0.831836
+ 1.288e+11Hz 0.529719 -0.832245
+ 1.289e+11Hz 0.529065 -0.832654
+ 1.29e+11Hz 0.52841 -0.833062
+ 1.291e+11Hz 0.527755 -0.833469
+ 1.292e+11Hz 0.5271 -0.833876
+ 1.293e+11Hz 0.526444 -0.834282
+ 1.294e+11Hz 0.525788 -0.834688
+ 1.295e+11Hz 0.525132 -0.835093
+ 1.296e+11Hz 0.524475 -0.835498
+ 1.297e+11Hz 0.523818 -0.835902
+ 1.298e+11Hz 0.52316 -0.836305
+ 1.299e+11Hz 0.522503 -0.836708
+ 1.3e+11Hz 0.521844 -0.837111
+ 1.301e+11Hz 0.521186 -0.837513
+ 1.302e+11Hz 0.520527 -0.837914
+ 1.303e+11Hz 0.519868 -0.838315
+ 1.304e+11Hz 0.519208 -0.838715
+ 1.305e+11Hz 0.518548 -0.839115
+ 1.306e+11Hz 0.517888 -0.839514
+ 1.307e+11Hz 0.517228 -0.839912
+ 1.308e+11Hz 0.516567 -0.84031
+ 1.309e+11Hz 0.515905 -0.840708
+ 1.31e+11Hz 0.515244 -0.841105
+ 1.311e+11Hz 0.514582 -0.841501
+ 1.312e+11Hz 0.513919 -0.841897
+ 1.313e+11Hz 0.513257 -0.842292
+ 1.314e+11Hz 0.512594 -0.842687
+ 1.315e+11Hz 0.51193 -0.843081
+ 1.316e+11Hz 0.511267 -0.843475
+ 1.317e+11Hz 0.510603 -0.843868
+ 1.318e+11Hz 0.509938 -0.84426
+ 1.319e+11Hz 0.509274 -0.844652
+ 1.32e+11Hz 0.508609 -0.845043
+ 1.321e+11Hz 0.507943 -0.845434
+ 1.322e+11Hz 0.507278 -0.845824
+ 1.323e+11Hz 0.506612 -0.846214
+ 1.324e+11Hz 0.505945 -0.846603
+ 1.325e+11Hz 0.505279 -0.846992
+ 1.326e+11Hz 0.504612 -0.847379
+ 1.327e+11Hz 0.503944 -0.847767
+ 1.328e+11Hz 0.503277 -0.848154
+ 1.329e+11Hz 0.502609 -0.84854
+ 1.33e+11Hz 0.501941 -0.848925
+ 1.331e+11Hz 0.501272 -0.84931
+ 1.332e+11Hz 0.500603 -0.849695
+ 1.333e+11Hz 0.499934 -0.850079
+ 1.334e+11Hz 0.499265 -0.850462
+ 1.335e+11Hz 0.498595 -0.850845
+ 1.336e+11Hz 0.497925 -0.851227
+ 1.337e+11Hz 0.497254 -0.851609
+ 1.338e+11Hz 0.496584 -0.85199
+ 1.339e+11Hz 0.495913 -0.85237
+ 1.34e+11Hz 0.495241 -0.85275
+ 1.341e+11Hz 0.49457 -0.85313
+ 1.342e+11Hz 0.493898 -0.853509
+ 1.343e+11Hz 0.493225 -0.853887
+ 1.344e+11Hz 0.492553 -0.854264
+ 1.345e+11Hz 0.49188 -0.854641
+ 1.346e+11Hz 0.491207 -0.855018
+ 1.347e+11Hz 0.490534 -0.855394
+ 1.348e+11Hz 0.48986 -0.855769
+ 1.349e+11Hz 0.489186 -0.856144
+ 1.35e+11Hz 0.488512 -0.856518
+ 1.351e+11Hz 0.487837 -0.856892
+ 1.352e+11Hz 0.487162 -0.857265
+ 1.353e+11Hz 0.486487 -0.857637
+ 1.354e+11Hz 0.485812 -0.858009
+ 1.355e+11Hz 0.485136 -0.858381
+ 1.356e+11Hz 0.48446 -0.858751
+ 1.357e+11Hz 0.483784 -0.859122
+ 1.358e+11Hz 0.483107 -0.859491
+ 1.359e+11Hz 0.48243 -0.85986
+ 1.36e+11Hz 0.481753 -0.860229
+ 1.361e+11Hz 0.481076 -0.860597
+ 1.362e+11Hz 0.480398 -0.860964
+ 1.363e+11Hz 0.47972 -0.861331
+ 1.364e+11Hz 0.479042 -0.861697
+ 1.365e+11Hz 0.478363 -0.862063
+ 1.366e+11Hz 0.477684 -0.862428
+ 1.367e+11Hz 0.477005 -0.862792
+ 1.368e+11Hz 0.476326 -0.863156
+ 1.369e+11Hz 0.475646 -0.86352
+ 1.37e+11Hz 0.474967 -0.863882
+ 1.371e+11Hz 0.474286 -0.864245
+ 1.372e+11Hz 0.473606 -0.864606
+ 1.373e+11Hz 0.472925 -0.864967
+ 1.374e+11Hz 0.472244 -0.865328
+ 1.375e+11Hz 0.471563 -0.865688
+ 1.376e+11Hz 0.470882 -0.866047
+ 1.377e+11Hz 0.4702 -0.866406
+ 1.378e+11Hz 0.469518 -0.866765
+ 1.379e+11Hz 0.468836 -0.867122
+ 1.38e+11Hz 0.468153 -0.867479
+ 1.381e+11Hz 0.46747 -0.867836
+ 1.382e+11Hz 0.466787 -0.868192
+ 1.383e+11Hz 0.466104 -0.868548
+ 1.384e+11Hz 0.46542 -0.868903
+ 1.385e+11Hz 0.464737 -0.869257
+ 1.386e+11Hz 0.464053 -0.869611
+ 1.387e+11Hz 0.463368 -0.869964
+ 1.388e+11Hz 0.462684 -0.870317
+ 1.389e+11Hz 0.461999 -0.870669
+ 1.39e+11Hz 0.461314 -0.871021
+ 1.391e+11Hz 0.460628 -0.871372
+ 1.392e+11Hz 0.459942 -0.871722
+ 1.393e+11Hz 0.459257 -0.872072
+ 1.394e+11Hz 0.45857 -0.872422
+ 1.395e+11Hz 0.457884 -0.87277
+ 1.396e+11Hz 0.457197 -0.873119
+ 1.397e+11Hz 0.45651 -0.873466
+ 1.398e+11Hz 0.455823 -0.873814
+ 1.399e+11Hz 0.455136 -0.87416
+ 1.4e+11Hz 0.454448 -0.874506
+ 1.401e+11Hz 0.45376 -0.874852
+ 1.402e+11Hz 0.453072 -0.875197
+ 1.403e+11Hz 0.452383 -0.875541
+ 1.404e+11Hz 0.451694 -0.875885
+ 1.405e+11Hz 0.451005 -0.876229
+ 1.406e+11Hz 0.450316 -0.876571
+ 1.407e+11Hz 0.449627 -0.876914
+ 1.408e+11Hz 0.448937 -0.877255
+ 1.409e+11Hz 0.448247 -0.877597
+ 1.41e+11Hz 0.447556 -0.877937
+ 1.411e+11Hz 0.446866 -0.878277
+ 1.412e+11Hz 0.446175 -0.878617
+ 1.413e+11Hz 0.445484 -0.878956
+ 1.414e+11Hz 0.444793 -0.879294
+ 1.415e+11Hz 0.444101 -0.879632
+ 1.416e+11Hz 0.443409 -0.879969
+ 1.417e+11Hz 0.442717 -0.880306
+ 1.418e+11Hz 0.442025 -0.880642
+ 1.419e+11Hz 0.441332 -0.880978
+ 1.42e+11Hz 0.440639 -0.881313
+ 1.421e+11Hz 0.439946 -0.881648
+ 1.422e+11Hz 0.439252 -0.881982
+ 1.423e+11Hz 0.438559 -0.882316
+ 1.424e+11Hz 0.437865 -0.882649
+ 1.425e+11Hz 0.437171 -0.882981
+ 1.426e+11Hz 0.436476 -0.883313
+ 1.427e+11Hz 0.435781 -0.883644
+ 1.428e+11Hz 0.435086 -0.883975
+ 1.429e+11Hz 0.434391 -0.884305
+ 1.43e+11Hz 0.433695 -0.884635
+ 1.431e+11Hz 0.433 -0.884964
+ 1.432e+11Hz 0.432304 -0.885293
+ 1.433e+11Hz 0.431607 -0.885621
+ 1.434e+11Hz 0.430911 -0.885948
+ 1.435e+11Hz 0.430214 -0.886275
+ 1.436e+11Hz 0.429517 -0.886602
+ 1.437e+11Hz 0.428819 -0.886927
+ 1.438e+11Hz 0.428121 -0.887253
+ 1.439e+11Hz 0.427423 -0.887578
+ 1.44e+11Hz 0.426725 -0.887902
+ 1.441e+11Hz 0.426027 -0.888225
+ 1.442e+11Hz 0.425328 -0.888548
+ 1.443e+11Hz 0.424629 -0.888871
+ 1.444e+11Hz 0.42393 -0.889193
+ 1.445e+11Hz 0.42323 -0.889514
+ 1.446e+11Hz 0.42253 -0.889835
+ 1.447e+11Hz 0.42183 -0.890156
+ 1.448e+11Hz 0.42113 -0.890476
+ 1.449e+11Hz 0.420429 -0.890795
+ 1.45e+11Hz 0.419728 -0.891113
+ 1.451e+11Hz 0.419027 -0.891432
+ 1.452e+11Hz 0.418325 -0.891749
+ 1.453e+11Hz 0.417623 -0.892066
+ 1.454e+11Hz 0.416921 -0.892382
+ 1.455e+11Hz 0.416219 -0.892698
+ 1.456e+11Hz 0.415517 -0.893014
+ 1.457e+11Hz 0.414814 -0.893328
+ 1.458e+11Hz 0.41411 -0.893643
+ 1.459e+11Hz 0.413407 -0.893956
+ 1.46e+11Hz 0.412703 -0.894269
+ 1.461e+11Hz 0.411999 -0.894582
+ 1.462e+11Hz 0.411295 -0.894894
+ 1.463e+11Hz 0.410591 -0.895205
+ 1.464e+11Hz 0.409886 -0.895516
+ 1.465e+11Hz 0.409181 -0.895826
+ 1.466e+11Hz 0.408475 -0.896136
+ 1.467e+11Hz 0.40777 -0.896445
+ 1.468e+11Hz 0.407064 -0.896753
+ 1.469e+11Hz 0.406358 -0.897061
+ 1.47e+11Hz 0.405651 -0.897368
+ 1.471e+11Hz 0.404944 -0.897675
+ 1.472e+11Hz 0.404237 -0.897981
+ 1.473e+11Hz 0.40353 -0.898287
+ 1.474e+11Hz 0.402823 -0.898592
+ 1.475e+11Hz 0.402115 -0.898896
+ 1.476e+11Hz 0.401407 -0.8992
+ 1.477e+11Hz 0.400698 -0.899503
+ 1.478e+11Hz 0.39999 -0.899806
+ 1.479e+11Hz 0.399281 -0.900108
+ 1.48e+11Hz 0.398572 -0.900409
+ 1.481e+11Hz 0.397862 -0.90071
+ 1.482e+11Hz 0.397152 -0.90101
+ 1.483e+11Hz 0.396442 -0.90131
+ 1.484e+11Hz 0.395732 -0.901609
+ 1.485e+11Hz 0.395021 -0.901908
+ 1.486e+11Hz 0.394311 -0.902205
+ 1.487e+11Hz 0.393599 -0.902503
+ 1.488e+11Hz 0.392888 -0.902799
+ 1.489e+11Hz 0.392176 -0.903095
+ 1.49e+11Hz 0.391465 -0.903391
+ 1.491e+11Hz 0.390752 -0.903686
+ 1.492e+11Hz 0.39004 -0.90398
+ 1.493e+11Hz 0.389327 -0.904274
+ 1.494e+11Hz 0.388614 -0.904567
+ 1.495e+11Hz 0.387901 -0.904859
+ 1.496e+11Hz 0.387187 -0.905151
+ 1.497e+11Hz 0.386474 -0.905442
+ 1.498e+11Hz 0.38576 -0.905733
+ 1.499e+11Hz 0.385045 -0.906023
+ 1.5e+11Hz 0.384331 -0.906312
+ 1.501e+11Hz 0.383616 -0.906601
+ 1.502e+11Hz 0.382901 -0.906889
+ 1.503e+11Hz 0.382186 -0.907176
+ 1.504e+11Hz 0.38147 -0.907463
+ 1.505e+11Hz 0.380754 -0.907749
+ 1.506e+11Hz 0.380038 -0.908035
+ 1.507e+11Hz 0.379322 -0.90832
+ 1.508e+11Hz 0.378605 -0.908604
+ 1.509e+11Hz 0.377888 -0.908888
+ 1.51e+11Hz 0.377171 -0.909171
+ 1.511e+11Hz 0.376454 -0.909453
+ 1.512e+11Hz 0.375736 -0.909735
+ 1.513e+11Hz 0.375018 -0.910016
+ 1.514e+11Hz 0.3743 -0.910297
+ 1.515e+11Hz 0.373582 -0.910577
+ 1.516e+11Hz 0.372863 -0.910856
+ 1.517e+11Hz 0.372145 -0.911135
+ 1.518e+11Hz 0.371426 -0.911413
+ 1.519e+11Hz 0.370706 -0.91169
+ 1.52e+11Hz 0.369987 -0.911967
+ 1.521e+11Hz 0.369267 -0.912243
+ 1.522e+11Hz 0.368547 -0.912518
+ 1.523e+11Hz 0.367827 -0.912793
+ 1.524e+11Hz 0.367107 -0.913067
+ 1.525e+11Hz 0.366386 -0.91334
+ 1.526e+11Hz 0.365665 -0.913613
+ 1.527e+11Hz 0.364944 -0.913885
+ 1.528e+11Hz 0.364223 -0.914157
+ 1.529e+11Hz 0.363501 -0.914428
+ 1.53e+11Hz 0.362779 -0.914698
+ 1.531e+11Hz 0.362057 -0.914967
+ 1.532e+11Hz 0.361335 -0.915236
+ 1.533e+11Hz 0.360613 -0.915504
+ 1.534e+11Hz 0.35989 -0.915772
+ 1.535e+11Hz 0.359167 -0.916039
+ 1.536e+11Hz 0.358444 -0.916305
+ 1.537e+11Hz 0.357721 -0.916571
+ 1.538e+11Hz 0.356997 -0.916836
+ 1.539e+11Hz 0.356274 -0.9171
+ 1.54e+11Hz 0.35555 -0.917364
+ 1.541e+11Hz 0.354826 -0.917627
+ 1.542e+11Hz 0.354102 -0.917889
+ 1.543e+11Hz 0.353377 -0.91815
+ 1.544e+11Hz 0.352652 -0.918411
+ 1.545e+11Hz 0.351928 -0.918672
+ 1.546e+11Hz 0.351203 -0.918931
+ 1.547e+11Hz 0.350477 -0.91919
+ 1.548e+11Hz 0.349752 -0.919449
+ 1.549e+11Hz 0.349026 -0.919706
+ 1.55e+11Hz 0.348301 -0.919963
+ 1.551e+11Hz 0.347575 -0.92022
+ 1.552e+11Hz 0.346849 -0.920475
+ 1.553e+11Hz 0.346122 -0.920731
+ 1.554e+11Hz 0.345396 -0.920985
+ 1.555e+11Hz 0.344669 -0.921239
+ 1.556e+11Hz 0.343942 -0.921492
+ 1.557e+11Hz 0.343215 -0.921744
+ 1.558e+11Hz 0.342488 -0.921996
+ 1.559e+11Hz 0.341761 -0.922247
+ 1.56e+11Hz 0.341033 -0.922497
+ 1.561e+11Hz 0.340306 -0.922747
+ 1.562e+11Hz 0.339578 -0.922996
+ 1.563e+11Hz 0.33885 -0.923244
+ 1.564e+11Hz 0.338122 -0.923492
+ 1.565e+11Hz 0.337393 -0.923739
+ 1.566e+11Hz 0.336665 -0.923985
+ 1.567e+11Hz 0.335936 -0.924231
+ 1.568e+11Hz 0.335207 -0.924476
+ 1.569e+11Hz 0.334479 -0.924721
+ 1.57e+11Hz 0.33375 -0.924964
+ 1.571e+11Hz 0.33302 -0.925207
+ 1.572e+11Hz 0.332291 -0.92545
+ 1.573e+11Hz 0.331561 -0.925692
+ 1.574e+11Hz 0.330832 -0.925933
+ 1.575e+11Hz 0.330102 -0.926173
+ 1.576e+11Hz 0.329372 -0.926413
+ 1.577e+11Hz 0.328642 -0.926652
+ 1.578e+11Hz 0.327912 -0.92689
+ 1.579e+11Hz 0.327182 -0.927128
+ 1.58e+11Hz 0.326451 -0.927365
+ 1.581e+11Hz 0.325721 -0.927602
+ 1.582e+11Hz 0.32499 -0.927838
+ 1.583e+11Hz 0.324259 -0.928073
+ 1.584e+11Hz 0.323528 -0.928307
+ 1.585e+11Hz 0.322797 -0.928541
+ 1.586e+11Hz 0.322066 -0.928774
+ 1.587e+11Hz 0.321335 -0.929007
+ 1.588e+11Hz 0.320603 -0.929239
+ 1.589e+11Hz 0.319872 -0.92947
+ 1.59e+11Hz 0.31914 -0.929701
+ 1.591e+11Hz 0.318408 -0.929931
+ 1.592e+11Hz 0.317676 -0.93016
+ 1.593e+11Hz 0.316944 -0.930389
+ 1.594e+11Hz 0.316212 -0.930617
+ 1.595e+11Hz 0.31548 -0.930844
+ 1.596e+11Hz 0.314747 -0.931071
+ 1.597e+11Hz 0.314015 -0.931297
+ 1.598e+11Hz 0.313282 -0.931522
+ 1.599e+11Hz 0.31255 -0.931747
+ 1.6e+11Hz 0.311817 -0.931971
+ 1.601e+11Hz 0.311084 -0.932194
+ 1.602e+11Hz 0.310351 -0.932417
+ 1.603e+11Hz 0.309618 -0.932639
+ 1.604e+11Hz 0.308885 -0.932861
+ 1.605e+11Hz 0.308152 -0.933082
+ 1.606e+11Hz 0.307418 -0.933302
+ 1.607e+11Hz 0.306685 -0.933522
+ 1.608e+11Hz 0.305951 -0.933741
+ 1.609e+11Hz 0.305217 -0.933959
+ 1.61e+11Hz 0.304484 -0.934177
+ 1.611e+11Hz 0.30375 -0.934394
+ 1.612e+11Hz 0.303016 -0.93461
+ 1.613e+11Hz 0.302282 -0.934826
+ 1.614e+11Hz 0.301548 -0.935041
+ 1.615e+11Hz 0.300813 -0.935256
+ 1.616e+11Hz 0.300079 -0.935469
+ 1.617e+11Hz 0.299345 -0.935683
+ 1.618e+11Hz 0.29861 -0.935895
+ 1.619e+11Hz 0.297876 -0.936107
+ 1.62e+11Hz 0.297141 -0.936319
+ 1.621e+11Hz 0.296406 -0.936529
+ 1.622e+11Hz 0.295671 -0.936739
+ 1.623e+11Hz 0.294937 -0.936949
+ 1.624e+11Hz 0.294202 -0.937158
+ 1.625e+11Hz 0.293466 -0.937366
+ 1.626e+11Hz 0.292731 -0.937574
+ 1.627e+11Hz 0.291996 -0.93778
+ 1.628e+11Hz 0.291261 -0.937987
+ 1.629e+11Hz 0.290525 -0.938193
+ 1.63e+11Hz 0.28979 -0.938398
+ 1.631e+11Hz 0.289054 -0.938602
+ 1.632e+11Hz 0.288319 -0.938806
+ 1.633e+11Hz 0.287583 -0.939009
+ 1.634e+11Hz 0.286847 -0.939212
+ 1.635e+11Hz 0.286111 -0.939414
+ 1.636e+11Hz 0.285375 -0.939615
+ 1.637e+11Hz 0.284639 -0.939816
+ 1.638e+11Hz 0.283903 -0.940016
+ 1.639e+11Hz 0.283167 -0.940215
+ 1.64e+11Hz 0.282431 -0.940414
+ 1.641e+11Hz 0.281694 -0.940612
+ 1.642e+11Hz 0.280958 -0.94081
+ 1.643e+11Hz 0.280221 -0.941007
+ 1.644e+11Hz 0.279485 -0.941203
+ 1.645e+11Hz 0.278748 -0.941399
+ 1.646e+11Hz 0.278012 -0.941594
+ 1.647e+11Hz 0.277275 -0.941789
+ 1.648e+11Hz 0.276538 -0.941983
+ 1.649e+11Hz 0.275801 -0.942176
+ 1.65e+11Hz 0.275064 -0.942369
+ 1.651e+11Hz 0.274327 -0.942561
+ 1.652e+11Hz 0.27359 -0.942752
+ 1.653e+11Hz 0.272853 -0.942943
+ 1.654e+11Hz 0.272116 -0.943133
+ 1.655e+11Hz 0.271378 -0.943323
+ 1.656e+11Hz 0.270641 -0.943512
+ 1.657e+11Hz 0.269903 -0.9437
+ 1.658e+11Hz 0.269166 -0.943888
+ 1.659e+11Hz 0.268428 -0.944075
+ 1.66e+11Hz 0.267691 -0.944262
+ 1.661e+11Hz 0.266953 -0.944448
+ 1.662e+11Hz 0.266215 -0.944633
+ 1.663e+11Hz 0.265478 -0.944818
+ 1.664e+11Hz 0.26474 -0.945002
+ 1.665e+11Hz 0.264002 -0.945185
+ 1.666e+11Hz 0.263264 -0.945368
+ 1.667e+11Hz 0.262526 -0.945551
+ 1.668e+11Hz 0.261788 -0.945732
+ 1.669e+11Hz 0.261049 -0.945913
+ 1.67e+11Hz 0.260311 -0.946094
+ 1.671e+11Hz 0.259573 -0.946273
+ 1.672e+11Hz 0.258834 -0.946453
+ 1.673e+11Hz 0.258096 -0.946631
+ 1.674e+11Hz 0.257358 -0.946809
+ 1.675e+11Hz 0.256619 -0.946987
+ 1.676e+11Hz 0.255881 -0.947163
+ 1.677e+11Hz 0.255142 -0.94734
+ 1.678e+11Hz 0.254403 -0.947515
+ 1.679e+11Hz 0.253665 -0.94769
+ 1.68e+11Hz 0.252926 -0.947864
+ 1.681e+11Hz 0.252187 -0.948038
+ 1.682e+11Hz 0.251448 -0.948211
+ 1.683e+11Hz 0.250709 -0.948384
+ 1.684e+11Hz 0.24997 -0.948556
+ 1.685e+11Hz 0.249231 -0.948727
+ 1.686e+11Hz 0.248492 -0.948898
+ 1.687e+11Hz 0.247753 -0.949068
+ 1.688e+11Hz 0.247014 -0.949237
+ 1.689e+11Hz 0.246275 -0.949406
+ 1.69e+11Hz 0.245535 -0.949574
+ 1.691e+11Hz 0.244796 -0.949742
+ 1.692e+11Hz 0.244057 -0.949909
+ 1.693e+11Hz 0.243317 -0.950075
+ 1.694e+11Hz 0.242578 -0.950241
+ 1.695e+11Hz 0.241839 -0.950406
+ 1.696e+11Hz 0.241099 -0.950571
+ 1.697e+11Hz 0.24036 -0.950735
+ 1.698e+11Hz 0.23962 -0.950898
+ 1.699e+11Hz 0.23888 -0.951061
+ 1.7e+11Hz 0.238141 -0.951223
+ 1.701e+11Hz 0.237401 -0.951384
+ 1.702e+11Hz 0.236662 -0.951545
+ 1.703e+11Hz 0.235922 -0.951706
+ 1.704e+11Hz 0.235182 -0.951865
+ 1.705e+11Hz 0.234442 -0.952024
+ 1.706e+11Hz 0.233703 -0.952183
+ 1.707e+11Hz 0.232963 -0.952341
+ 1.708e+11Hz 0.232223 -0.952498
+ 1.709e+11Hz 0.231483 -0.952655
+ 1.71e+11Hz 0.230743 -0.952811
+ 1.711e+11Hz 0.230003 -0.952966
+ 1.712e+11Hz 0.229263 -0.953121
+ 1.713e+11Hz 0.228523 -0.953275
+ 1.714e+11Hz 0.227783 -0.953429
+ 1.715e+11Hz 0.227043 -0.953582
+ 1.716e+11Hz 0.226303 -0.953735
+ 1.717e+11Hz 0.225563 -0.953886
+ 1.718e+11Hz 0.224823 -0.954038
+ 1.719e+11Hz 0.224083 -0.954188
+ 1.72e+11Hz 0.223343 -0.954338
+ 1.721e+11Hz 0.222603 -0.954488
+ 1.722e+11Hz 0.221863 -0.954637
+ 1.723e+11Hz 0.221123 -0.954785
+ 1.724e+11Hz 0.220383 -0.954933
+ 1.725e+11Hz 0.219643 -0.95508
+ 1.726e+11Hz 0.218903 -0.955226
+ 1.727e+11Hz 0.218163 -0.955372
+ 1.728e+11Hz 0.217423 -0.955517
+ 1.729e+11Hz 0.216683 -0.955662
+ 1.73e+11Hz 0.215943 -0.955806
+ 1.731e+11Hz 0.215203 -0.955949
+ 1.732e+11Hz 0.214463 -0.956092
+ 1.733e+11Hz 0.213723 -0.956234
+ 1.734e+11Hz 0.212983 -0.956376
+ 1.735e+11Hz 0.212243 -0.956517
+ 1.736e+11Hz 0.211503 -0.956658
+ 1.737e+11Hz 0.210763 -0.956798
+ 1.738e+11Hz 0.210023 -0.956937
+ 1.739e+11Hz 0.209283 -0.957076
+ 1.74e+11Hz 0.208543 -0.957214
+ 1.741e+11Hz 0.207803 -0.957352
+ 1.742e+11Hz 0.207063 -0.957489
+ 1.743e+11Hz 0.206323 -0.957625
+ 1.744e+11Hz 0.205583 -0.957761
+ 1.745e+11Hz 0.204844 -0.957896
+ 1.746e+11Hz 0.204104 -0.958031
+ 1.747e+11Hz 0.203364 -0.958165
+ 1.748e+11Hz 0.202624 -0.958298
+ 1.749e+11Hz 0.201884 -0.958431
+ 1.75e+11Hz 0.201145 -0.958564
+ 1.751e+11Hz 0.200405 -0.958696
+ 1.752e+11Hz 0.199665 -0.958827
+ 1.753e+11Hz 0.198926 -0.958957
+ 1.754e+11Hz 0.198186 -0.959088
+ 1.755e+11Hz 0.197447 -0.959217
+ 1.756e+11Hz 0.196707 -0.959346
+ 1.757e+11Hz 0.195968 -0.959474
+ 1.758e+11Hz 0.195228 -0.959602
+ 1.759e+11Hz 0.194489 -0.95973
+ 1.76e+11Hz 0.19375 -0.959856
+ 1.761e+11Hz 0.19301 -0.959983
+ 1.762e+11Hz 0.192271 -0.960108
+ 1.763e+11Hz 0.191532 -0.960233
+ 1.764e+11Hz 0.190792 -0.960358
+ 1.765e+11Hz 0.190053 -0.960482
+ 1.766e+11Hz 0.189314 -0.960605
+ 1.767e+11Hz 0.188575 -0.960728
+ 1.768e+11Hz 0.187836 -0.96085
+ 1.769e+11Hz 0.187097 -0.960972
+ 1.77e+11Hz 0.186358 -0.961093
+ 1.771e+11Hz 0.185619 -0.961214
+ 1.772e+11Hz 0.18488 -0.961334
+ 1.773e+11Hz 0.184142 -0.961454
+ 1.774e+11Hz 0.183403 -0.961573
+ 1.775e+11Hz 0.182664 -0.961692
+ 1.776e+11Hz 0.181926 -0.96181
+ 1.777e+11Hz 0.181187 -0.961927
+ 1.778e+11Hz 0.180448 -0.962044
+ 1.779e+11Hz 0.17971 -0.962161
+ 1.78e+11Hz 0.178971 -0.962277
+ 1.781e+11Hz 0.178233 -0.962392
+ 1.782e+11Hz 0.177495 -0.962507
+ 1.783e+11Hz 0.176756 -0.962622
+ 1.784e+11Hz 0.176018 -0.962735
+ 1.785e+11Hz 0.17528 -0.962849
+ 1.786e+11Hz 0.174542 -0.962962
+ 1.787e+11Hz 0.173804 -0.963074
+ 1.788e+11Hz 0.173066 -0.963186
+ 1.789e+11Hz 0.172328 -0.963297
+ 1.79e+11Hz 0.17159 -0.963408
+ 1.791e+11Hz 0.170852 -0.963518
+ 1.792e+11Hz 0.170114 -0.963628
+ 1.793e+11Hz 0.169376 -0.963738
+ 1.794e+11Hz 0.168638 -0.963847
+ 1.795e+11Hz 0.167901 -0.963955
+ 1.796e+11Hz 0.167163 -0.964063
+ 1.797e+11Hz 0.166425 -0.96417
+ 1.798e+11Hz 0.165688 -0.964277
+ 1.799e+11Hz 0.16495 -0.964384
+ 1.8e+11Hz 0.164213 -0.96449
+ 1.801e+11Hz 0.163475 -0.964595
+ 1.802e+11Hz 0.162738 -0.9647
+ 1.803e+11Hz 0.162001 -0.964805
+ 1.804e+11Hz 0.161263 -0.964909
+ 1.805e+11Hz 0.160526 -0.965012
+ 1.806e+11Hz 0.159789 -0.965115
+ 1.807e+11Hz 0.159052 -0.965218
+ 1.808e+11Hz 0.158314 -0.96532
+ 1.809e+11Hz 0.157577 -0.965422
+ 1.81e+11Hz 0.15684 -0.965523
+ 1.811e+11Hz 0.156103 -0.965624
+ 1.812e+11Hz 0.155366 -0.965724
+ 1.813e+11Hz 0.154629 -0.965824
+ 1.814e+11Hz 0.153892 -0.965923
+ 1.815e+11Hz 0.153155 -0.966022
+ 1.816e+11Hz 0.152418 -0.966121
+ 1.817e+11Hz 0.151682 -0.966219
+ 1.818e+11Hz 0.150945 -0.966317
+ 1.819e+11Hz 0.150208 -0.966414
+ 1.82e+11Hz 0.149471 -0.96651
+ 1.821e+11Hz 0.148734 -0.966607
+ 1.822e+11Hz 0.147998 -0.966703
+ 1.823e+11Hz 0.147261 -0.966798
+ 1.824e+11Hz 0.146524 -0.966893
+ 1.825e+11Hz 0.145787 -0.966987
+ 1.826e+11Hz 0.145051 -0.967081
+ 1.827e+11Hz 0.144314 -0.967175
+ 1.828e+11Hz 0.143577 -0.967268
+ 1.829e+11Hz 0.142841 -0.967361
+ 1.83e+11Hz 0.142104 -0.967453
+ 1.831e+11Hz 0.141367 -0.967545
+ 1.832e+11Hz 0.140631 -0.967637
+ 1.833e+11Hz 0.139894 -0.967728
+ 1.834e+11Hz 0.139158 -0.967818
+ 1.835e+11Hz 0.138421 -0.967908
+ 1.836e+11Hz 0.137684 -0.967998
+ 1.837e+11Hz 0.136948 -0.968088
+ 1.838e+11Hz 0.136211 -0.968176
+ 1.839e+11Hz 0.135474 -0.968265
+ 1.84e+11Hz 0.134738 -0.968353
+ 1.841e+11Hz 0.134001 -0.968441
+ 1.842e+11Hz 0.133264 -0.968528
+ 1.843e+11Hz 0.132527 -0.968615
+ 1.844e+11Hz 0.131791 -0.968701
+ 1.845e+11Hz 0.131054 -0.968787
+ 1.846e+11Hz 0.130317 -0.968872
+ 1.847e+11Hz 0.12958 -0.968957
+ 1.848e+11Hz 0.128843 -0.969042
+ 1.849e+11Hz 0.128106 -0.969126
+ 1.85e+11Hz 0.127369 -0.96921
+ 1.851e+11Hz 0.126632 -0.969293
+ 1.852e+11Hz 0.125895 -0.969376
+ 1.853e+11Hz 0.125158 -0.969459
+ 1.854e+11Hz 0.124421 -0.969541
+ 1.855e+11Hz 0.123684 -0.969623
+ 1.856e+11Hz 0.122947 -0.969704
+ 1.857e+11Hz 0.12221 -0.969785
+ 1.858e+11Hz 0.121472 -0.969866
+ 1.859e+11Hz 0.120735 -0.969946
+ 1.86e+11Hz 0.119998 -0.970025
+ 1.861e+11Hz 0.11926 -0.970104
+ 1.862e+11Hz 0.118523 -0.970183
+ 1.863e+11Hz 0.117785 -0.970261
+ 1.864e+11Hz 0.117047 -0.970339
+ 1.865e+11Hz 0.11631 -0.970417
+ 1.866e+11Hz 0.115572 -0.970494
+ 1.867e+11Hz 0.114834 -0.970571
+ 1.868e+11Hz 0.114096 -0.970647
+ 1.869e+11Hz 0.113358 -0.970723
+ 1.87e+11Hz 0.11262 -0.970798
+ 1.871e+11Hz 0.111882 -0.970873
+ 1.872e+11Hz 0.111144 -0.970947
+ 1.873e+11Hz 0.110405 -0.971021
+ 1.874e+11Hz 0.109667 -0.971095
+ 1.875e+11Hz 0.108928 -0.971168
+ 1.876e+11Hz 0.10819 -0.971241
+ 1.877e+11Hz 0.107451 -0.971313
+ 1.878e+11Hz 0.106712 -0.971385
+ 1.879e+11Hz 0.105973 -0.971457
+ 1.88e+11Hz 0.105234 -0.971528
+ 1.881e+11Hz 0.104495 -0.971598
+ 1.882e+11Hz 0.103756 -0.971668
+ 1.883e+11Hz 0.103017 -0.971738
+ 1.884e+11Hz 0.102277 -0.971807
+ 1.885e+11Hz 0.101538 -0.971876
+ 1.886e+11Hz 0.100798 -0.971944
+ 1.887e+11Hz 0.100059 -0.972012
+ 1.888e+11Hz 0.0993189 -0.972079
+ 1.889e+11Hz 0.098579 -0.972146
+ 1.89e+11Hz 0.097839 -0.972213
+ 1.891e+11Hz 0.0970988 -0.972279
+ 1.892e+11Hz 0.0963586 -0.972344
+ 1.893e+11Hz 0.0956182 -0.97241
+ 1.894e+11Hz 0.0948777 -0.972474
+ 1.895e+11Hz 0.0941371 -0.972538
+ 1.896e+11Hz 0.0933963 -0.972602
+ 1.897e+11Hz 0.0926555 -0.972665
+ 1.898e+11Hz 0.0919145 -0.972728
+ 1.899e+11Hz 0.0911734 -0.97279
+ 1.9e+11Hz 0.0904321 -0.972852
+ 1.901e+11Hz 0.0896908 -0.972914
+ 1.902e+11Hz 0.0889493 -0.972974
+ 1.903e+11Hz 0.0882077 -0.973035
+ 1.904e+11Hz 0.0874659 -0.973095
+ 1.905e+11Hz 0.0867241 -0.973154
+ 1.906e+11Hz 0.0859821 -0.973213
+ 1.907e+11Hz 0.0852399 -0.973271
+ 1.908e+11Hz 0.0844977 -0.973329
+ 1.909e+11Hz 0.0837553 -0.973387
+ 1.91e+11Hz 0.0830128 -0.973444
+ 1.911e+11Hz 0.0822701 -0.9735
+ 1.912e+11Hz 0.0815273 -0.973556
+ 1.913e+11Hz 0.0807844 -0.973611
+ 1.914e+11Hz 0.0800413 -0.973666
+ 1.915e+11Hz 0.0792981 -0.97372
+ 1.916e+11Hz 0.0785548 -0.973774
+ 1.917e+11Hz 0.0778114 -0.973828
+ 1.918e+11Hz 0.0770678 -0.97388
+ 1.919e+11Hz 0.076324 -0.973933
+ 1.92e+11Hz 0.0755802 -0.973985
+ 1.921e+11Hz 0.0748362 -0.974036
+ 1.922e+11Hz 0.074092 -0.974086
+ 1.923e+11Hz 0.0733478 -0.974137
+ 1.924e+11Hz 0.0726034 -0.974186
+ 1.925e+11Hz 0.0718589 -0.974235
+ 1.926e+11Hz 0.0711142 -0.974284
+ 1.927e+11Hz 0.0703694 -0.974332
+ 1.928e+11Hz 0.0696245 -0.974379
+ 1.929e+11Hz 0.0688794 -0.974426
+ 1.93e+11Hz 0.0681342 -0.974473
+ 1.931e+11Hz 0.0673889 -0.974519
+ 1.932e+11Hz 0.0666435 -0.974564
+ 1.933e+11Hz 0.0658979 -0.974609
+ 1.934e+11Hz 0.0651522 -0.974653
+ 1.935e+11Hz 0.0644063 -0.974696
+ 1.936e+11Hz 0.0636604 -0.974739
+ 1.937e+11Hz 0.0629143 -0.974782
+ 1.938e+11Hz 0.0621681 -0.974824
+ 1.939e+11Hz 0.0614217 -0.974865
+ 1.94e+11Hz 0.0606753 -0.974906
+ 1.941e+11Hz 0.0599287 -0.974946
+ 1.942e+11Hz 0.059182 -0.974985
+ 1.943e+11Hz 0.0584352 -0.975025
+ 1.944e+11Hz 0.0576883 -0.975063
+ 1.945e+11Hz 0.0569412 -0.975101
+ 1.946e+11Hz 0.056194 -0.975138
+ 1.947e+11Hz 0.0554468 -0.975175
+ 1.948e+11Hz 0.0546994 -0.975211
+ 1.949e+11Hz 0.0539519 -0.975246
+ 1.95e+11Hz 0.0532043 -0.975281
+ 1.951e+11Hz 0.0524565 -0.975316
+ 1.952e+11Hz 0.0517087 -0.975349
+ 1.953e+11Hz 0.0509608 -0.975382
+ 1.954e+11Hz 0.0502128 -0.975415
+ 1.955e+11Hz 0.0494646 -0.975447
+ 1.956e+11Hz 0.0487164 -0.975478
+ 1.957e+11Hz 0.0479681 -0.975509
+ 1.958e+11Hz 0.0472196 -0.975539
+ 1.959e+11Hz 0.0464711 -0.975568
+ 1.96e+11Hz 0.0457225 -0.975597
+ 1.961e+11Hz 0.0449738 -0.975625
+ 1.962e+11Hz 0.044225 -0.975653
+ 1.963e+11Hz 0.0434761 -0.97568
+ 1.964e+11Hz 0.0427272 -0.975706
+ 1.965e+11Hz 0.0419781 -0.975732
+ 1.966e+11Hz 0.041229 -0.975757
+ 1.967e+11Hz 0.0404798 -0.975782
+ 1.968e+11Hz 0.0397305 -0.975806
+ 1.969e+11Hz 0.0389812 -0.975829
+ 1.97e+11Hz 0.0382317 -0.975852
+ 1.971e+11Hz 0.0374822 -0.975874
+ 1.972e+11Hz 0.0367327 -0.975895
+ 1.973e+11Hz 0.035983 -0.975916
+ 1.974e+11Hz 0.0352333 -0.975936
+ 1.975e+11Hz 0.0344836 -0.975955
+ 1.976e+11Hz 0.0337338 -0.975974
+ 1.977e+11Hz 0.0329839 -0.975992
+ 1.978e+11Hz 0.032234 -0.97601
+ 1.979e+11Hz 0.031484 -0.976027
+ 1.98e+11Hz 0.0307339 -0.976043
+ 1.981e+11Hz 0.0299839 -0.976059
+ 1.982e+11Hz 0.0292337 -0.976074
+ 1.983e+11Hz 0.0284836 -0.976088
+ 1.984e+11Hz 0.0277334 -0.976102
+ 1.985e+11Hz 0.0269831 -0.976115
+ 1.986e+11Hz 0.0262328 -0.976128
+ 1.987e+11Hz 0.0254825 -0.97614
+ 1.988e+11Hz 0.0247321 -0.976151
+ 1.989e+11Hz 0.0239817 -0.976161
+ 1.99e+11Hz 0.0232313 -0.976171
+ 1.991e+11Hz 0.0224809 -0.976181
+ 1.992e+11Hz 0.0217304 -0.976189
+ 1.993e+11Hz 0.0209799 -0.976197
+ 1.994e+11Hz 0.0202294 -0.976205
+ 1.995e+11Hz 0.0194789 -0.976211
+ 1.996e+11Hz 0.0187284 -0.976217
+ 1.997e+11Hz 0.0179778 -0.976223
+ 1.998e+11Hz 0.0172273 -0.976227
+ 1.999e+11Hz 0.0164767 -0.976232
+ 2e+11Hz 0.0157261 -0.976235
+ 2.001e+11Hz 0.0149755 -0.976238
+ 2.002e+11Hz 0.014225 -0.97624
+ 2.003e+11Hz 0.0134744 -0.976242
+ 2.004e+11Hz 0.0127238 -0.976242
+ 2.005e+11Hz 0.0119732 -0.976243
+ 2.006e+11Hz 0.0112227 -0.976242
+ 2.007e+11Hz 0.0104721 -0.976241
+ 2.008e+11Hz 0.00972156 -0.97624
+ 2.009e+11Hz 0.00897103 -0.976237
+ 2.01e+11Hz 0.00822051 -0.976234
+ 2.011e+11Hz 0.00747001 -0.976231
+ 2.012e+11Hz 0.00671953 -0.976226
+ 2.013e+11Hz 0.00596907 -0.976222
+ 2.014e+11Hz 0.00521864 -0.976216
+ 2.015e+11Hz 0.00446823 -0.97621
+ 2.016e+11Hz 0.00371784 -0.976203
+ 2.017e+11Hz 0.00296749 -0.976196
+ 2.018e+11Hz 0.00221717 -0.976187
+ 2.019e+11Hz 0.00146688 -0.976179
+ 2.02e+11Hz 0.00071662 -0.976169
+ 2.021e+11Hz -3.35995e-05 -0.976159
+ 2.022e+11Hz -0.00078378 -0.976149
+ 2.023e+11Hz -0.00153392 -0.976137
+ 2.024e+11Hz -0.00228402 -0.976125
+ 2.025e+11Hz -0.00303408 -0.976113
+ 2.026e+11Hz -0.00378409 -0.9761
+ 2.027e+11Hz -0.00453405 -0.976086
+ 2.028e+11Hz -0.00528396 -0.976071
+ 2.029e+11Hz -0.00603383 -0.976056
+ 2.03e+11Hz -0.00678364 -0.97604
+ 2.031e+11Hz -0.0075334 -0.976024
+ 2.032e+11Hz -0.0082831 -0.976007
+ 2.033e+11Hz -0.00903275 -0.975989
+ 2.034e+11Hz -0.00978234 -0.975971
+ 2.035e+11Hz -0.0105319 -0.975952
+ 2.036e+11Hz -0.0112813 -0.975933
+ 2.037e+11Hz -0.0120307 -0.975913
+ 2.038e+11Hz -0.0127801 -0.975892
+ 2.039e+11Hz -0.0135294 -0.97587
+ 2.04e+11Hz -0.0142786 -0.975848
+ 2.041e+11Hz -0.0150277 -0.975826
+ 2.042e+11Hz -0.0157768 -0.975802
+ 2.043e+11Hz -0.0165258 -0.975779
+ 2.044e+11Hz -0.0172747 -0.975754
+ 2.045e+11Hz -0.0180236 -0.975729
+ 2.046e+11Hz -0.0187723 -0.975703
+ 2.047e+11Hz -0.019521 -0.975677
+ 2.048e+11Hz -0.0202697 -0.97565
+ 2.049e+11Hz -0.0210182 -0.975622
+ 2.05e+11Hz -0.0217667 -0.975594
+ 2.051e+11Hz -0.0225151 -0.975565
+ 2.052e+11Hz -0.0232634 -0.975536
+ 2.053e+11Hz -0.0240116 -0.975506
+ 2.054e+11Hz -0.0247597 -0.975475
+ 2.055e+11Hz -0.0255078 -0.975444
+ 2.056e+11Hz -0.0262557 -0.975412
+ 2.057e+11Hz -0.0270036 -0.975379
+ 2.058e+11Hz -0.0277514 -0.975346
+ 2.059e+11Hz -0.0284991 -0.975312
+ 2.06e+11Hz -0.0292467 -0.975278
+ 2.061e+11Hz -0.0299942 -0.975243
+ 2.062e+11Hz -0.0307416 -0.975208
+ 2.063e+11Hz -0.0314889 -0.975171
+ 2.064e+11Hz -0.0322361 -0.975135
+ 2.065e+11Hz -0.0329833 -0.975097
+ 2.066e+11Hz -0.0337303 -0.975059
+ 2.067e+11Hz -0.0344772 -0.975021
+ 2.068e+11Hz -0.0352241 -0.974982
+ 2.069e+11Hz -0.0359708 -0.974942
+ 2.07e+11Hz -0.0367175 -0.974901
+ 2.071e+11Hz -0.037464 -0.97486
+ 2.072e+11Hz -0.0382104 -0.974819
+ 2.073e+11Hz -0.0389567 -0.974777
+ 2.074e+11Hz -0.039703 -0.974734
+ 2.075e+11Hz -0.0404491 -0.974691
+ 2.076e+11Hz -0.0411951 -0.974647
+ 2.077e+11Hz -0.041941 -0.974602
+ 2.078e+11Hz -0.0426868 -0.974557
+ 2.079e+11Hz -0.0434324 -0.974511
+ 2.08e+11Hz -0.044178 -0.974465
+ 2.081e+11Hz -0.0449235 -0.974418
+ 2.082e+11Hz -0.0456688 -0.97437
+ 2.083e+11Hz -0.046414 -0.974322
+ 2.084e+11Hz -0.0471591 -0.974274
+ 2.085e+11Hz -0.0479041 -0.974224
+ 2.086e+11Hz -0.048649 -0.974174
+ 2.087e+11Hz -0.0493938 -0.974124
+ 2.088e+11Hz -0.0501384 -0.974073
+ 2.089e+11Hz -0.050883 -0.974021
+ 2.09e+11Hz -0.0516274 -0.973969
+ 2.091e+11Hz -0.0523716 -0.973916
+ 2.092e+11Hz -0.0531158 -0.973863
+ 2.093e+11Hz -0.0538598 -0.973809
+ 2.094e+11Hz -0.0546038 -0.973754
+ 2.095e+11Hz -0.0553475 -0.973699
+ 2.096e+11Hz -0.0560912 -0.973644
+ 2.097e+11Hz -0.0568347 -0.973587
+ 2.098e+11Hz -0.0575781 -0.97353
+ 2.099e+11Hz -0.0583214 -0.973473
+ 2.1e+11Hz -0.0590646 -0.973415
+ 2.101e+11Hz -0.0598076 -0.973356
+ 2.102e+11Hz -0.0605504 -0.973297
+ 2.103e+11Hz -0.0612932 -0.973237
+ 2.104e+11Hz -0.0620358 -0.973177
+ 2.105e+11Hz -0.0627783 -0.973116
+ 2.106e+11Hz -0.0635206 -0.973055
+ 2.107e+11Hz -0.0642628 -0.972992
+ 2.108e+11Hz -0.0650049 -0.97293
+ 2.109e+11Hz -0.0657468 -0.972867
+ 2.11e+11Hz -0.0664885 -0.972803
+ 2.111e+11Hz -0.0672302 -0.972739
+ 2.112e+11Hz -0.0679717 -0.972674
+ 2.113e+11Hz -0.068713 -0.972608
+ 2.114e+11Hz -0.0694542 -0.972542
+ 2.115e+11Hz -0.0701952 -0.972475
+ 2.116e+11Hz -0.0709361 -0.972408
+ 2.117e+11Hz -0.0716769 -0.97234
+ 2.118e+11Hz -0.0724175 -0.972272
+ 2.119e+11Hz -0.0731579 -0.972203
+ 2.12e+11Hz -0.0738982 -0.972134
+ 2.121e+11Hz -0.0746383 -0.972064
+ 2.122e+11Hz -0.0753783 -0.971993
+ 2.123e+11Hz -0.0761181 -0.971922
+ 2.124e+11Hz -0.0768577 -0.97185
+ 2.125e+11Hz -0.0775972 -0.971778
+ 2.126e+11Hz -0.0783366 -0.971705
+ 2.127e+11Hz -0.0790757 -0.971632
+ 2.128e+11Hz -0.0798147 -0.971558
+ 2.129e+11Hz -0.0805536 -0.971484
+ 2.13e+11Hz -0.0812922 -0.971409
+ 2.131e+11Hz -0.0820307 -0.971333
+ 2.132e+11Hz -0.0827691 -0.971257
+ 2.133e+11Hz -0.0835072 -0.97118
+ 2.134e+11Hz -0.0842452 -0.971103
+ 2.135e+11Hz -0.084983 -0.971026
+ 2.136e+11Hz -0.0857206 -0.970947
+ 2.137e+11Hz -0.0864581 -0.970868
+ 2.138e+11Hz -0.0871954 -0.970789
+ 2.139e+11Hz -0.0879325 -0.970709
+ 2.14e+11Hz -0.0886694 -0.970629
+ 2.141e+11Hz -0.0894061 -0.970548
+ 2.142e+11Hz -0.0901427 -0.970466
+ 2.143e+11Hz -0.090879 -0.970384
+ 2.144e+11Hz -0.0916152 -0.970302
+ 2.145e+11Hz -0.0923512 -0.970219
+ 2.146e+11Hz -0.093087 -0.970135
+ 2.147e+11Hz -0.0938226 -0.970051
+ 2.148e+11Hz -0.0945581 -0.969966
+ 2.149e+11Hz -0.0952933 -0.969881
+ 2.15e+11Hz -0.0960283 -0.969795
+ 2.151e+11Hz -0.0967632 -0.969709
+ 2.152e+11Hz -0.0974978 -0.969622
+ 2.153e+11Hz -0.0982323 -0.969535
+ 2.154e+11Hz -0.0989665 -0.969447
+ 2.155e+11Hz -0.0997006 -0.969359
+ 2.156e+11Hz -0.100434 -0.96927
+ 2.157e+11Hz -0.101168 -0.969181
+ 2.158e+11Hz -0.101902 -0.969091
+ 2.159e+11Hz -0.102635 -0.969001
+ 2.16e+11Hz -0.103368 -0.96891
+ 2.161e+11Hz -0.104101 -0.968819
+ 2.162e+11Hz -0.104833 -0.968727
+ 2.163e+11Hz -0.105566 -0.968635
+ 2.164e+11Hz -0.106298 -0.968542
+ 2.165e+11Hz -0.10703 -0.968449
+ 2.166e+11Hz -0.107762 -0.968355
+ 2.167e+11Hz -0.108493 -0.968261
+ 2.168e+11Hz -0.109225 -0.968166
+ 2.169e+11Hz -0.109956 -0.968071
+ 2.17e+11Hz -0.110687 -0.967976
+ 2.171e+11Hz -0.111418 -0.96788
+ 2.172e+11Hz -0.112148 -0.967783
+ 2.173e+11Hz -0.112878 -0.967686
+ 2.174e+11Hz -0.113608 -0.967589
+ 2.175e+11Hz -0.114338 -0.967491
+ 2.176e+11Hz -0.115068 -0.967392
+ 2.177e+11Hz -0.115797 -0.967294
+ 2.178e+11Hz -0.116527 -0.967194
+ 2.179e+11Hz -0.117256 -0.967095
+ 2.18e+11Hz -0.117984 -0.966995
+ 2.181e+11Hz -0.118713 -0.966894
+ 2.182e+11Hz -0.119441 -0.966793
+ 2.183e+11Hz -0.12017 -0.966691
+ 2.184e+11Hz -0.120898 -0.96659
+ 2.185e+11Hz -0.121625 -0.966487
+ 2.186e+11Hz -0.122353 -0.966385
+ 2.187e+11Hz -0.12308 -0.966281
+ 2.188e+11Hz -0.123807 -0.966178
+ 2.189e+11Hz -0.124534 -0.966074
+ 2.19e+11Hz -0.125261 -0.96597
+ 2.191e+11Hz -0.125987 -0.965865
+ 2.192e+11Hz -0.126713 -0.96576
+ 2.193e+11Hz -0.127439 -0.965654
+ 2.194e+11Hz -0.128165 -0.965548
+ 2.195e+11Hz -0.128891 -0.965442
+ 2.196e+11Hz -0.129616 -0.965335
+ 2.197e+11Hz -0.130341 -0.965228
+ 2.198e+11Hz -0.131066 -0.96512
+ 2.199e+11Hz -0.131791 -0.965012
+ 2.2e+11Hz -0.132516 -0.964904
+ 2.201e+11Hz -0.13324 -0.964795
+ 2.202e+11Hz -0.133964 -0.964686
+ 2.203e+11Hz -0.134688 -0.964577
+ 2.204e+11Hz -0.135412 -0.964467
+ 2.205e+11Hz -0.136136 -0.964357
+ 2.206e+11Hz -0.136859 -0.964247
+ 2.207e+11Hz -0.137582 -0.964136
+ 2.208e+11Hz -0.138305 -0.964025
+ 2.209e+11Hz -0.139028 -0.963913
+ 2.21e+11Hz -0.139751 -0.963801
+ 2.211e+11Hz -0.140473 -0.963689
+ 2.212e+11Hz -0.141195 -0.963576
+ 2.213e+11Hz -0.141917 -0.963464
+ 2.214e+11Hz -0.142639 -0.96335
+ 2.215e+11Hz -0.143361 -0.963237
+ 2.216e+11Hz -0.144083 -0.963123
+ 2.217e+11Hz -0.144804 -0.963009
+ 2.218e+11Hz -0.145525 -0.962894
+ 2.219e+11Hz -0.146246 -0.96278
+ 2.22e+11Hz -0.146967 -0.962665
+ 2.221e+11Hz -0.147688 -0.962549
+ 2.222e+11Hz -0.148409 -0.962433
+ 2.223e+11Hz -0.149129 -0.962317
+ 2.224e+11Hz -0.149849 -0.962201
+ 2.225e+11Hz -0.15057 -0.962085
+ 2.226e+11Hz -0.15129 -0.961968
+ 2.227e+11Hz -0.152009 -0.96185
+ 2.228e+11Hz -0.152729 -0.961733
+ 2.229e+11Hz -0.153449 -0.961615
+ 2.23e+11Hz -0.154168 -0.961497
+ 2.231e+11Hz -0.154888 -0.961379
+ 2.232e+11Hz -0.155607 -0.96126
+ 2.233e+11Hz -0.156326 -0.961141
+ 2.234e+11Hz -0.157045 -0.961022
+ 2.235e+11Hz -0.157764 -0.960903
+ 2.236e+11Hz -0.158483 -0.960783
+ 2.237e+11Hz -0.159202 -0.960663
+ 2.238e+11Hz -0.15992 -0.960543
+ 2.239e+11Hz -0.160639 -0.960422
+ 2.24e+11Hz -0.161357 -0.960302
+ 2.241e+11Hz -0.162076 -0.960181
+ 2.242e+11Hz -0.162794 -0.960059
+ 2.243e+11Hz -0.163512 -0.959938
+ 2.244e+11Hz -0.16423 -0.959816
+ 2.245e+11Hz -0.164948 -0.959694
+ 2.246e+11Hz -0.165667 -0.959572
+ 2.247e+11Hz -0.166385 -0.959449
+ 2.248e+11Hz -0.167102 -0.959326
+ 2.249e+11Hz -0.16782 -0.959203
+ 2.25e+11Hz -0.168538 -0.95908
+ 2.251e+11Hz -0.169256 -0.958956
+ 2.252e+11Hz -0.169974 -0.958832
+ 2.253e+11Hz -0.170692 -0.958708
+ 2.254e+11Hz -0.17141 -0.958584
+ 2.255e+11Hz -0.172127 -0.958459
+ 2.256e+11Hz -0.172845 -0.958335
+ 2.257e+11Hz -0.173563 -0.95821
+ 2.258e+11Hz -0.174281 -0.958084
+ 2.259e+11Hz -0.174999 -0.957959
+ 2.26e+11Hz -0.175716 -0.957833
+ 2.261e+11Hz -0.176434 -0.957707
+ 2.262e+11Hz -0.177152 -0.95758
+ 2.263e+11Hz -0.17787 -0.957454
+ 2.264e+11Hz -0.178588 -0.957327
+ 2.265e+11Hz -0.179306 -0.9572
+ 2.266e+11Hz -0.180024 -0.957073
+ 2.267e+11Hz -0.180742 -0.956945
+ 2.268e+11Hz -0.18146 -0.956817
+ 2.269e+11Hz -0.182178 -0.956689
+ 2.27e+11Hz -0.182897 -0.956561
+ 2.271e+11Hz -0.183615 -0.956432
+ 2.272e+11Hz -0.184333 -0.956303
+ 2.273e+11Hz -0.185052 -0.956174
+ 2.274e+11Hz -0.18577 -0.956044
+ 2.275e+11Hz -0.186489 -0.955915
+ 2.276e+11Hz -0.187208 -0.955785
+ 2.277e+11Hz -0.187927 -0.955655
+ 2.278e+11Hz -0.188646 -0.955524
+ 2.279e+11Hz -0.189365 -0.955393
+ 2.28e+11Hz -0.190084 -0.955262
+ 2.281e+11Hz -0.190804 -0.955131
+ 2.282e+11Hz -0.191523 -0.954999
+ 2.283e+11Hz -0.192243 -0.954867
+ 2.284e+11Hz -0.192963 -0.954735
+ 2.285e+11Hz -0.193683 -0.954602
+ 2.286e+11Hz -0.194403 -0.954469
+ 2.287e+11Hz -0.195123 -0.954336
+ 2.288e+11Hz -0.195844 -0.954203
+ 2.289e+11Hz -0.196564 -0.954069
+ 2.29e+11Hz -0.197285 -0.953935
+ 2.291e+11Hz -0.198006 -0.9538
+ 2.292e+11Hz -0.198727 -0.953665
+ 2.293e+11Hz -0.199449 -0.95353
+ 2.294e+11Hz -0.20017 -0.953395
+ 2.295e+11Hz -0.200892 -0.953259
+ 2.296e+11Hz -0.201614 -0.953123
+ 2.297e+11Hz -0.202336 -0.952986
+ 2.298e+11Hz -0.203058 -0.952849
+ 2.299e+11Hz -0.203781 -0.952712
+ 2.3e+11Hz -0.204504 -0.952575
+ 2.301e+11Hz -0.205227 -0.952437
+ 2.302e+11Hz -0.20595 -0.952298
+ 2.303e+11Hz -0.206673 -0.952159
+ 2.304e+11Hz -0.207397 -0.95202
+ 2.305e+11Hz -0.208121 -0.951881
+ 2.306e+11Hz -0.208845 -0.951741
+ 2.307e+11Hz -0.209569 -0.951601
+ 2.308e+11Hz -0.210294 -0.95146
+ 2.309e+11Hz -0.211019 -0.951319
+ 2.31e+11Hz -0.211744 -0.951177
+ 2.311e+11Hz -0.212469 -0.951035
+ 2.312e+11Hz -0.213195 -0.950893
+ 2.313e+11Hz -0.213921 -0.95075
+ 2.314e+11Hz -0.214647 -0.950606
+ 2.315e+11Hz -0.215374 -0.950462
+ 2.316e+11Hz -0.2161 -0.950318
+ 2.317e+11Hz -0.216827 -0.950173
+ 2.318e+11Hz -0.217554 -0.950028
+ 2.319e+11Hz -0.218282 -0.949883
+ 2.32e+11Hz -0.21901 -0.949736
+ 2.321e+11Hz -0.219738 -0.94959
+ 2.322e+11Hz -0.220466 -0.949442
+ 2.323e+11Hz -0.221195 -0.949295
+ 2.324e+11Hz -0.221923 -0.949146
+ 2.325e+11Hz -0.222653 -0.948998
+ 2.326e+11Hz -0.223382 -0.948848
+ 2.327e+11Hz -0.224112 -0.948699
+ 2.328e+11Hz -0.224842 -0.948548
+ 2.329e+11Hz -0.225572 -0.948397
+ 2.33e+11Hz -0.226302 -0.948246
+ 2.331e+11Hz -0.227033 -0.948094
+ 2.332e+11Hz -0.227764 -0.947941
+ 2.333e+11Hz -0.228495 -0.947788
+ 2.334e+11Hz -0.229227 -0.947634
+ 2.335e+11Hz -0.229959 -0.947479
+ 2.336e+11Hz -0.230691 -0.947324
+ 2.337e+11Hz -0.231424 -0.947169
+ 2.338e+11Hz -0.232156 -0.947012
+ 2.339e+11Hz -0.232889 -0.946855
+ 2.34e+11Hz -0.233623 -0.946698
+ 2.341e+11Hz -0.234356 -0.94654
+ 2.342e+11Hz -0.23509 -0.946381
+ 2.343e+11Hz -0.235824 -0.946221
+ 2.344e+11Hz -0.236558 -0.946061
+ 2.345e+11Hz -0.237293 -0.9459
+ 2.346e+11Hz -0.238028 -0.945739
+ 2.347e+11Hz -0.238763 -0.945577
+ 2.348e+11Hz -0.239498 -0.945414
+ 2.349e+11Hz -0.240234 -0.94525
+ 2.35e+11Hz -0.240969 -0.945086
+ 2.351e+11Hz -0.241706 -0.944921
+ 2.352e+11Hz -0.242442 -0.944755
+ 2.353e+11Hz -0.243178 -0.944589
+ 2.354e+11Hz -0.243915 -0.944421
+ 2.355e+11Hz -0.244652 -0.944253
+ 2.356e+11Hz -0.245389 -0.944085
+ 2.357e+11Hz -0.246127 -0.943915
+ 2.358e+11Hz -0.246865 -0.943745
+ 2.359e+11Hz -0.247602 -0.943574
+ 2.36e+11Hz -0.248341 -0.943402
+ 2.361e+11Hz -0.249079 -0.94323
+ 2.362e+11Hz -0.249817 -0.943057
+ 2.363e+11Hz -0.250556 -0.942882
+ 2.364e+11Hz -0.251295 -0.942708
+ 2.365e+11Hz -0.252034 -0.942532
+ 2.366e+11Hz -0.252773 -0.942355
+ 2.367e+11Hz -0.253513 -0.942178
+ 2.368e+11Hz -0.254252 -0.942
+ 2.369e+11Hz -0.254992 -0.941821
+ 2.37e+11Hz -0.255732 -0.941641
+ 2.371e+11Hz -0.256472 -0.94146
+ 2.372e+11Hz -0.257212 -0.941279
+ 2.373e+11Hz -0.257952 -0.941096
+ 2.374e+11Hz -0.258693 -0.940913
+ 2.375e+11Hz -0.259433 -0.940729
+ 2.376e+11Hz -0.260174 -0.940544
+ 2.377e+11Hz -0.260915 -0.940359
+ 2.378e+11Hz -0.261656 -0.940172
+ 2.379e+11Hz -0.262397 -0.939984
+ 2.38e+11Hz -0.263138 -0.939796
+ 2.381e+11Hz -0.263879 -0.939607
+ 2.382e+11Hz -0.26462 -0.939417
+ 2.383e+11Hz -0.265362 -0.939225
+ 2.384e+11Hz -0.266103 -0.939034
+ 2.385e+11Hz -0.266845 -0.938841
+ 2.386e+11Hz -0.267586 -0.938647
+ 2.387e+11Hz -0.268328 -0.938452
+ 2.388e+11Hz -0.269069 -0.938257
+ 2.389e+11Hz -0.269811 -0.93806
+ 2.39e+11Hz -0.270553 -0.937863
+ 2.391e+11Hz -0.271294 -0.937665
+ 2.392e+11Hz -0.272036 -0.937465
+ 2.393e+11Hz -0.272778 -0.937265
+ 2.394e+11Hz -0.273519 -0.937064
+ 2.395e+11Hz -0.274261 -0.936862
+ 2.396e+11Hz -0.275003 -0.936659
+ 2.397e+11Hz -0.275744 -0.936456
+ 2.398e+11Hz -0.276486 -0.936251
+ 2.399e+11Hz -0.277227 -0.936045
+ 2.4e+11Hz -0.277969 -0.935839
+ 2.401e+11Hz -0.27871 -0.935631
+ 2.402e+11Hz -0.279451 -0.935423
+ 2.403e+11Hz -0.280193 -0.935213
+ 2.404e+11Hz -0.280934 -0.935003
+ 2.405e+11Hz -0.281675 -0.934792
+ 2.406e+11Hz -0.282416 -0.93458
+ 2.407e+11Hz -0.283157 -0.934367
+ 2.408e+11Hz -0.283898 -0.934153
+ 2.409e+11Hz -0.284638 -0.933938
+ 2.41e+11Hz -0.285379 -0.933722
+ 2.411e+11Hz -0.286119 -0.933505
+ 2.412e+11Hz -0.286859 -0.933287
+ 2.413e+11Hz -0.287599 -0.933069
+ 2.414e+11Hz -0.288339 -0.932849
+ 2.415e+11Hz -0.289079 -0.932629
+ 2.416e+11Hz -0.289819 -0.932407
+ 2.417e+11Hz -0.290558 -0.932185
+ 2.418e+11Hz -0.291297 -0.931962
+ 2.419e+11Hz -0.292036 -0.931737
+ 2.42e+11Hz -0.292775 -0.931512
+ 2.421e+11Hz -0.293514 -0.931286
+ 2.422e+11Hz -0.294252 -0.931059
+ 2.423e+11Hz -0.29499 -0.930832
+ 2.424e+11Hz -0.295728 -0.930603
+ 2.425e+11Hz -0.296466 -0.930373
+ 2.426e+11Hz -0.297203 -0.930143
+ 2.427e+11Hz -0.29794 -0.929911
+ 2.428e+11Hz -0.298677 -0.929679
+ 2.429e+11Hz -0.299414 -0.929446
+ 2.43e+11Hz -0.30015 -0.929212
+ 2.431e+11Hz -0.300887 -0.928977
+ 2.432e+11Hz -0.301622 -0.928741
+ 2.433e+11Hz -0.302358 -0.928504
+ 2.434e+11Hz -0.303093 -0.928267
+ 2.435e+11Hz -0.303828 -0.928028
+ 2.436e+11Hz -0.304563 -0.927789
+ 2.437e+11Hz -0.305297 -0.927549
+ 2.438e+11Hz -0.306031 -0.927308
+ 2.439e+11Hz -0.306765 -0.927066
+ 2.44e+11Hz -0.307498 -0.926823
+ 2.441e+11Hz -0.308231 -0.926579
+ 2.442e+11Hz -0.308964 -0.926335
+ 2.443e+11Hz -0.309697 -0.92609
+ 2.444e+11Hz -0.310429 -0.925844
+ 2.445e+11Hz -0.31116 -0.925597
+ 2.446e+11Hz -0.311892 -0.925349
+ 2.447e+11Hz -0.312623 -0.925101
+ 2.448e+11Hz -0.313353 -0.924851
+ 2.449e+11Hz -0.314083 -0.924601
+ 2.45e+11Hz -0.314813 -0.92435
+ 2.451e+11Hz -0.315543 -0.924099
+ 2.452e+11Hz -0.316272 -0.923846
+ 2.453e+11Hz -0.317001 -0.923593
+ 2.454e+11Hz -0.317729 -0.923339
+ 2.455e+11Hz -0.318457 -0.923084
+ 2.456e+11Hz -0.319185 -0.922828
+ 2.457e+11Hz -0.319912 -0.922572
+ 2.458e+11Hz -0.320639 -0.922315
+ 2.459e+11Hz -0.321365 -0.922057
+ 2.46e+11Hz -0.322091 -0.921798
+ 2.461e+11Hz -0.322817 -0.921539
+ 2.462e+11Hz -0.323542 -0.921279
+ 2.463e+11Hz -0.324267 -0.921018
+ 2.464e+11Hz -0.324991 -0.920756
+ 2.465e+11Hz -0.325715 -0.920494
+ 2.466e+11Hz -0.326439 -0.920231
+ 2.467e+11Hz -0.327162 -0.919968
+ 2.468e+11Hz -0.327884 -0.919703
+ 2.469e+11Hz -0.328607 -0.919438
+ 2.47e+11Hz -0.329329 -0.919172
+ 2.471e+11Hz -0.33005 -0.918906
+ 2.472e+11Hz -0.330771 -0.918639
+ 2.473e+11Hz -0.331492 -0.918371
+ 2.474e+11Hz -0.332212 -0.918103
+ 2.475e+11Hz -0.332932 -0.917833
+ 2.476e+11Hz -0.333651 -0.917564
+ 2.477e+11Hz -0.33437 -0.917293
+ 2.478e+11Hz -0.335089 -0.917022
+ 2.479e+11Hz -0.335807 -0.91675
+ 2.48e+11Hz -0.336524 -0.916478
+ 2.481e+11Hz -0.337242 -0.916205
+ 2.482e+11Hz -0.337958 -0.915931
+ 2.483e+11Hz -0.338675 -0.915657
+ 2.484e+11Hz -0.339391 -0.915382
+ 2.485e+11Hz -0.340106 -0.915107
+ 2.486e+11Hz -0.340821 -0.914831
+ 2.487e+11Hz -0.341536 -0.914554
+ 2.488e+11Hz -0.342251 -0.914277
+ 2.489e+11Hz -0.342964 -0.913999
+ 2.49e+11Hz -0.343678 -0.91372
+ 2.491e+11Hz -0.344391 -0.913441
+ 2.492e+11Hz -0.345104 -0.913162
+ 2.493e+11Hz -0.345816 -0.912881
+ 2.494e+11Hz -0.346528 -0.912601
+ 2.495e+11Hz -0.347239 -0.912319
+ 2.496e+11Hz -0.34795 -0.912037
+ 2.497e+11Hz -0.348661 -0.911755
+ 2.498e+11Hz -0.349371 -0.911472
+ 2.499e+11Hz -0.350081 -0.911188
+ 2.5e+11Hz -0.35079 -0.910904
+ 2.501e+11Hz -0.351499 -0.910619
+ 2.502e+11Hz -0.352208 -0.910334
+ 2.503e+11Hz -0.352916 -0.910048
+ 2.504e+11Hz -0.353624 -0.909762
+ 2.505e+11Hz -0.354332 -0.909475
+ 2.506e+11Hz -0.355039 -0.909187
+ 2.507e+11Hz -0.355745 -0.908899
+ 2.508e+11Hz -0.356452 -0.908611
+ 2.509e+11Hz -0.357158 -0.908322
+ 2.51e+11Hz -0.357863 -0.908032
+ 2.511e+11Hz -0.358568 -0.907742
+ 2.512e+11Hz -0.359273 -0.907452
+ 2.513e+11Hz -0.359978 -0.907161
+ 2.514e+11Hz -0.360682 -0.906869
+ 2.515e+11Hz -0.361386 -0.906577
+ 2.516e+11Hz -0.362089 -0.906284
+ 2.517e+11Hz -0.362792 -0.905991
+ 2.518e+11Hz -0.363495 -0.905697
+ 2.519e+11Hz -0.364197 -0.905403
+ 2.52e+11Hz -0.364899 -0.905108
+ 2.521e+11Hz -0.3656 -0.904813
+ 2.522e+11Hz -0.366302 -0.904517
+ 2.523e+11Hz -0.367003 -0.904221
+ 2.524e+11Hz -0.367703 -0.903924
+ 2.525e+11Hz -0.368404 -0.903627
+ 2.526e+11Hz -0.369103 -0.903329
+ 2.527e+11Hz -0.369803 -0.903031
+ 2.528e+11Hz -0.370502 -0.902732
+ 2.529e+11Hz -0.371201 -0.902433
+ 2.53e+11Hz -0.3719 -0.902133
+ 2.531e+11Hz -0.372598 -0.901833
+ 2.532e+11Hz -0.373296 -0.901532
+ 2.533e+11Hz -0.373994 -0.901231
+ 2.534e+11Hz -0.374691 -0.900929
+ 2.535e+11Hz -0.375388 -0.900627
+ 2.536e+11Hz -0.376085 -0.900324
+ 2.537e+11Hz -0.376781 -0.90002
+ 2.538e+11Hz -0.377477 -0.899717
+ 2.539e+11Hz -0.378173 -0.899412
+ 2.54e+11Hz -0.378868 -0.899107
+ 2.541e+11Hz -0.379564 -0.898802
+ 2.542e+11Hz -0.380258 -0.898496
+ 2.543e+11Hz -0.380953 -0.89819
+ 2.544e+11Hz -0.381647 -0.897883
+ 2.545e+11Hz -0.382341 -0.897575
+ 2.546e+11Hz -0.383035 -0.897267
+ 2.547e+11Hz -0.383728 -0.896959
+ 2.548e+11Hz -0.384421 -0.89665
+ 2.549e+11Hz -0.385114 -0.89634
+ 2.55e+11Hz -0.385806 -0.89603
+ 2.551e+11Hz -0.386498 -0.89572
+ 2.552e+11Hz -0.38719 -0.895409
+ 2.553e+11Hz -0.387882 -0.895097
+ 2.554e+11Hz -0.388573 -0.894785
+ 2.555e+11Hz -0.389264 -0.894472
+ 2.556e+11Hz -0.389955 -0.894159
+ 2.557e+11Hz -0.390645 -0.893845
+ 2.558e+11Hz -0.391335 -0.893531
+ 2.559e+11Hz -0.392025 -0.893216
+ 2.56e+11Hz -0.392715 -0.892901
+ 2.561e+11Hz -0.393404 -0.892585
+ 2.562e+11Hz -0.394093 -0.892269
+ 2.563e+11Hz -0.394782 -0.891952
+ 2.564e+11Hz -0.39547 -0.891634
+ 2.565e+11Hz -0.396158 -0.891316
+ 2.566e+11Hz -0.396846 -0.890997
+ 2.567e+11Hz -0.397533 -0.890678
+ 2.568e+11Hz -0.39822 -0.890359
+ 2.569e+11Hz -0.398907 -0.890038
+ 2.57e+11Hz -0.399594 -0.889717
+ 2.571e+11Hz -0.40028 -0.889396
+ 2.572e+11Hz -0.400966 -0.889074
+ 2.573e+11Hz -0.401652 -0.888751
+ 2.574e+11Hz -0.402337 -0.888428
+ 2.575e+11Hz -0.403022 -0.888105
+ 2.576e+11Hz -0.403707 -0.88778
+ 2.577e+11Hz -0.404391 -0.887456
+ 2.578e+11Hz -0.405075 -0.88713
+ 2.579e+11Hz -0.405759 -0.886804
+ 2.58e+11Hz -0.406442 -0.886478
+ 2.581e+11Hz -0.407125 -0.886151
+ 2.582e+11Hz -0.407808 -0.885823
+ 2.583e+11Hz -0.408491 -0.885495
+ 2.584e+11Hz -0.409173 -0.885166
+ 2.585e+11Hz -0.409855 -0.884837
+ 2.586e+11Hz -0.410536 -0.884507
+ 2.587e+11Hz -0.411217 -0.884176
+ 2.588e+11Hz -0.411898 -0.883845
+ 2.589e+11Hz -0.412578 -0.883513
+ 2.59e+11Hz -0.413258 -0.883181
+ 2.591e+11Hz -0.413938 -0.882848
+ 2.592e+11Hz -0.414617 -0.882515
+ 2.593e+11Hz -0.415296 -0.882181
+ 2.594e+11Hz -0.415975 -0.881846
+ 2.595e+11Hz -0.416653 -0.881511
+ 2.596e+11Hz -0.417331 -0.881175
+ 2.597e+11Hz -0.418009 -0.880839
+ 2.598e+11Hz -0.418686 -0.880502
+ 2.599e+11Hz -0.419363 -0.880164
+ 2.6e+11Hz -0.420039 -0.879826
+ 2.601e+11Hz -0.420715 -0.879487
+ 2.602e+11Hz -0.42139 -0.879148
+ 2.603e+11Hz -0.422066 -0.878808
+ 2.604e+11Hz -0.42274 -0.878468
+ 2.605e+11Hz -0.423415 -0.878127
+ 2.606e+11Hz -0.424089 -0.877785
+ 2.607e+11Hz -0.424762 -0.877443
+ 2.608e+11Hz -0.425435 -0.8771
+ 2.609e+11Hz -0.426108 -0.876757
+ 2.61e+11Hz -0.42678 -0.876413
+ 2.611e+11Hz -0.427452 -0.876069
+ 2.612e+11Hz -0.428124 -0.875724
+ 2.613e+11Hz -0.428794 -0.875378
+ 2.614e+11Hz -0.429465 -0.875032
+ 2.615e+11Hz -0.430135 -0.874686
+ 2.616e+11Hz -0.430805 -0.874338
+ 2.617e+11Hz -0.431474 -0.873991
+ 2.618e+11Hz -0.432143 -0.873642
+ 2.619e+11Hz -0.432811 -0.873293
+ 2.62e+11Hz -0.433479 -0.872944
+ 2.621e+11Hz -0.434146 -0.872594
+ 2.622e+11Hz -0.434813 -0.872244
+ 2.623e+11Hz -0.435479 -0.871893
+ 2.624e+11Hz -0.436145 -0.871541
+ 2.625e+11Hz -0.43681 -0.871189
+ 2.626e+11Hz -0.437475 -0.870837
+ 2.627e+11Hz -0.43814 -0.870484
+ 2.628e+11Hz -0.438803 -0.87013
+ 2.629e+11Hz -0.439467 -0.869776
+ 2.63e+11Hz -0.44013 -0.869422
+ 2.631e+11Hz -0.440792 -0.869067
+ 2.632e+11Hz -0.441454 -0.868711
+ 2.633e+11Hz -0.442115 -0.868355
+ 2.634e+11Hz -0.442776 -0.867999
+ 2.635e+11Hz -0.443437 -0.867642
+ 2.636e+11Hz -0.444096 -0.867284
+ 2.637e+11Hz -0.444756 -0.866926
+ 2.638e+11Hz -0.445415 -0.866568
+ 2.639e+11Hz -0.446073 -0.866209
+ 2.64e+11Hz -0.44673 -0.86585
+ 2.641e+11Hz -0.447388 -0.86549
+ 2.642e+11Hz -0.448044 -0.86513
+ 2.643e+11Hz -0.4487 -0.86477
+ 2.644e+11Hz -0.449356 -0.864409
+ 2.645e+11Hz -0.450011 -0.864048
+ 2.646e+11Hz -0.450666 -0.863686
+ 2.647e+11Hz -0.45132 -0.863324
+ 2.648e+11Hz -0.451973 -0.862961
+ 2.649e+11Hz -0.452626 -0.862598
+ 2.65e+11Hz -0.453278 -0.862235
+ 2.651e+11Hz -0.45393 -0.861871
+ 2.652e+11Hz -0.454581 -0.861507
+ 2.653e+11Hz -0.455232 -0.861143
+ 2.654e+11Hz -0.455882 -0.860778
+ 2.655e+11Hz -0.456532 -0.860413
+ 2.656e+11Hz -0.457181 -0.860048
+ 2.657e+11Hz -0.45783 -0.859682
+ 2.658e+11Hz -0.458478 -0.859316
+ 2.659e+11Hz -0.459125 -0.858949
+ 2.66e+11Hz -0.459772 -0.858583
+ 2.661e+11Hz -0.460419 -0.858216
+ 2.662e+11Hz -0.461065 -0.857848
+ 2.663e+11Hz -0.46171 -0.857481
+ 2.664e+11Hz -0.462355 -0.857113
+ 2.665e+11Hz -0.462999 -0.856745
+ 2.666e+11Hz -0.463643 -0.856377
+ 2.667e+11Hz -0.464286 -0.856008
+ 2.668e+11Hz -0.464929 -0.855639
+ 2.669e+11Hz -0.465571 -0.85527
+ 2.67e+11Hz -0.466213 -0.854901
+ 2.671e+11Hz -0.466854 -0.854531
+ 2.672e+11Hz -0.467495 -0.854161
+ 2.673e+11Hz -0.468135 -0.853791
+ 2.674e+11Hz -0.468775 -0.853421
+ 2.675e+11Hz -0.469414 -0.85305
+ 2.676e+11Hz -0.470053 -0.85268
+ 2.677e+11Hz -0.470691 -0.852309
+ 2.678e+11Hz -0.471329 -0.851938
+ 2.679e+11Hz -0.471966 -0.851567
+ 2.68e+11Hz -0.472603 -0.851196
+ 2.681e+11Hz -0.473239 -0.850824
+ 2.682e+11Hz -0.473875 -0.850452
+ 2.683e+11Hz -0.47451 -0.850081
+ 2.684e+11Hz -0.475145 -0.849709
+ 2.685e+11Hz -0.47578 -0.849337
+ 2.686e+11Hz -0.476414 -0.848964
+ 2.687e+11Hz -0.477048 -0.848592
+ 2.688e+11Hz -0.477681 -0.84822
+ 2.689e+11Hz -0.478314 -0.847847
+ 2.69e+11Hz -0.478946 -0.847475
+ 2.691e+11Hz -0.479578 -0.847102
+ 2.692e+11Hz -0.48021 -0.846729
+ 2.693e+11Hz -0.480841 -0.846356
+ 2.694e+11Hz -0.481472 -0.845983
+ 2.695e+11Hz -0.482102 -0.84561
+ 2.696e+11Hz -0.482732 -0.845237
+ 2.697e+11Hz -0.483362 -0.844864
+ 2.698e+11Hz -0.483992 -0.84449
+ 2.699e+11Hz -0.484621 -0.844117
+ 2.7e+11Hz -0.48525 -0.843743
+ 2.701e+11Hz -0.485878 -0.84337
+ 2.702e+11Hz -0.486506 -0.842996
+ 2.703e+11Hz -0.487134 -0.842623
+ 2.704e+11Hz -0.487761 -0.842249
+ 2.705e+11Hz -0.488389 -0.841875
+ 2.706e+11Hz -0.489016 -0.841502
+ 2.707e+11Hz -0.489642 -0.841128
+ 2.708e+11Hz -0.490269 -0.840754
+ 2.709e+11Hz -0.490895 -0.84038
+ 2.71e+11Hz -0.491521 -0.840006
+ 2.711e+11Hz -0.492147 -0.839633
+ 2.712e+11Hz -0.492772 -0.839259
+ 2.713e+11Hz -0.493398 -0.838885
+ 2.714e+11Hz -0.494023 -0.838511
+ 2.715e+11Hz -0.494648 -0.838137
+ 2.716e+11Hz -0.495272 -0.837763
+ 2.717e+11Hz -0.495897 -0.837388
+ 2.718e+11Hz -0.496522 -0.837014
+ 2.719e+11Hz -0.497146 -0.83664
+ 2.72e+11Hz -0.49777 -0.836266
+ 2.721e+11Hz -0.498394 -0.835892
+ 2.722e+11Hz -0.499018 -0.835517
+ 2.723e+11Hz -0.499642 -0.835143
+ 2.724e+11Hz -0.500265 -0.834769
+ 2.725e+11Hz -0.500889 -0.834394
+ 2.726e+11Hz -0.501513 -0.83402
+ 2.727e+11Hz -0.502136 -0.833646
+ 2.728e+11Hz -0.502759 -0.833271
+ 2.729e+11Hz -0.503383 -0.832897
+ 2.73e+11Hz -0.504006 -0.832522
+ 2.731e+11Hz -0.50463 -0.832147
+ 2.732e+11Hz -0.505253 -0.831772
+ 2.733e+11Hz -0.505876 -0.831398
+ 2.734e+11Hz -0.506499 -0.831023
+ 2.735e+11Hz -0.507123 -0.830648
+ 2.736e+11Hz -0.507746 -0.830273
+ 2.737e+11Hz -0.50837 -0.829898
+ 2.738e+11Hz -0.508993 -0.829522
+ 2.739e+11Hz -0.509616 -0.829147
+ 2.74e+11Hz -0.51024 -0.828772
+ 2.741e+11Hz -0.510864 -0.828396
+ 2.742e+11Hz -0.511487 -0.828021
+ 2.743e+11Hz -0.512111 -0.827645
+ 2.744e+11Hz -0.512735 -0.827269
+ 2.745e+11Hz -0.513359 -0.826893
+ 2.746e+11Hz -0.513983 -0.826517
+ 2.747e+11Hz -0.514607 -0.82614
+ 2.748e+11Hz -0.515232 -0.825764
+ 2.749e+11Hz -0.515856 -0.825387
+ 2.75e+11Hz -0.516481 -0.82501
+ 2.751e+11Hz -0.517106 -0.824633
+ 2.752e+11Hz -0.517731 -0.824256
+ 2.753e+11Hz -0.518356 -0.823879
+ 2.754e+11Hz -0.518981 -0.823501
+ 2.755e+11Hz -0.519607 -0.823123
+ 2.756e+11Hz -0.520232 -0.822745
+ 2.757e+11Hz -0.520858 -0.822367
+ 2.758e+11Hz -0.521484 -0.821988
+ 2.759e+11Hz -0.522111 -0.821609
+ 2.76e+11Hz -0.522737 -0.82123
+ 2.761e+11Hz -0.523364 -0.820851
+ 2.762e+11Hz -0.523991 -0.820471
+ 2.763e+11Hz -0.524618 -0.820091
+ 2.764e+11Hz -0.525246 -0.819711
+ 2.765e+11Hz -0.525873 -0.81933
+ 2.766e+11Hz -0.526501 -0.818949
+ 2.767e+11Hz -0.527129 -0.818568
+ 2.768e+11Hz -0.527758 -0.818186
+ 2.769e+11Hz -0.528386 -0.817804
+ 2.77e+11Hz -0.529015 -0.817422
+ 2.771e+11Hz -0.529645 -0.817039
+ 2.772e+11Hz -0.530274 -0.816655
+ 2.773e+11Hz -0.530904 -0.816272
+ 2.774e+11Hz -0.531534 -0.815888
+ 2.775e+11Hz -0.532164 -0.815503
+ 2.776e+11Hz -0.532795 -0.815118
+ 2.777e+11Hz -0.533426 -0.814733
+ 2.778e+11Hz -0.534057 -0.814347
+ 2.779e+11Hz -0.534688 -0.81396
+ 2.78e+11Hz -0.53532 -0.813573
+ 2.781e+11Hz -0.535952 -0.813186
+ 2.782e+11Hz -0.536584 -0.812798
+ 2.783e+11Hz -0.537217 -0.812409
+ 2.784e+11Hz -0.537849 -0.81202
+ 2.785e+11Hz -0.538482 -0.81163
+ 2.786e+11Hz -0.539116 -0.81124
+ 2.787e+11Hz -0.539749 -0.810849
+ 2.788e+11Hz -0.540383 -0.810457
+ 2.789e+11Hz -0.541017 -0.810065
+ 2.79e+11Hz -0.541652 -0.809673
+ 2.791e+11Hz -0.542287 -0.809279
+ 2.792e+11Hz -0.542921 -0.808885
+ 2.793e+11Hz -0.543557 -0.80849
+ 2.794e+11Hz -0.544192 -0.808095
+ 2.795e+11Hz -0.544828 -0.807699
+ 2.796e+11Hz -0.545464 -0.807302
+ 2.797e+11Hz -0.5461 -0.806904
+ 2.798e+11Hz -0.546736 -0.806506
+ 2.799e+11Hz -0.547373 -0.806107
+ 2.8e+11Hz -0.54801 -0.805707
+ 2.801e+11Hz -0.548647 -0.805307
+ 2.802e+11Hz -0.549284 -0.804905
+ 2.803e+11Hz -0.549921 -0.804503
+ 2.804e+11Hz -0.550559 -0.8041
+ 2.805e+11Hz -0.551197 -0.803697
+ 2.806e+11Hz -0.551835 -0.803292
+ 2.807e+11Hz -0.552473 -0.802887
+ 2.808e+11Hz -0.553111 -0.80248
+ 2.809e+11Hz -0.55375 -0.802073
+ 2.81e+11Hz -0.554389 -0.801665
+ 2.811e+11Hz -0.555027 -0.801256
+ 2.812e+11Hz -0.555666 -0.800847
+ 2.813e+11Hz -0.556305 -0.800436
+ 2.814e+11Hz -0.556945 -0.800024
+ 2.815e+11Hz -0.557584 -0.799612
+ 2.816e+11Hz -0.558223 -0.799198
+ 2.817e+11Hz -0.558863 -0.798784
+ 2.818e+11Hz -0.559502 -0.798369
+ 2.819e+11Hz -0.560142 -0.797953
+ 2.82e+11Hz -0.560781 -0.797535
+ 2.821e+11Hz -0.561421 -0.797117
+ 2.822e+11Hz -0.562061 -0.796698
+ 2.823e+11Hz -0.5627 -0.796278
+ 2.824e+11Hz -0.56334 -0.795857
+ 2.825e+11Hz -0.56398 -0.795435
+ 2.826e+11Hz -0.564619 -0.795012
+ 2.827e+11Hz -0.565259 -0.794588
+ 2.828e+11Hz -0.565899 -0.794162
+ 2.829e+11Hz -0.566538 -0.793736
+ 2.83e+11Hz -0.567178 -0.793309
+ 2.831e+11Hz -0.567817 -0.792881
+ 2.832e+11Hz -0.568456 -0.792452
+ 2.833e+11Hz -0.569096 -0.792021
+ 2.834e+11Hz -0.569735 -0.79159
+ 2.835e+11Hz -0.570374 -0.791158
+ 2.836e+11Hz -0.571012 -0.790724
+ 2.837e+11Hz -0.571651 -0.79029
+ 2.838e+11Hz -0.572289 -0.789854
+ 2.839e+11Hz -0.572928 -0.789418
+ 2.84e+11Hz -0.573566 -0.78898
+ 2.841e+11Hz -0.574204 -0.788541
+ 2.842e+11Hz -0.574841 -0.788102
+ 2.843e+11Hz -0.575479 -0.787661
+ 2.844e+11Hz -0.576116 -0.787219
+ 2.845e+11Hz -0.576753 -0.786776
+ 2.846e+11Hz -0.577389 -0.786332
+ 2.847e+11Hz -0.578026 -0.785887
+ 2.848e+11Hz -0.578662 -0.78544
+ 2.849e+11Hz -0.579297 -0.784993
+ 2.85e+11Hz -0.579933 -0.784545
+ 2.851e+11Hz -0.580568 -0.784095
+ 2.852e+11Hz -0.581202 -0.783645
+ 2.853e+11Hz -0.581836 -0.783193
+ 2.854e+11Hz -0.58247 -0.782741
+ 2.855e+11Hz -0.583104 -0.782287
+ 2.856e+11Hz -0.583737 -0.781833
+ 2.857e+11Hz -0.58437 -0.781377
+ 2.858e+11Hz -0.585002 -0.78092
+ 2.859e+11Hz -0.585633 -0.780462
+ 2.86e+11Hz -0.586265 -0.780003
+ 2.861e+11Hz -0.586896 -0.779544
+ 2.862e+11Hz -0.587526 -0.779083
+ 2.863e+11Hz -0.588156 -0.778621
+ 2.864e+11Hz -0.588785 -0.778158
+ 2.865e+11Hz -0.589414 -0.777694
+ 2.866e+11Hz -0.590042 -0.777229
+ 2.867e+11Hz -0.59067 -0.776763
+ 2.868e+11Hz -0.591297 -0.776296
+ 2.869e+11Hz -0.591923 -0.775828
+ 2.87e+11Hz -0.592549 -0.775359
+ 2.871e+11Hz -0.593175 -0.774889
+ 2.872e+11Hz -0.593799 -0.774418
+ 2.873e+11Hz -0.594423 -0.773946
+ 2.874e+11Hz -0.595047 -0.773473
+ 2.875e+11Hz -0.59567 -0.773
+ 2.876e+11Hz -0.596292 -0.772525
+ 2.877e+11Hz -0.596914 -0.772049
+ 2.878e+11Hz -0.597535 -0.771573
+ 2.879e+11Hz -0.598155 -0.771095
+ 2.88e+11Hz -0.598774 -0.770617
+ 2.881e+11Hz -0.599393 -0.770138
+ 2.882e+11Hz -0.600011 -0.769658
+ 2.883e+11Hz -0.600629 -0.769177
+ 2.884e+11Hz -0.601246 -0.768695
+ 2.885e+11Hz -0.601862 -0.768212
+ 2.886e+11Hz -0.602477 -0.767729
+ 2.887e+11Hz -0.603091 -0.767245
+ 2.888e+11Hz -0.603705 -0.766759
+ 2.889e+11Hz -0.604318 -0.766273
+ 2.89e+11Hz -0.604931 -0.765787
+ 2.891e+11Hz -0.605542 -0.765299
+ 2.892e+11Hz -0.606153 -0.764811
+ 2.893e+11Hz -0.606763 -0.764322
+ 2.894e+11Hz -0.607372 -0.763832
+ 2.895e+11Hz -0.607981 -0.763341
+ 2.896e+11Hz -0.608588 -0.76285
+ 2.897e+11Hz -0.609195 -0.762358
+ 2.898e+11Hz -0.609801 -0.761865
+ 2.899e+11Hz -0.610407 -0.761372
+ 2.9e+11Hz -0.611011 -0.760878
+ 2.901e+11Hz -0.611615 -0.760383
+ 2.902e+11Hz -0.612218 -0.759888
+ 2.903e+11Hz -0.61282 -0.759392
+ 2.904e+11Hz -0.613421 -0.758895
+ 2.905e+11Hz -0.614021 -0.758398
+ 2.906e+11Hz -0.614621 -0.7579
+ 2.907e+11Hz -0.61522 -0.757401
+ 2.908e+11Hz -0.615818 -0.756902
+ 2.909e+11Hz -0.616415 -0.756402
+ 2.91e+11Hz -0.617011 -0.755902
+ 2.911e+11Hz -0.617607 -0.755401
+ 2.912e+11Hz -0.618202 -0.7549
+ 2.913e+11Hz -0.618796 -0.754398
+ 2.914e+11Hz -0.619389 -0.753896
+ 2.915e+11Hz -0.619981 -0.753393
+ 2.916e+11Hz -0.620573 -0.752889
+ 2.917e+11Hz -0.621163 -0.752385
+ 2.918e+11Hz -0.621753 -0.751881
+ 2.919e+11Hz -0.622342 -0.751376
+ 2.92e+11Hz -0.622931 -0.750871
+ 2.921e+11Hz -0.623518 -0.750365
+ 2.922e+11Hz -0.624105 -0.749859
+ 2.923e+11Hz -0.624691 -0.749352
+ 2.924e+11Hz -0.625276 -0.748845
+ 2.925e+11Hz -0.625861 -0.748338
+ 2.926e+11Hz -0.626444 -0.74783
+ 2.927e+11Hz -0.627027 -0.747322
+ 2.928e+11Hz -0.627609 -0.746813
+ 2.929e+11Hz -0.628191 -0.746304
+ 2.93e+11Hz -0.628771 -0.745795
+ 2.931e+11Hz -0.629351 -0.745285
+ 2.932e+11Hz -0.62993 -0.744775
+ 2.933e+11Hz -0.630509 -0.744264
+ 2.934e+11Hz -0.631086 -0.743754
+ 2.935e+11Hz -0.631663 -0.743243
+ 2.936e+11Hz -0.63224 -0.742731
+ 2.937e+11Hz -0.632815 -0.74222
+ 2.938e+11Hz -0.63339 -0.741708
+ 2.939e+11Hz -0.633964 -0.741195
+ 2.94e+11Hz -0.634538 -0.740683
+ 2.941e+11Hz -0.63511 -0.74017
+ 2.942e+11Hz -0.635683 -0.739657
+ 2.943e+11Hz -0.636254 -0.739143
+ 2.944e+11Hz -0.636825 -0.73863
+ 2.945e+11Hz -0.637395 -0.738116
+ 2.946e+11Hz -0.637965 -0.737602
+ 2.947e+11Hz -0.638533 -0.737087
+ 2.948e+11Hz -0.639102 -0.736573
+ 2.949e+11Hz -0.639669 -0.736058
+ 2.95e+11Hz -0.640237 -0.735543
+ 2.951e+11Hz -0.640803 -0.735027
+ 2.952e+11Hz -0.641369 -0.734512
+ 2.953e+11Hz -0.641934 -0.733996
+ 2.954e+11Hz -0.642499 -0.73348
+ 2.955e+11Hz -0.643063 -0.732963
+ 2.956e+11Hz -0.643627 -0.732447
+ 2.957e+11Hz -0.64419 -0.73193
+ 2.958e+11Hz -0.644752 -0.731413
+ 2.959e+11Hz -0.645314 -0.730896
+ 2.96e+11Hz -0.645876 -0.730378
+ 2.961e+11Hz -0.646437 -0.729861
+ 2.962e+11Hz -0.646997 -0.729343
+ 2.963e+11Hz -0.647557 -0.728825
+ 2.964e+11Hz -0.648117 -0.728307
+ 2.965e+11Hz -0.648676 -0.727788
+ 2.966e+11Hz -0.649235 -0.727269
+ 2.967e+11Hz -0.649793 -0.72675
+ 2.968e+11Hz -0.65035 -0.726231
+ 2.969e+11Hz -0.650908 -0.725712
+ 2.97e+11Hz -0.651464 -0.725192
+ 2.971e+11Hz -0.652021 -0.724672
+ 2.972e+11Hz -0.652577 -0.724152
+ 2.973e+11Hz -0.653132 -0.723631
+ 2.974e+11Hz -0.653687 -0.723111
+ 2.975e+11Hz -0.654242 -0.72259
+ 2.976e+11Hz -0.654797 -0.722069
+ 2.977e+11Hz -0.655351 -0.721547
+ 2.978e+11Hz -0.655904 -0.721026
+ 2.979e+11Hz -0.656457 -0.720504
+ 2.98e+11Hz -0.65701 -0.719981
+ 2.981e+11Hz -0.657563 -0.719459
+ 2.982e+11Hz -0.658115 -0.718936
+ 2.983e+11Hz -0.658667 -0.718413
+ 2.984e+11Hz -0.659218 -0.71789
+ 2.985e+11Hz -0.659769 -0.717366
+ 2.986e+11Hz -0.66032 -0.716842
+ 2.987e+11Hz -0.66087 -0.716318
+ 2.988e+11Hz -0.66142 -0.715793
+ 2.989e+11Hz -0.66197 -0.715268
+ 2.99e+11Hz -0.66252 -0.714743
+ 2.991e+11Hz -0.663069 -0.714218
+ 2.992e+11Hz -0.663618 -0.713692
+ 2.993e+11Hz -0.664166 -0.713165
+ 2.994e+11Hz -0.664715 -0.712639
+ 2.995e+11Hz -0.665262 -0.712112
+ 2.996e+11Hz -0.66581 -0.711584
+ 2.997e+11Hz -0.666357 -0.711057
+ 2.998e+11Hz -0.666905 -0.710528
+ 2.999e+11Hz -0.667451 -0.71
+ 3e+11Hz -0.667998 -0.709471
+ ]

A21 %vd(10 3) %vd(21, 22) xfer3
.model xfer3 xfer R_I=true table=[
+ 0Hz 0.995382 0
+ 1e+08Hz 0.995382 -0.000812217
+ 2e+08Hz 0.99538 -0.00162442
+ 3e+08Hz 0.995377 -0.0024366
+ 4e+08Hz 0.995372 -0.00324873
+ 5e+08Hz 0.995367 -0.00406082
+ 6e+08Hz 0.99536 -0.00487284
+ 7e+08Hz 0.995352 -0.00568478
+ 8e+08Hz 0.995343 -0.00649662
+ 9e+08Hz 0.995333 -0.00730836
+ 1e+09Hz 0.995321 -0.00811999
+ 1.1e+09Hz 0.995308 -0.00893148
+ 1.2e+09Hz 0.995294 -0.00974282
+ 1.3e+09Hz 0.995279 -0.010554
+ 1.4e+09Hz 0.995263 -0.011365
+ 1.5e+09Hz 0.995245 -0.0121759
+ 1.6e+09Hz 0.995226 -0.0129865
+ 1.7e+09Hz 0.995206 -0.013797
+ 1.8e+09Hz 0.995185 -0.0146072
+ 1.9e+09Hz 0.995163 -0.0154172
+ 2e+09Hz 0.995139 -0.0162269
+ 2.1e+09Hz 0.995115 -0.0170364
+ 2.2e+09Hz 0.995089 -0.0178456
+ 2.3e+09Hz 0.995062 -0.0186546
+ 2.4e+09Hz 0.995034 -0.0194632
+ 2.5e+09Hz 0.995005 -0.0202716
+ 2.6e+09Hz 0.994974 -0.0210796
+ 2.7e+09Hz 0.994943 -0.0218873
+ 2.8e+09Hz 0.99491 -0.0226947
+ 2.9e+09Hz 0.994876 -0.0235018
+ 3e+09Hz 0.994841 -0.0243085
+ 3.1e+09Hz 0.994806 -0.0251148
+ 3.2e+09Hz 0.994768 -0.0259208
+ 3.3e+09Hz 0.99473 -0.0267263
+ 3.4e+09Hz 0.994691 -0.0275315
+ 3.5e+09Hz 0.994651 -0.0283363
+ 3.6e+09Hz 0.99461 -0.0291407
+ 3.7e+09Hz 0.994567 -0.0299446
+ 3.8e+09Hz 0.994524 -0.0307482
+ 3.9e+09Hz 0.99448 -0.0315512
+ 4e+09Hz 0.994434 -0.0323539
+ 4.1e+09Hz 0.994388 -0.0331561
+ 4.2e+09Hz 0.99434 -0.0339578
+ 4.3e+09Hz 0.994292 -0.0347591
+ 4.4e+09Hz 0.994243 -0.0355599
+ 4.5e+09Hz 0.994192 -0.0363602
+ 4.6e+09Hz 0.994141 -0.0371601
+ 4.7e+09Hz 0.994089 -0.0379594
+ 4.8e+09Hz 0.994036 -0.0387583
+ 4.9e+09Hz 0.993982 -0.0395566
+ 5e+09Hz 0.993927 -0.0403545
+ 5.1e+09Hz 0.993871 -0.0411518
+ 5.2e+09Hz 0.993814 -0.0419486
+ 5.3e+09Hz 0.993757 -0.0427449
+ 5.4e+09Hz 0.993698 -0.0435407
+ 5.5e+09Hz 0.993639 -0.0443359
+ 5.6e+09Hz 0.993579 -0.0451306
+ 5.7e+09Hz 0.993518 -0.0459248
+ 5.8e+09Hz 0.993456 -0.0467184
+ 5.9e+09Hz 0.993394 -0.0475115
+ 6e+09Hz 0.99333 -0.048304
+ 6.1e+09Hz 0.993266 -0.049096
+ 6.2e+09Hz 0.993201 -0.0498875
+ 6.3e+09Hz 0.993135 -0.0506783
+ 6.4e+09Hz 0.993069 -0.0514687
+ 6.5e+09Hz 0.993002 -0.0522585
+ 6.6e+09Hz 0.992934 -0.0530477
+ 6.7e+09Hz 0.992865 -0.0538364
+ 6.8e+09Hz 0.992796 -0.0546245
+ 6.9e+09Hz 0.992726 -0.0554121
+ 7e+09Hz 0.992655 -0.0561991
+ 7.1e+09Hz 0.992584 -0.0569855
+ 7.2e+09Hz 0.992512 -0.0577714
+ 7.3e+09Hz 0.992439 -0.0585568
+ 7.4e+09Hz 0.992366 -0.0593416
+ 7.5e+09Hz 0.992292 -0.0601258
+ 7.6e+09Hz 0.992217 -0.0609095
+ 7.7e+09Hz 0.992142 -0.0616927
+ 7.8e+09Hz 0.992066 -0.0624753
+ 7.9e+09Hz 0.99199 -0.0632574
+ 8e+09Hz 0.991913 -0.0640389
+ 8.1e+09Hz 0.991836 -0.0648199
+ 8.2e+09Hz 0.991758 -0.0656004
+ 8.3e+09Hz 0.991679 -0.0663804
+ 8.4e+09Hz 0.9916 -0.0671598
+ 8.5e+09Hz 0.991521 -0.0679387
+ 8.6e+09Hz 0.99144 -0.0687171
+ 8.7e+09Hz 0.99136 -0.0694949
+ 8.8e+09Hz 0.991279 -0.0702723
+ 8.9e+09Hz 0.991197 -0.0710492
+ 9e+09Hz 0.991115 -0.0718255
+ 9.1e+09Hz 0.991033 -0.0726014
+ 9.2e+09Hz 0.99095 -0.0733768
+ 9.3e+09Hz 0.990866 -0.0741517
+ 9.4e+09Hz 0.990782 -0.0749261
+ 9.5e+09Hz 0.990698 -0.0757001
+ 9.6e+09Hz 0.990613 -0.0764736
+ 9.7e+09Hz 0.990528 -0.0772466
+ 9.8e+09Hz 0.990443 -0.0780192
+ 9.9e+09Hz 0.990357 -0.0787913
+ 1e+10Hz 0.99027 -0.079563
+ 1.01e+10Hz 0.990184 -0.0803343
+ 1.02e+10Hz 0.990097 -0.0811051
+ 1.03e+10Hz 0.990009 -0.0818755
+ 1.04e+10Hz 0.989921 -0.0826455
+ 1.05e+10Hz 0.989833 -0.0834151
+ 1.06e+10Hz 0.989744 -0.0841844
+ 1.07e+10Hz 0.989655 -0.0849532
+ 1.08e+10Hz 0.989566 -0.0857216
+ 1.09e+10Hz 0.989477 -0.0864897
+ 1.1e+10Hz 0.989387 -0.0872574
+ 1.11e+10Hz 0.989296 -0.0880247
+ 1.12e+10Hz 0.989206 -0.0887917
+ 1.13e+10Hz 0.989115 -0.0895584
+ 1.14e+10Hz 0.989023 -0.0903247
+ 1.15e+10Hz 0.988932 -0.0910906
+ 1.16e+10Hz 0.98884 -0.0918563
+ 1.17e+10Hz 0.988748 -0.0926217
+ 1.18e+10Hz 0.988655 -0.0933867
+ 1.19e+10Hz 0.988563 -0.0941515
+ 1.2e+10Hz 0.988469 -0.0949159
+ 1.21e+10Hz 0.988376 -0.0956801
+ 1.22e+10Hz 0.988282 -0.096444
+ 1.23e+10Hz 0.988188 -0.0972077
+ 1.24e+10Hz 0.988094 -0.0979711
+ 1.25e+10Hz 0.988 -0.0987343
+ 1.26e+10Hz 0.987905 -0.0994972
+ 1.27e+10Hz 0.98781 -0.10026
+ 1.28e+10Hz 0.987714 -0.101022
+ 1.29e+10Hz 0.987618 -0.101785
+ 1.3e+10Hz 0.987523 -0.102547
+ 1.31e+10Hz 0.987426 -0.103309
+ 1.32e+10Hz 0.98733 -0.10407
+ 1.33e+10Hz 0.987233 -0.104832
+ 1.34e+10Hz 0.987136 -0.105593
+ 1.35e+10Hz 0.987038 -0.106354
+ 1.36e+10Hz 0.986941 -0.107115
+ 1.37e+10Hz 0.986843 -0.107876
+ 1.38e+10Hz 0.986744 -0.108637
+ 1.39e+10Hz 0.986646 -0.109397
+ 1.4e+10Hz 0.986547 -0.110158
+ 1.41e+10Hz 0.986448 -0.110918
+ 1.42e+10Hz 0.986348 -0.111678
+ 1.43e+10Hz 0.986249 -0.112438
+ 1.44e+10Hz 0.986149 -0.113198
+ 1.45e+10Hz 0.986048 -0.113958
+ 1.46e+10Hz 0.985948 -0.114718
+ 1.47e+10Hz 0.985847 -0.115478
+ 1.48e+10Hz 0.985745 -0.116237
+ 1.49e+10Hz 0.985644 -0.116997
+ 1.5e+10Hz 0.985542 -0.117756
+ 1.51e+10Hz 0.98544 -0.118516
+ 1.52e+10Hz 0.985337 -0.119275
+ 1.53e+10Hz 0.985234 -0.120035
+ 1.54e+10Hz 0.985131 -0.120794
+ 1.55e+10Hz 0.985028 -0.121554
+ 1.56e+10Hz 0.984924 -0.122313
+ 1.57e+10Hz 0.98482 -0.123072
+ 1.58e+10Hz 0.984715 -0.123831
+ 1.59e+10Hz 0.98461 -0.124591
+ 1.6e+10Hz 0.984505 -0.12535
+ 1.61e+10Hz 0.984399 -0.126109
+ 1.62e+10Hz 0.984293 -0.126869
+ 1.63e+10Hz 0.984187 -0.127628
+ 1.64e+10Hz 0.98408 -0.128387
+ 1.65e+10Hz 0.983973 -0.129147
+ 1.66e+10Hz 0.983865 -0.129906
+ 1.67e+10Hz 0.983758 -0.130665
+ 1.68e+10Hz 0.983649 -0.131425
+ 1.69e+10Hz 0.983541 -0.132184
+ 1.7e+10Hz 0.983431 -0.132944
+ 1.71e+10Hz 0.983322 -0.133703
+ 1.72e+10Hz 0.983212 -0.134463
+ 1.73e+10Hz 0.983102 -0.135222
+ 1.74e+10Hz 0.982991 -0.135982
+ 1.75e+10Hz 0.98288 -0.136742
+ 1.76e+10Hz 0.982768 -0.137502
+ 1.77e+10Hz 0.982656 -0.138262
+ 1.78e+10Hz 0.982543 -0.139021
+ 1.79e+10Hz 0.98243 -0.139781
+ 1.8e+10Hz 0.982317 -0.140541
+ 1.81e+10Hz 0.982203 -0.141302
+ 1.82e+10Hz 0.982088 -0.142062
+ 1.83e+10Hz 0.981973 -0.142822
+ 1.84e+10Hz 0.981858 -0.143582
+ 1.85e+10Hz 0.981742 -0.144343
+ 1.86e+10Hz 0.981625 -0.145103
+ 1.87e+10Hz 0.981508 -0.145863
+ 1.88e+10Hz 0.981391 -0.146624
+ 1.89e+10Hz 0.981273 -0.147385
+ 1.9e+10Hz 0.981154 -0.148145
+ 1.91e+10Hz 0.981035 -0.148906
+ 1.92e+10Hz 0.980916 -0.149667
+ 1.93e+10Hz 0.980796 -0.150428
+ 1.94e+10Hz 0.980675 -0.151189
+ 1.95e+10Hz 0.980554 -0.15195
+ 1.96e+10Hz 0.980432 -0.152711
+ 1.97e+10Hz 0.980309 -0.153472
+ 1.98e+10Hz 0.980186 -0.154233
+ 1.99e+10Hz 0.980063 -0.154995
+ 2e+10Hz 0.979939 -0.155756
+ 2.01e+10Hz 0.979814 -0.156517
+ 2.02e+10Hz 0.979689 -0.157279
+ 2.03e+10Hz 0.979563 -0.15804
+ 2.04e+10Hz 0.979436 -0.158802
+ 2.05e+10Hz 0.979309 -0.159563
+ 2.06e+10Hz 0.979182 -0.160325
+ 2.07e+10Hz 0.979053 -0.161087
+ 2.08e+10Hz 0.978924 -0.161848
+ 2.09e+10Hz 0.978795 -0.16261
+ 2.1e+10Hz 0.978665 -0.163372
+ 2.11e+10Hz 0.978534 -0.164134
+ 2.12e+10Hz 0.978402 -0.164896
+ 2.13e+10Hz 0.97827 -0.165657
+ 2.14e+10Hz 0.978137 -0.166419
+ 2.15e+10Hz 0.978004 -0.167181
+ 2.16e+10Hz 0.97787 -0.167943
+ 2.17e+10Hz 0.977735 -0.168705
+ 2.18e+10Hz 0.977599 -0.169467
+ 2.19e+10Hz 0.977463 -0.170229
+ 2.2e+10Hz 0.977327 -0.170991
+ 2.21e+10Hz 0.977189 -0.171753
+ 2.22e+10Hz 0.977051 -0.172515
+ 2.23e+10Hz 0.976912 -0.173276
+ 2.24e+10Hz 0.976773 -0.174038
+ 2.25e+10Hz 0.976633 -0.1748
+ 2.26e+10Hz 0.976492 -0.175562
+ 2.27e+10Hz 0.97635 -0.176324
+ 2.28e+10Hz 0.976208 -0.177085
+ 2.29e+10Hz 0.976065 -0.177847
+ 2.3e+10Hz 0.975921 -0.178609
+ 2.31e+10Hz 0.975777 -0.17937
+ 2.32e+10Hz 0.975632 -0.180132
+ 2.33e+10Hz 0.975486 -0.180893
+ 2.34e+10Hz 0.97534 -0.181655
+ 2.35e+10Hz 0.975192 -0.182416
+ 2.36e+10Hz 0.975045 -0.183177
+ 2.37e+10Hz 0.974896 -0.183938
+ 2.38e+10Hz 0.974747 -0.184699
+ 2.39e+10Hz 0.974597 -0.18546
+ 2.4e+10Hz 0.974446 -0.186221
+ 2.41e+10Hz 0.974294 -0.186982
+ 2.42e+10Hz 0.974142 -0.187743
+ 2.43e+10Hz 0.973989 -0.188503
+ 2.44e+10Hz 0.973836 -0.189263
+ 2.45e+10Hz 0.973682 -0.190024
+ 2.46e+10Hz 0.973527 -0.190784
+ 2.47e+10Hz 0.973371 -0.191544
+ 2.48e+10Hz 0.973214 -0.192304
+ 2.49e+10Hz 0.973057 -0.193064
+ 2.5e+10Hz 0.9729 -0.193823
+ 2.51e+10Hz 0.972741 -0.194583
+ 2.52e+10Hz 0.972582 -0.195342
+ 2.53e+10Hz 0.972422 -0.196101
+ 2.54e+10Hz 0.972261 -0.19686
+ 2.55e+10Hz 0.9721 -0.197619
+ 2.56e+10Hz 0.971938 -0.198378
+ 2.57e+10Hz 0.971775 -0.199136
+ 2.58e+10Hz 0.971611 -0.199894
+ 2.59e+10Hz 0.971447 -0.200652
+ 2.6e+10Hz 0.971282 -0.20141
+ 2.61e+10Hz 0.971117 -0.202168
+ 2.62e+10Hz 0.970951 -0.202925
+ 2.63e+10Hz 0.970784 -0.203683
+ 2.64e+10Hz 0.970616 -0.20444
+ 2.65e+10Hz 0.970448 -0.205197
+ 2.66e+10Hz 0.970279 -0.205953
+ 2.67e+10Hz 0.970109 -0.20671
+ 2.68e+10Hz 0.969939 -0.207466
+ 2.69e+10Hz 0.969768 -0.208222
+ 2.7e+10Hz 0.969596 -0.208978
+ 2.71e+10Hz 0.969424 -0.209733
+ 2.72e+10Hz 0.969251 -0.210489
+ 2.73e+10Hz 0.969077 -0.211244
+ 2.74e+10Hz 0.968903 -0.211998
+ 2.75e+10Hz 0.968728 -0.212753
+ 2.76e+10Hz 0.968552 -0.213507
+ 2.77e+10Hz 0.968376 -0.214261
+ 2.78e+10Hz 0.968199 -0.215015
+ 2.79e+10Hz 0.968021 -0.215769
+ 2.8e+10Hz 0.967843 -0.216522
+ 2.81e+10Hz 0.967664 -0.217275
+ 2.82e+10Hz 0.967485 -0.218028
+ 2.83e+10Hz 0.967304 -0.21878
+ 2.84e+10Hz 0.967124 -0.219533
+ 2.85e+10Hz 0.966942 -0.220285
+ 2.86e+10Hz 0.96676 -0.221036
+ 2.87e+10Hz 0.966578 -0.221788
+ 2.88e+10Hz 0.966395 -0.222539
+ 2.89e+10Hz 0.966211 -0.22329
+ 2.9e+10Hz 0.966026 -0.22404
+ 2.91e+10Hz 0.965842 -0.224791
+ 2.92e+10Hz 0.965656 -0.225541
+ 2.93e+10Hz 0.96547 -0.226291
+ 2.94e+10Hz 0.965283 -0.22704
+ 2.95e+10Hz 0.965096 -0.227789
+ 2.96e+10Hz 0.964908 -0.228538
+ 2.97e+10Hz 0.964719 -0.229287
+ 2.98e+10Hz 0.96453 -0.230035
+ 2.99e+10Hz 0.964341 -0.230784
+ 3e+10Hz 0.96415 -0.231531
+ 3.01e+10Hz 0.96396 -0.232279
+ 3.02e+10Hz 0.963768 -0.233026
+ 3.03e+10Hz 0.963577 -0.233773
+ 3.04e+10Hz 0.963384 -0.23452
+ 3.05e+10Hz 0.963191 -0.235266
+ 3.06e+10Hz 0.962998 -0.236013
+ 3.07e+10Hz 0.962804 -0.236758
+ 3.08e+10Hz 0.962609 -0.237504
+ 3.09e+10Hz 0.962414 -0.238249
+ 3.1e+10Hz 0.962219 -0.238994
+ 3.11e+10Hz 0.962023 -0.239739
+ 3.12e+10Hz 0.961826 -0.240484
+ 3.13e+10Hz 0.961629 -0.241228
+ 3.14e+10Hz 0.961431 -0.241972
+ 3.15e+10Hz 0.961233 -0.242716
+ 3.16e+10Hz 0.961034 -0.243459
+ 3.17e+10Hz 0.960835 -0.244202
+ 3.18e+10Hz 0.960636 -0.244945
+ 3.19e+10Hz 0.960435 -0.245688
+ 3.2e+10Hz 0.960235 -0.24643
+ 3.21e+10Hz 0.960034 -0.247172
+ 3.22e+10Hz 0.959832 -0.247914
+ 3.23e+10Hz 0.95963 -0.248656
+ 3.24e+10Hz 0.959427 -0.249397
+ 3.25e+10Hz 0.959224 -0.250138
+ 3.26e+10Hz 0.959021 -0.250879
+ 3.27e+10Hz 0.958817 -0.25162
+ 3.28e+10Hz 0.958612 -0.25236
+ 3.29e+10Hz 0.958407 -0.2531
+ 3.3e+10Hz 0.958202 -0.25384
+ 3.31e+10Hz 0.957996 -0.25458
+ 3.32e+10Hz 0.957789 -0.255319
+ 3.33e+10Hz 0.957583 -0.256058
+ 3.34e+10Hz 0.957375 -0.256797
+ 3.35e+10Hz 0.957168 -0.257536
+ 3.36e+10Hz 0.956959 -0.258275
+ 3.37e+10Hz 0.956751 -0.259013
+ 3.38e+10Hz 0.956542 -0.259751
+ 3.39e+10Hz 0.956332 -0.260489
+ 3.4e+10Hz 0.956122 -0.261227
+ 3.41e+10Hz 0.955911 -0.261964
+ 3.42e+10Hz 0.955701 -0.262701
+ 3.43e+10Hz 0.955489 -0.263438
+ 3.44e+10Hz 0.955277 -0.264175
+ 3.45e+10Hz 0.955065 -0.264912
+ 3.46e+10Hz 0.954852 -0.265649
+ 3.47e+10Hz 0.954639 -0.266385
+ 3.48e+10Hz 0.954426 -0.267121
+ 3.49e+10Hz 0.954212 -0.267857
+ 3.5e+10Hz 0.953997 -0.268593
+ 3.51e+10Hz 0.953782 -0.269328
+ 3.52e+10Hz 0.953567 -0.270064
+ 3.53e+10Hz 0.953351 -0.270799
+ 3.54e+10Hz 0.953134 -0.271534
+ 3.55e+10Hz 0.952918 -0.272269
+ 3.56e+10Hz 0.952701 -0.273003
+ 3.57e+10Hz 0.952483 -0.273738
+ 3.58e+10Hz 0.952265 -0.274472
+ 3.59e+10Hz 0.952046 -0.275207
+ 3.6e+10Hz 0.951827 -0.275941
+ 3.61e+10Hz 0.951608 -0.276675
+ 3.62e+10Hz 0.951388 -0.277409
+ 3.63e+10Hz 0.951168 -0.278142
+ 3.64e+10Hz 0.950947 -0.278876
+ 3.65e+10Hz 0.950725 -0.279609
+ 3.66e+10Hz 0.950504 -0.280342
+ 3.67e+10Hz 0.950282 -0.281075
+ 3.68e+10Hz 0.950059 -0.281808
+ 3.69e+10Hz 0.949836 -0.282541
+ 3.7e+10Hz 0.949612 -0.283274
+ 3.71e+10Hz 0.949388 -0.284007
+ 3.72e+10Hz 0.949164 -0.284739
+ 3.73e+10Hz 0.948939 -0.285471
+ 3.74e+10Hz 0.948713 -0.286204
+ 3.75e+10Hz 0.948487 -0.286936
+ 3.76e+10Hz 0.948261 -0.287668
+ 3.77e+10Hz 0.948034 -0.2884
+ 3.78e+10Hz 0.947807 -0.289132
+ 3.79e+10Hz 0.947579 -0.289863
+ 3.8e+10Hz 0.947351 -0.290595
+ 3.81e+10Hz 0.947122 -0.291326
+ 3.82e+10Hz 0.946893 -0.292058
+ 3.83e+10Hz 0.946663 -0.292789
+ 3.84e+10Hz 0.946433 -0.29352
+ 3.85e+10Hz 0.946202 -0.294251
+ 3.86e+10Hz 0.945971 -0.294982
+ 3.87e+10Hz 0.945739 -0.295713
+ 3.88e+10Hz 0.945507 -0.296444
+ 3.89e+10Hz 0.945274 -0.297175
+ 3.9e+10Hz 0.945041 -0.297905
+ 3.91e+10Hz 0.944807 -0.298636
+ 3.92e+10Hz 0.944573 -0.299366
+ 3.93e+10Hz 0.944338 -0.300097
+ 3.94e+10Hz 0.944103 -0.300827
+ 3.95e+10Hz 0.943867 -0.301557
+ 3.96e+10Hz 0.94363 -0.302287
+ 3.97e+10Hz 0.943394 -0.303017
+ 3.98e+10Hz 0.943156 -0.303747
+ 3.99e+10Hz 0.942918 -0.304477
+ 4e+10Hz 0.94268 -0.305206
+ 4.01e+10Hz 0.942441 -0.305936
+ 4.02e+10Hz 0.942201 -0.306666
+ 4.03e+10Hz 0.941961 -0.307395
+ 4.04e+10Hz 0.94172 -0.308124
+ 4.05e+10Hz 0.941479 -0.308854
+ 4.06e+10Hz 0.941237 -0.309583
+ 4.07e+10Hz 0.940995 -0.310312
+ 4.08e+10Hz 0.940752 -0.311041
+ 4.09e+10Hz 0.940509 -0.31177
+ 4.1e+10Hz 0.940265 -0.312499
+ 4.11e+10Hz 0.94002 -0.313227
+ 4.12e+10Hz 0.939775 -0.313956
+ 4.13e+10Hz 0.939529 -0.314685
+ 4.14e+10Hz 0.939283 -0.315413
+ 4.15e+10Hz 0.939036 -0.316141
+ 4.16e+10Hz 0.938789 -0.31687
+ 4.17e+10Hz 0.938541 -0.317598
+ 4.18e+10Hz 0.938292 -0.318326
+ 4.19e+10Hz 0.938043 -0.319054
+ 4.2e+10Hz 0.937793 -0.319782
+ 4.21e+10Hz 0.937543 -0.320509
+ 4.22e+10Hz 0.937292 -0.321237
+ 4.23e+10Hz 0.93704 -0.321965
+ 4.24e+10Hz 0.936788 -0.322692
+ 4.25e+10Hz 0.936535 -0.323419
+ 4.26e+10Hz 0.936282 -0.324146
+ 4.27e+10Hz 0.936028 -0.324874
+ 4.28e+10Hz 0.935773 -0.3256
+ 4.29e+10Hz 0.935518 -0.326327
+ 4.3e+10Hz 0.935262 -0.327054
+ 4.31e+10Hz 0.935006 -0.327781
+ 4.32e+10Hz 0.934749 -0.328507
+ 4.33e+10Hz 0.934491 -0.329233
+ 4.34e+10Hz 0.934233 -0.32996
+ 4.35e+10Hz 0.933974 -0.330686
+ 4.36e+10Hz 0.933714 -0.331412
+ 4.37e+10Hz 0.933454 -0.332137
+ 4.38e+10Hz 0.933193 -0.332863
+ 4.39e+10Hz 0.932932 -0.333589
+ 4.4e+10Hz 0.932669 -0.334314
+ 4.41e+10Hz 0.932407 -0.335039
+ 4.42e+10Hz 0.932143 -0.335764
+ 4.43e+10Hz 0.931879 -0.336489
+ 4.44e+10Hz 0.931615 -0.337214
+ 4.45e+10Hz 0.93135 -0.337938
+ 4.46e+10Hz 0.931084 -0.338663
+ 4.47e+10Hz 0.930817 -0.339387
+ 4.48e+10Hz 0.93055 -0.340111
+ 4.49e+10Hz 0.930282 -0.340835
+ 4.5e+10Hz 0.930014 -0.341559
+ 4.51e+10Hz 0.929744 -0.342282
+ 4.52e+10Hz 0.929475 -0.343006
+ 4.53e+10Hz 0.929204 -0.343729
+ 4.54e+10Hz 0.928933 -0.344452
+ 4.55e+10Hz 0.928662 -0.345175
+ 4.56e+10Hz 0.928389 -0.345897
+ 4.57e+10Hz 0.928116 -0.34662
+ 4.58e+10Hz 0.927843 -0.347342
+ 4.59e+10Hz 0.927568 -0.348064
+ 4.6e+10Hz 0.927293 -0.348786
+ 4.61e+10Hz 0.927018 -0.349507
+ 4.62e+10Hz 0.926742 -0.350229
+ 4.63e+10Hz 0.926465 -0.35095
+ 4.64e+10Hz 0.926187 -0.351671
+ 4.65e+10Hz 0.925909 -0.352391
+ 4.66e+10Hz 0.92563 -0.353112
+ 4.67e+10Hz 0.925351 -0.353832
+ 4.68e+10Hz 0.925071 -0.354552
+ 4.69e+10Hz 0.92479 -0.355272
+ 4.7e+10Hz 0.924509 -0.355992
+ 4.71e+10Hz 0.924227 -0.356711
+ 4.72e+10Hz 0.923944 -0.35743
+ 4.73e+10Hz 0.923661 -0.358149
+ 4.74e+10Hz 0.923377 -0.358867
+ 4.75e+10Hz 0.923092 -0.359586
+ 4.76e+10Hz 0.922807 -0.360304
+ 4.77e+10Hz 0.922521 -0.361022
+ 4.78e+10Hz 0.922235 -0.361739
+ 4.79e+10Hz 0.921948 -0.362457
+ 4.8e+10Hz 0.92166 -0.363174
+ 4.81e+10Hz 0.921371 -0.36389
+ 4.82e+10Hz 0.921082 -0.364607
+ 4.83e+10Hz 0.920793 -0.365323
+ 4.84e+10Hz 0.920503 -0.366039
+ 4.85e+10Hz 0.920212 -0.366755
+ 4.86e+10Hz 0.91992 -0.36747
+ 4.87e+10Hz 0.919628 -0.368185
+ 4.88e+10Hz 0.919335 -0.3689
+ 4.89e+10Hz 0.919042 -0.369615
+ 4.9e+10Hz 0.918748 -0.370329
+ 4.91e+10Hz 0.918454 -0.371043
+ 4.92e+10Hz 0.918158 -0.371756
+ 4.93e+10Hz 0.917863 -0.37247
+ 4.94e+10Hz 0.917566 -0.373183
+ 4.95e+10Hz 0.917269 -0.373896
+ 4.96e+10Hz 0.916972 -0.374608
+ 4.97e+10Hz 0.916673 -0.37532
+ 4.98e+10Hz 0.916375 -0.376032
+ 4.99e+10Hz 0.916075 -0.376744
+ 5e+10Hz 0.915775 -0.377455
+ 5.01e+10Hz 0.915475 -0.378166
+ 5.02e+10Hz 0.915174 -0.378877
+ 5.03e+10Hz 0.914872 -0.379587
+ 5.04e+10Hz 0.914569 -0.380297
+ 5.05e+10Hz 0.914267 -0.381007
+ 5.06e+10Hz 0.913963 -0.381716
+ 5.07e+10Hz 0.913659 -0.382425
+ 5.08e+10Hz 0.913354 -0.383134
+ 5.09e+10Hz 0.913049 -0.383842
+ 5.1e+10Hz 0.912743 -0.38455
+ 5.11e+10Hz 0.912437 -0.385258
+ 5.12e+10Hz 0.91213 -0.385966
+ 5.13e+10Hz 0.911823 -0.386673
+ 5.14e+10Hz 0.911515 -0.38738
+ 5.15e+10Hz 0.911206 -0.388086
+ 5.16e+10Hz 0.910897 -0.388792
+ 5.17e+10Hz 0.910587 -0.389498
+ 5.18e+10Hz 0.910277 -0.390204
+ 5.19e+10Hz 0.909967 -0.390909
+ 5.2e+10Hz 0.909655 -0.391614
+ 5.21e+10Hz 0.909343 -0.392318
+ 5.22e+10Hz 0.909031 -0.393023
+ 5.23e+10Hz 0.908718 -0.393726
+ 5.24e+10Hz 0.908405 -0.39443
+ 5.25e+10Hz 0.908091 -0.395133
+ 5.26e+10Hz 0.907776 -0.395836
+ 5.27e+10Hz 0.907461 -0.396539
+ 5.28e+10Hz 0.907146 -0.397241
+ 5.29e+10Hz 0.90683 -0.397943
+ 5.3e+10Hz 0.906513 -0.398645
+ 5.31e+10Hz 0.906196 -0.399346
+ 5.32e+10Hz 0.905878 -0.400047
+ 5.33e+10Hz 0.90556 -0.400748
+ 5.34e+10Hz 0.905242 -0.401448
+ 5.35e+10Hz 0.904922 -0.402148
+ 5.36e+10Hz 0.904603 -0.402848
+ 5.37e+10Hz 0.904283 -0.403547
+ 5.38e+10Hz 0.903962 -0.404246
+ 5.39e+10Hz 0.903641 -0.404945
+ 5.4e+10Hz 0.903319 -0.405643
+ 5.41e+10Hz 0.902997 -0.406341
+ 5.42e+10Hz 0.902675 -0.407039
+ 5.43e+10Hz 0.902351 -0.407737
+ 5.44e+10Hz 0.902028 -0.408434
+ 5.45e+10Hz 0.901704 -0.409131
+ 5.46e+10Hz 0.901379 -0.409827
+ 5.47e+10Hz 0.901054 -0.410523
+ 5.48e+10Hz 0.900729 -0.411219
+ 5.49e+10Hz 0.900403 -0.411915
+ 5.5e+10Hz 0.900076 -0.41261
+ 5.51e+10Hz 0.899749 -0.413305
+ 5.52e+10Hz 0.899422 -0.414
+ 5.53e+10Hz 0.899094 -0.414694
+ 5.54e+10Hz 0.898765 -0.415388
+ 5.55e+10Hz 0.898437 -0.416082
+ 5.56e+10Hz 0.898107 -0.416776
+ 5.57e+10Hz 0.897778 -0.417469
+ 5.58e+10Hz 0.897447 -0.418162
+ 5.59e+10Hz 0.897117 -0.418854
+ 5.6e+10Hz 0.896785 -0.419547
+ 5.61e+10Hz 0.896454 -0.420239
+ 5.62e+10Hz 0.896122 -0.420931
+ 5.63e+10Hz 0.895789 -0.421622
+ 5.64e+10Hz 0.895456 -0.422313
+ 5.65e+10Hz 0.895122 -0.423004
+ 5.66e+10Hz 0.894788 -0.423695
+ 5.67e+10Hz 0.894454 -0.424385
+ 5.68e+10Hz 0.894119 -0.425075
+ 5.69e+10Hz 0.893784 -0.425765
+ 5.7e+10Hz 0.893448 -0.426455
+ 5.71e+10Hz 0.893112 -0.427144
+ 5.72e+10Hz 0.892775 -0.427833
+ 5.73e+10Hz 0.892438 -0.428522
+ 5.74e+10Hz 0.8921 -0.42921
+ 5.75e+10Hz 0.891762 -0.429898
+ 5.76e+10Hz 0.891424 -0.430586
+ 5.77e+10Hz 0.891085 -0.431274
+ 5.78e+10Hz 0.890745 -0.431961
+ 5.79e+10Hz 0.890405 -0.432648
+ 5.8e+10Hz 0.890065 -0.433335
+ 5.81e+10Hz 0.889724 -0.434022
+ 5.82e+10Hz 0.889383 -0.434708
+ 5.83e+10Hz 0.889041 -0.435394
+ 5.84e+10Hz 0.888699 -0.43608
+ 5.85e+10Hz 0.888356 -0.436766
+ 5.86e+10Hz 0.888013 -0.437451
+ 5.87e+10Hz 0.887669 -0.438137
+ 5.88e+10Hz 0.887325 -0.438821
+ 5.89e+10Hz 0.886981 -0.439506
+ 5.9e+10Hz 0.886636 -0.440191
+ 5.91e+10Hz 0.88629 -0.440875
+ 5.92e+10Hz 0.885944 -0.441559
+ 5.93e+10Hz 0.885598 -0.442242
+ 5.94e+10Hz 0.885251 -0.442926
+ 5.95e+10Hz 0.884904 -0.443609
+ 5.96e+10Hz 0.884556 -0.444292
+ 5.97e+10Hz 0.884208 -0.444975
+ 5.98e+10Hz 0.883859 -0.445658
+ 5.99e+10Hz 0.88351 -0.44634
+ 6e+10Hz 0.88316 -0.447022
+ 6.01e+10Hz 0.88281 -0.447704
+ 6.02e+10Hz 0.88246 -0.448385
+ 6.03e+10Hz 0.882108 -0.449067
+ 6.04e+10Hz 0.881757 -0.449748
+ 6.05e+10Hz 0.881405 -0.450429
+ 6.06e+10Hz 0.881052 -0.45111
+ 6.07e+10Hz 0.880699 -0.45179
+ 6.08e+10Hz 0.880346 -0.452471
+ 6.09e+10Hz 0.879992 -0.453151
+ 6.1e+10Hz 0.879637 -0.453831
+ 6.11e+10Hz 0.879282 -0.45451
+ 6.12e+10Hz 0.878927 -0.45519
+ 6.13e+10Hz 0.878571 -0.455869
+ 6.14e+10Hz 0.878215 -0.456548
+ 6.15e+10Hz 0.877858 -0.457227
+ 6.16e+10Hz 0.8775 -0.457905
+ 6.17e+10Hz 0.877142 -0.458584
+ 6.18e+10Hz 0.876784 -0.459262
+ 6.19e+10Hz 0.876425 -0.45994
+ 6.2e+10Hz 0.876066 -0.460618
+ 6.21e+10Hz 0.875706 -0.461295
+ 6.22e+10Hz 0.875345 -0.461972
+ 6.23e+10Hz 0.874984 -0.462649
+ 6.24e+10Hz 0.874623 -0.463326
+ 6.25e+10Hz 0.874261 -0.464003
+ 6.26e+10Hz 0.873899 -0.464679
+ 6.27e+10Hz 0.873536 -0.465356
+ 6.28e+10Hz 0.873172 -0.466032
+ 6.29e+10Hz 0.872808 -0.466707
+ 6.3e+10Hz 0.872444 -0.467383
+ 6.31e+10Hz 0.872079 -0.468058
+ 6.32e+10Hz 0.871713 -0.468734
+ 6.33e+10Hz 0.871347 -0.469408
+ 6.34e+10Hz 0.87098 -0.470083
+ 6.35e+10Hz 0.870613 -0.470758
+ 6.36e+10Hz 0.870245 -0.471432
+ 6.37e+10Hz 0.869877 -0.472106
+ 6.38e+10Hz 0.869508 -0.47278
+ 6.39e+10Hz 0.869139 -0.473453
+ 6.4e+10Hz 0.868769 -0.474127
+ 6.41e+10Hz 0.868399 -0.4748
+ 6.42e+10Hz 0.868028 -0.475473
+ 6.43e+10Hz 0.867657 -0.476145
+ 6.44e+10Hz 0.867285 -0.476818
+ 6.45e+10Hz 0.866912 -0.47749
+ 6.46e+10Hz 0.866539 -0.478162
+ 6.47e+10Hz 0.866165 -0.478834
+ 6.48e+10Hz 0.865791 -0.479506
+ 6.49e+10Hz 0.865416 -0.480177
+ 6.5e+10Hz 0.865041 -0.480848
+ 6.51e+10Hz 0.864665 -0.481519
+ 6.52e+10Hz 0.864289 -0.482189
+ 6.53e+10Hz 0.863912 -0.48286
+ 6.54e+10Hz 0.863534 -0.48353
+ 6.55e+10Hz 0.863156 -0.4842
+ 6.56e+10Hz 0.862778 -0.484869
+ 6.57e+10Hz 0.862399 -0.485539
+ 6.58e+10Hz 0.862019 -0.486208
+ 6.59e+10Hz 0.861639 -0.486877
+ 6.6e+10Hz 0.861258 -0.487546
+ 6.61e+10Hz 0.860876 -0.488214
+ 6.62e+10Hz 0.860494 -0.488882
+ 6.63e+10Hz 0.860112 -0.48955
+ 6.64e+10Hz 0.859729 -0.490218
+ 6.65e+10Hz 0.859345 -0.490885
+ 6.66e+10Hz 0.858961 -0.491552
+ 6.67e+10Hz 0.858576 -0.492219
+ 6.68e+10Hz 0.85819 -0.492886
+ 6.69e+10Hz 0.857804 -0.493552
+ 6.7e+10Hz 0.857418 -0.494218
+ 6.71e+10Hz 0.857031 -0.494884
+ 6.72e+10Hz 0.856643 -0.495549
+ 6.73e+10Hz 0.856255 -0.496214
+ 6.74e+10Hz 0.855866 -0.496879
+ 6.75e+10Hz 0.855476 -0.497544
+ 6.76e+10Hz 0.855086 -0.498208
+ 6.77e+10Hz 0.854696 -0.498872
+ 6.78e+10Hz 0.854305 -0.499536
+ 6.79e+10Hz 0.853913 -0.5002
+ 6.8e+10Hz 0.853521 -0.500863
+ 6.81e+10Hz 0.853128 -0.501526
+ 6.82e+10Hz 0.852734 -0.502189
+ 6.83e+10Hz 0.85234 -0.502851
+ 6.84e+10Hz 0.851946 -0.503513
+ 6.85e+10Hz 0.851551 -0.504175
+ 6.86e+10Hz 0.851155 -0.504836
+ 6.87e+10Hz 0.850759 -0.505497
+ 6.88e+10Hz 0.850362 -0.506158
+ 6.89e+10Hz 0.849964 -0.506819
+ 6.9e+10Hz 0.849566 -0.507479
+ 6.91e+10Hz 0.849168 -0.508139
+ 6.92e+10Hz 0.848768 -0.508798
+ 6.93e+10Hz 0.848369 -0.509457
+ 6.94e+10Hz 0.847968 -0.510116
+ 6.95e+10Hz 0.847567 -0.510775
+ 6.96e+10Hz 0.847166 -0.511433
+ 6.97e+10Hz 0.846764 -0.512091
+ 6.98e+10Hz 0.846361 -0.512749
+ 6.99e+10Hz 0.845958 -0.513406
+ 7e+10Hz 0.845554 -0.514063
+ 7.01e+10Hz 0.84515 -0.51472
+ 7.02e+10Hz 0.844745 -0.515376
+ 7.03e+10Hz 0.84434 -0.516032
+ 7.04e+10Hz 0.843934 -0.516687
+ 7.05e+10Hz 0.843527 -0.517343
+ 7.06e+10Hz 0.84312 -0.517998
+ 7.07e+10Hz 0.842712 -0.518652
+ 7.08e+10Hz 0.842304 -0.519306
+ 7.09e+10Hz 0.841895 -0.51996
+ 7.1e+10Hz 0.841486 -0.520614
+ 7.11e+10Hz 0.841076 -0.521267
+ 7.12e+10Hz 0.840665 -0.52192
+ 7.13e+10Hz 0.840254 -0.522572
+ 7.14e+10Hz 0.839843 -0.523224
+ 7.15e+10Hz 0.83943 -0.523876
+ 7.16e+10Hz 0.839018 -0.524527
+ 7.17e+10Hz 0.838605 -0.525178
+ 7.18e+10Hz 0.838191 -0.525829
+ 7.19e+10Hz 0.837776 -0.526479
+ 7.2e+10Hz 0.837362 -0.527129
+ 7.21e+10Hz 0.836946 -0.527779
+ 7.22e+10Hz 0.83653 -0.528428
+ 7.23e+10Hz 0.836114 -0.529077
+ 7.24e+10Hz 0.835697 -0.529725
+ 7.25e+10Hz 0.835279 -0.530373
+ 7.26e+10Hz 0.834861 -0.531021
+ 7.27e+10Hz 0.834442 -0.531668
+ 7.28e+10Hz 0.834023 -0.532315
+ 7.29e+10Hz 0.833604 -0.532961
+ 7.3e+10Hz 0.833183 -0.533608
+ 7.31e+10Hz 0.832763 -0.534253
+ 7.32e+10Hz 0.832341 -0.534899
+ 7.33e+10Hz 0.83192 -0.535544
+ 7.34e+10Hz 0.831497 -0.536188
+ 7.35e+10Hz 0.831075 -0.536833
+ 7.36e+10Hz 0.830651 -0.537476
+ 7.37e+10Hz 0.830227 -0.53812
+ 7.38e+10Hz 0.829803 -0.538763
+ 7.39e+10Hz 0.829378 -0.539406
+ 7.4e+10Hz 0.828953 -0.540048
+ 7.41e+10Hz 0.828527 -0.54069
+ 7.42e+10Hz 0.828101 -0.541331
+ 7.43e+10Hz 0.827674 -0.541972
+ 7.44e+10Hz 0.827246 -0.542613
+ 7.45e+10Hz 0.826818 -0.543254
+ 7.46e+10Hz 0.82639 -0.543894
+ 7.47e+10Hz 0.825961 -0.544533
+ 7.48e+10Hz 0.825532 -0.545172
+ 7.49e+10Hz 0.825102 -0.545811
+ 7.5e+10Hz 0.824672 -0.546449
+ 7.51e+10Hz 0.824241 -0.547087
+ 7.52e+10Hz 0.82381 -0.547725
+ 7.53e+10Hz 0.823378 -0.548362
+ 7.54e+10Hz 0.822946 -0.548999
+ 7.55e+10Hz 0.822513 -0.549636
+ 7.56e+10Hz 0.82208 -0.550272
+ 7.57e+10Hz 0.821646 -0.550907
+ 7.58e+10Hz 0.821212 -0.551542
+ 7.59e+10Hz 0.820777 -0.552177
+ 7.6e+10Hz 0.820342 -0.552812
+ 7.61e+10Hz 0.819906 -0.553446
+ 7.62e+10Hz 0.81947 -0.55408
+ 7.63e+10Hz 0.819034 -0.554713
+ 7.64e+10Hz 0.818597 -0.555346
+ 7.65e+10Hz 0.818159 -0.555978
+ 7.66e+10Hz 0.817721 -0.556611
+ 7.67e+10Hz 0.817283 -0.557242
+ 7.68e+10Hz 0.816844 -0.557874
+ 7.69e+10Hz 0.816405 -0.558505
+ 7.7e+10Hz 0.815965 -0.559135
+ 7.71e+10Hz 0.815525 -0.559765
+ 7.72e+10Hz 0.815084 -0.560395
+ 7.73e+10Hz 0.814643 -0.561025
+ 7.74e+10Hz 0.814202 -0.561654
+ 7.75e+10Hz 0.81376 -0.562282
+ 7.76e+10Hz 0.813317 -0.562911
+ 7.77e+10Hz 0.812874 -0.563539
+ 7.78e+10Hz 0.812431 -0.564166
+ 7.79e+10Hz 0.811987 -0.564793
+ 7.8e+10Hz 0.811543 -0.56542
+ 7.81e+10Hz 0.811098 -0.566047
+ 7.82e+10Hz 0.810653 -0.566673
+ 7.83e+10Hz 0.810208 -0.567298
+ 7.84e+10Hz 0.809762 -0.567924
+ 7.85e+10Hz 0.809315 -0.568549
+ 7.86e+10Hz 0.808868 -0.569173
+ 7.87e+10Hz 0.808421 -0.569797
+ 7.88e+10Hz 0.807973 -0.570421
+ 7.89e+10Hz 0.807525 -0.571044
+ 7.9e+10Hz 0.807076 -0.571668
+ 7.91e+10Hz 0.806627 -0.57229
+ 7.92e+10Hz 0.806178 -0.572913
+ 7.93e+10Hz 0.805728 -0.573535
+ 7.94e+10Hz 0.805278 -0.574156
+ 7.95e+10Hz 0.804827 -0.574777
+ 7.96e+10Hz 0.804376 -0.575398
+ 7.97e+10Hz 0.803924 -0.576019
+ 7.98e+10Hz 0.803472 -0.576639
+ 7.99e+10Hz 0.80302 -0.577259
+ 8e+10Hz 0.802567 -0.577878
+ 8.01e+10Hz 0.802113 -0.578497
+ 8.02e+10Hz 0.80166 -0.579116
+ 8.03e+10Hz 0.801205 -0.579734
+ 8.04e+10Hz 0.800751 -0.580352
+ 8.05e+10Hz 0.800296 -0.58097
+ 8.06e+10Hz 0.79984 -0.581587
+ 8.07e+10Hz 0.799384 -0.582204
+ 8.08e+10Hz 0.798928 -0.582821
+ 8.09e+10Hz 0.798471 -0.583437
+ 8.1e+10Hz 0.798014 -0.584053
+ 8.11e+10Hz 0.797556 -0.584669
+ 8.12e+10Hz 0.797098 -0.585284
+ 8.13e+10Hz 0.79664 -0.585899
+ 8.14e+10Hz 0.796181 -0.586514
+ 8.15e+10Hz 0.795721 -0.587128
+ 8.16e+10Hz 0.795262 -0.587742
+ 8.17e+10Hz 0.794801 -0.588355
+ 8.18e+10Hz 0.794341 -0.588969
+ 8.19e+10Hz 0.79388 -0.589581
+ 8.2e+10Hz 0.793418 -0.590194
+ 8.21e+10Hz 0.792956 -0.590806
+ 8.22e+10Hz 0.792494 -0.591418
+ 8.23e+10Hz 0.792031 -0.59203
+ 8.24e+10Hz 0.791568 -0.592641
+ 8.25e+10Hz 0.791104 -0.593252
+ 8.26e+10Hz 0.79064 -0.593862
+ 8.27e+10Hz 0.790176 -0.594472
+ 8.28e+10Hz 0.789711 -0.595082
+ 8.29e+10Hz 0.789245 -0.595692
+ 8.3e+10Hz 0.788779 -0.596301
+ 8.31e+10Hz 0.788313 -0.59691
+ 8.32e+10Hz 0.787846 -0.597518
+ 8.33e+10Hz 0.787379 -0.598127
+ 8.34e+10Hz 0.786912 -0.598735
+ 8.35e+10Hz 0.786444 -0.599342
+ 8.36e+10Hz 0.785975 -0.599949
+ 8.37e+10Hz 0.785506 -0.600556
+ 8.38e+10Hz 0.785037 -0.601163
+ 8.39e+10Hz 0.784567 -0.601769
+ 8.4e+10Hz 0.784097 -0.602375
+ 8.41e+10Hz 0.783626 -0.602981
+ 8.42e+10Hz 0.783155 -0.603586
+ 8.43e+10Hz 0.782683 -0.604191
+ 8.44e+10Hz 0.782211 -0.604796
+ 8.45e+10Hz 0.781739 -0.6054
+ 8.46e+10Hz 0.781266 -0.606004
+ 8.47e+10Hz 0.780792 -0.606608
+ 8.48e+10Hz 0.780319 -0.607211
+ 8.49e+10Hz 0.779844 -0.607814
+ 8.5e+10Hz 0.779369 -0.608417
+ 8.51e+10Hz 0.778894 -0.609019
+ 8.52e+10Hz 0.778419 -0.609621
+ 8.53e+10Hz 0.777942 -0.610223
+ 8.54e+10Hz 0.777466 -0.610825
+ 8.55e+10Hz 0.776989 -0.611426
+ 8.56e+10Hz 0.776511 -0.612026
+ 8.57e+10Hz 0.776033 -0.612627
+ 8.58e+10Hz 0.775555 -0.613227
+ 8.59e+10Hz 0.775076 -0.613827
+ 8.6e+10Hz 0.774596 -0.614426
+ 8.61e+10Hz 0.774117 -0.615025
+ 8.62e+10Hz 0.773636 -0.615624
+ 8.63e+10Hz 0.773155 -0.616223
+ 8.64e+10Hz 0.772674 -0.616821
+ 8.65e+10Hz 0.772192 -0.617419
+ 8.66e+10Hz 0.77171 -0.618016
+ 8.67e+10Hz 0.771228 -0.618614
+ 8.68e+10Hz 0.770744 -0.61921
+ 8.69e+10Hz 0.770261 -0.619807
+ 8.7e+10Hz 0.769777 -0.620403
+ 8.71e+10Hz 0.769292 -0.620999
+ 8.72e+10Hz 0.768807 -0.621594
+ 8.73e+10Hz 0.768321 -0.62219
+ 8.74e+10Hz 0.767835 -0.622784
+ 8.75e+10Hz 0.767349 -0.623379
+ 8.76e+10Hz 0.766862 -0.623973
+ 8.77e+10Hz 0.766374 -0.624567
+ 8.78e+10Hz 0.765886 -0.625161
+ 8.79e+10Hz 0.765398 -0.625754
+ 8.8e+10Hz 0.764909 -0.626346
+ 8.81e+10Hz 0.76442 -0.626939
+ 8.82e+10Hz 0.76393 -0.627531
+ 8.83e+10Hz 0.763439 -0.628123
+ 8.84e+10Hz 0.762948 -0.628714
+ 8.85e+10Hz 0.762457 -0.629305
+ 8.86e+10Hz 0.761965 -0.629896
+ 8.87e+10Hz 0.761473 -0.630487
+ 8.88e+10Hz 0.76098 -0.631077
+ 8.89e+10Hz 0.760487 -0.631666
+ 8.9e+10Hz 0.759993 -0.632256
+ 8.91e+10Hz 0.759499 -0.632845
+ 8.92e+10Hz 0.759004 -0.633433
+ 8.93e+10Hz 0.758508 -0.634021
+ 8.94e+10Hz 0.758013 -0.634609
+ 8.95e+10Hz 0.757516 -0.635197
+ 8.96e+10Hz 0.757019 -0.635784
+ 8.97e+10Hz 0.756522 -0.636371
+ 8.98e+10Hz 0.756024 -0.636957
+ 8.99e+10Hz 0.755526 -0.637543
+ 9e+10Hz 0.755027 -0.638129
+ 9.01e+10Hz 0.754528 -0.638715
+ 9.02e+10Hz 0.754028 -0.639299
+ 9.03e+10Hz 0.753528 -0.639884
+ 9.04e+10Hz 0.753027 -0.640468
+ 9.05e+10Hz 0.752526 -0.641052
+ 9.06e+10Hz 0.752024 -0.641636
+ 9.07e+10Hz 0.751522 -0.642219
+ 9.08e+10Hz 0.751019 -0.642801
+ 9.09e+10Hz 0.750516 -0.643384
+ 9.1e+10Hz 0.750012 -0.643966
+ 9.11e+10Hz 0.749508 -0.644547
+ 9.12e+10Hz 0.749003 -0.645128
+ 9.13e+10Hz 0.748498 -0.645709
+ 9.14e+10Hz 0.747992 -0.64629
+ 9.15e+10Hz 0.747486 -0.64687
+ 9.16e+10Hz 0.74698 -0.647449
+ 9.17e+10Hz 0.746472 -0.648028
+ 9.18e+10Hz 0.745965 -0.648607
+ 9.19e+10Hz 0.745456 -0.649186
+ 9.2e+10Hz 0.744948 -0.649764
+ 9.21e+10Hz 0.744439 -0.650341
+ 9.22e+10Hz 0.743929 -0.650919
+ 9.23e+10Hz 0.743419 -0.651495
+ 9.24e+10Hz 0.742908 -0.652072
+ 9.25e+10Hz 0.742397 -0.652648
+ 9.26e+10Hz 0.741885 -0.653223
+ 9.27e+10Hz 0.741373 -0.653799
+ 9.28e+10Hz 0.740861 -0.654373
+ 9.29e+10Hz 0.740347 -0.654948
+ 9.3e+10Hz 0.739834 -0.655522
+ 9.31e+10Hz 0.73932 -0.656095
+ 9.32e+10Hz 0.738805 -0.656668
+ 9.33e+10Hz 0.73829 -0.657241
+ 9.34e+10Hz 0.737775 -0.657813
+ 9.35e+10Hz 0.737259 -0.658385
+ 9.36e+10Hz 0.736742 -0.658956
+ 9.37e+10Hz 0.736225 -0.659527
+ 9.38e+10Hz 0.735708 -0.660098
+ 9.39e+10Hz 0.73519 -0.660668
+ 9.4e+10Hz 0.734671 -0.661238
+ 9.41e+10Hz 0.734153 -0.661807
+ 9.42e+10Hz 0.733633 -0.662376
+ 9.43e+10Hz 0.733113 -0.662944
+ 9.44e+10Hz 0.732593 -0.663512
+ 9.45e+10Hz 0.732072 -0.66408
+ 9.46e+10Hz 0.731551 -0.664647
+ 9.47e+10Hz 0.731029 -0.665214
+ 9.48e+10Hz 0.730507 -0.66578
+ 9.49e+10Hz 0.729984 -0.666346
+ 9.5e+10Hz 0.729461 -0.666911
+ 9.51e+10Hz 0.728938 -0.667476
+ 9.52e+10Hz 0.728414 -0.66804
+ 9.53e+10Hz 0.727889 -0.668605
+ 9.54e+10Hz 0.727364 -0.669168
+ 9.55e+10Hz 0.726839 -0.669731
+ 9.56e+10Hz 0.726313 -0.670294
+ 9.57e+10Hz 0.725787 -0.670856
+ 9.58e+10Hz 0.72526 -0.671418
+ 9.59e+10Hz 0.724733 -0.671979
+ 9.6e+10Hz 0.724205 -0.67254
+ 9.61e+10Hz 0.723677 -0.673101
+ 9.62e+10Hz 0.723148 -0.673661
+ 9.63e+10Hz 0.722619 -0.67422
+ 9.64e+10Hz 0.72209 -0.674779
+ 9.65e+10Hz 0.72156 -0.675338
+ 9.66e+10Hz 0.721029 -0.675896
+ 9.67e+10Hz 0.720498 -0.676454
+ 9.68e+10Hz 0.719967 -0.677011
+ 9.69e+10Hz 0.719436 -0.677568
+ 9.7e+10Hz 0.718903 -0.678125
+ 9.71e+10Hz 0.718371 -0.678681
+ 9.72e+10Hz 0.717838 -0.679236
+ 9.73e+10Hz 0.717304 -0.679791
+ 9.74e+10Hz 0.71677 -0.680346
+ 9.75e+10Hz 0.716236 -0.6809
+ 9.76e+10Hz 0.715701 -0.681453
+ 9.77e+10Hz 0.715166 -0.682007
+ 9.78e+10Hz 0.714631 -0.682559
+ 9.79e+10Hz 0.714095 -0.683112
+ 9.8e+10Hz 0.713558 -0.683664
+ 9.81e+10Hz 0.713021 -0.684215
+ 9.82e+10Hz 0.712484 -0.684766
+ 9.83e+10Hz 0.711946 -0.685316
+ 9.84e+10Hz 0.711408 -0.685866
+ 9.85e+10Hz 0.71087 -0.686416
+ 9.86e+10Hz 0.710331 -0.686965
+ 9.87e+10Hz 0.709791 -0.687514
+ 9.88e+10Hz 0.709252 -0.688062
+ 9.89e+10Hz 0.708712 -0.68861
+ 9.9e+10Hz 0.708171 -0.689157
+ 9.91e+10Hz 0.70763 -0.689704
+ 9.92e+10Hz 0.707089 -0.69025
+ 9.93e+10Hz 0.706547 -0.690796
+ 9.94e+10Hz 0.706004 -0.691342
+ 9.95e+10Hz 0.705462 -0.691887
+ 9.96e+10Hz 0.704919 -0.692431
+ 9.97e+10Hz 0.704375 -0.692975
+ 9.98e+10Hz 0.703832 -0.693519
+ 9.99e+10Hz 0.703287 -0.694062
+ 1e+11Hz 0.702743 -0.694605
+ 1.001e+11Hz 0.702198 -0.695147
+ 1.002e+11Hz 0.701652 -0.695689
+ 1.003e+11Hz 0.701106 -0.696231
+ 1.004e+11Hz 0.70056 -0.696772
+ 1.005e+11Hz 0.700014 -0.697312
+ 1.006e+11Hz 0.699467 -0.697852
+ 1.007e+11Hz 0.698919 -0.698392
+ 1.008e+11Hz 0.698372 -0.698931
+ 1.009e+11Hz 0.697823 -0.69947
+ 1.01e+11Hz 0.697275 -0.700008
+ 1.011e+11Hz 0.696726 -0.700546
+ 1.012e+11Hz 0.696177 -0.701083
+ 1.013e+11Hz 0.695627 -0.70162
+ 1.014e+11Hz 0.695077 -0.702157
+ 1.015e+11Hz 0.694526 -0.702693
+ 1.016e+11Hz 0.693975 -0.703229
+ 1.017e+11Hz 0.693424 -0.703764
+ 1.018e+11Hz 0.692873 -0.704299
+ 1.019e+11Hz 0.692321 -0.704833
+ 1.02e+11Hz 0.691768 -0.705367
+ 1.021e+11Hz 0.691215 -0.7059
+ 1.022e+11Hz 0.690662 -0.706433
+ 1.023e+11Hz 0.690109 -0.706966
+ 1.024e+11Hz 0.689555 -0.707498
+ 1.025e+11Hz 0.689 -0.70803
+ 1.026e+11Hz 0.688446 -0.708561
+ 1.027e+11Hz 0.687891 -0.709092
+ 1.028e+11Hz 0.687335 -0.709622
+ 1.029e+11Hz 0.686779 -0.710152
+ 1.03e+11Hz 0.686223 -0.710682
+ 1.031e+11Hz 0.685667 -0.711211
+ 1.032e+11Hz 0.68511 -0.71174
+ 1.033e+11Hz 0.684552 -0.712268
+ 1.034e+11Hz 0.683995 -0.712796
+ 1.035e+11Hz 0.683437 -0.713323
+ 1.036e+11Hz 0.682878 -0.71385
+ 1.037e+11Hz 0.682319 -0.714377
+ 1.038e+11Hz 0.68176 -0.714903
+ 1.039e+11Hz 0.681201 -0.715428
+ 1.04e+11Hz 0.680641 -0.715954
+ 1.041e+11Hz 0.68008 -0.716479
+ 1.042e+11Hz 0.67952 -0.717003
+ 1.043e+11Hz 0.678958 -0.717527
+ 1.044e+11Hz 0.678397 -0.718051
+ 1.045e+11Hz 0.677835 -0.718574
+ 1.046e+11Hz 0.677273 -0.719097
+ 1.047e+11Hz 0.67671 -0.719619
+ 1.048e+11Hz 0.676147 -0.720141
+ 1.049e+11Hz 0.675584 -0.720662
+ 1.05e+11Hz 0.67502 -0.721183
+ 1.051e+11Hz 0.674456 -0.721704
+ 1.052e+11Hz 0.673891 -0.722224
+ 1.053e+11Hz 0.673327 -0.722744
+ 1.054e+11Hz 0.672761 -0.723264
+ 1.055e+11Hz 0.672196 -0.723783
+ 1.056e+11Hz 0.67163 -0.724301
+ 1.057e+11Hz 0.671063 -0.72482
+ 1.058e+11Hz 0.670496 -0.725337
+ 1.059e+11Hz 0.669929 -0.725855
+ 1.06e+11Hz 0.669362 -0.726372
+ 1.061e+11Hz 0.668794 -0.726888
+ 1.062e+11Hz 0.668225 -0.727404
+ 1.063e+11Hz 0.667657 -0.72792
+ 1.064e+11Hz 0.667087 -0.728435
+ 1.065e+11Hz 0.666518 -0.72895
+ 1.066e+11Hz 0.665948 -0.729465
+ 1.067e+11Hz 0.665378 -0.729979
+ 1.068e+11Hz 0.664807 -0.730493
+ 1.069e+11Hz 0.664236 -0.731006
+ 1.07e+11Hz 0.663665 -0.731519
+ 1.071e+11Hz 0.663093 -0.732031
+ 1.072e+11Hz 0.662521 -0.732543
+ 1.073e+11Hz 0.661948 -0.733055
+ 1.074e+11Hz 0.661375 -0.733566
+ 1.075e+11Hz 0.660801 -0.734077
+ 1.076e+11Hz 0.660228 -0.734587
+ 1.077e+11Hz 0.659653 -0.735097
+ 1.078e+11Hz 0.659079 -0.735607
+ 1.079e+11Hz 0.658504 -0.736116
+ 1.08e+11Hz 0.657928 -0.736625
+ 1.081e+11Hz 0.657353 -0.737133
+ 1.082e+11Hz 0.656776 -0.737641
+ 1.083e+11Hz 0.6562 -0.738148
+ 1.084e+11Hz 0.655623 -0.738655
+ 1.085e+11Hz 0.655045 -0.739162
+ 1.086e+11Hz 0.654468 -0.739668
+ 1.087e+11Hz 0.653889 -0.740174
+ 1.088e+11Hz 0.653311 -0.74068
+ 1.089e+11Hz 0.652732 -0.741185
+ 1.09e+11Hz 0.652152 -0.741689
+ 1.091e+11Hz 0.651573 -0.742194
+ 1.092e+11Hz 0.650992 -0.742697
+ 1.093e+11Hz 0.650412 -0.743201
+ 1.094e+11Hz 0.649831 -0.743704
+ 1.095e+11Hz 0.649249 -0.744206
+ 1.096e+11Hz 0.648667 -0.744708
+ 1.097e+11Hz 0.648085 -0.74521
+ 1.098e+11Hz 0.647502 -0.745711
+ 1.099e+11Hz 0.646919 -0.746212
+ 1.1e+11Hz 0.646336 -0.746713
+ 1.101e+11Hz 0.645752 -0.747213
+ 1.102e+11Hz 0.645167 -0.747712
+ 1.103e+11Hz 0.644583 -0.748212
+ 1.104e+11Hz 0.643998 -0.74871
+ 1.105e+11Hz 0.643412 -0.749209
+ 1.106e+11Hz 0.642826 -0.749706
+ 1.107e+11Hz 0.64224 -0.750204
+ 1.108e+11Hz 0.641653 -0.750701
+ 1.109e+11Hz 0.641065 -0.751198
+ 1.11e+11Hz 0.640478 -0.751694
+ 1.111e+11Hz 0.63989 -0.75219
+ 1.112e+11Hz 0.639301 -0.752685
+ 1.113e+11Hz 0.638712 -0.75318
+ 1.114e+11Hz 0.638123 -0.753674
+ 1.115e+11Hz 0.637533 -0.754168
+ 1.116e+11Hz 0.636943 -0.754662
+ 1.117e+11Hz 0.636352 -0.755155
+ 1.118e+11Hz 0.635761 -0.755648
+ 1.119e+11Hz 0.63517 -0.75614
+ 1.12e+11Hz 0.634578 -0.756632
+ 1.121e+11Hz 0.633986 -0.757123
+ 1.122e+11Hz 0.633393 -0.757614
+ 1.123e+11Hz 0.6328 -0.758105
+ 1.124e+11Hz 0.632206 -0.758595
+ 1.125e+11Hz 0.631612 -0.759084
+ 1.126e+11Hz 0.631018 -0.759573
+ 1.127e+11Hz 0.630423 -0.760062
+ 1.128e+11Hz 0.629828 -0.76055
+ 1.129e+11Hz 0.629232 -0.761038
+ 1.13e+11Hz 0.628636 -0.761526
+ 1.131e+11Hz 0.628039 -0.762012
+ 1.132e+11Hz 0.627442 -0.762499
+ 1.133e+11Hz 0.626845 -0.762985
+ 1.134e+11Hz 0.626247 -0.76347
+ 1.135e+11Hz 0.625649 -0.763955
+ 1.136e+11Hz 0.62505 -0.76444
+ 1.137e+11Hz 0.624451 -0.764924
+ 1.138e+11Hz 0.623852 -0.765408
+ 1.139e+11Hz 0.623252 -0.765891
+ 1.14e+11Hz 0.622651 -0.766374
+ 1.141e+11Hz 0.622051 -0.766856
+ 1.142e+11Hz 0.621449 -0.767338
+ 1.143e+11Hz 0.620848 -0.767819
+ 1.144e+11Hz 0.620246 -0.7683
+ 1.145e+11Hz 0.619643 -0.76878
+ 1.146e+11Hz 0.61904 -0.76926
+ 1.147e+11Hz 0.618437 -0.76974
+ 1.148e+11Hz 0.617833 -0.770218
+ 1.149e+11Hz 0.617229 -0.770697
+ 1.15e+11Hz 0.616625 -0.771175
+ 1.151e+11Hz 0.61602 -0.771652
+ 1.152e+11Hz 0.615414 -0.772129
+ 1.153e+11Hz 0.614808 -0.772606
+ 1.154e+11Hz 0.614202 -0.773082
+ 1.155e+11Hz 0.613596 -0.773557
+ 1.156e+11Hz 0.612989 -0.774032
+ 1.157e+11Hz 0.612381 -0.774507
+ 1.158e+11Hz 0.611773 -0.774981
+ 1.159e+11Hz 0.611165 -0.775455
+ 1.16e+11Hz 0.610556 -0.775928
+ 1.161e+11Hz 0.609947 -0.7764
+ 1.162e+11Hz 0.609338 -0.776872
+ 1.163e+11Hz 0.608728 -0.777344
+ 1.164e+11Hz 0.608117 -0.777815
+ 1.165e+11Hz 0.607507 -0.778286
+ 1.166e+11Hz 0.606895 -0.778756
+ 1.167e+11Hz 0.606284 -0.779225
+ 1.168e+11Hz 0.605672 -0.779694
+ 1.169e+11Hz 0.60506 -0.780163
+ 1.17e+11Hz 0.604447 -0.780631
+ 1.171e+11Hz 0.603834 -0.781099
+ 1.172e+11Hz 0.60322 -0.781566
+ 1.173e+11Hz 0.602606 -0.782032
+ 1.174e+11Hz 0.601992 -0.782498
+ 1.175e+11Hz 0.601377 -0.782964
+ 1.176e+11Hz 0.600762 -0.783429
+ 1.177e+11Hz 0.600146 -0.783893
+ 1.178e+11Hz 0.59953 -0.784357
+ 1.179e+11Hz 0.598914 -0.784821
+ 1.18e+11Hz 0.598297 -0.785284
+ 1.181e+11Hz 0.59768 -0.785746
+ 1.182e+11Hz 0.597063 -0.786208
+ 1.183e+11Hz 0.596445 -0.786669
+ 1.184e+11Hz 0.595827 -0.78713
+ 1.185e+11Hz 0.595208 -0.78759
+ 1.186e+11Hz 0.594589 -0.78805
+ 1.187e+11Hz 0.593969 -0.78851
+ 1.188e+11Hz 0.59335 -0.788968
+ 1.189e+11Hz 0.592729 -0.789427
+ 1.19e+11Hz 0.592109 -0.789884
+ 1.191e+11Hz 0.591488 -0.790342
+ 1.192e+11Hz 0.590867 -0.790798
+ 1.193e+11Hz 0.590245 -0.791254
+ 1.194e+11Hz 0.589623 -0.79171
+ 1.195e+11Hz 0.589001 -0.792165
+ 1.196e+11Hz 0.588378 -0.79262
+ 1.197e+11Hz 0.587755 -0.793074
+ 1.198e+11Hz 0.587131 -0.793527
+ 1.199e+11Hz 0.586507 -0.79398
+ 1.2e+11Hz 0.585883 -0.794433
+ 1.201e+11Hz 0.585258 -0.794885
+ 1.202e+11Hz 0.584633 -0.795336
+ 1.203e+11Hz 0.584008 -0.795787
+ 1.204e+11Hz 0.583382 -0.796237
+ 1.205e+11Hz 0.582756 -0.796687
+ 1.206e+11Hz 0.58213 -0.797137
+ 1.207e+11Hz 0.581503 -0.797585
+ 1.208e+11Hz 0.580876 -0.798033
+ 1.209e+11Hz 0.580248 -0.798481
+ 1.21e+11Hz 0.579621 -0.798928
+ 1.211e+11Hz 0.578993 -0.799375
+ 1.212e+11Hz 0.578364 -0.799821
+ 1.213e+11Hz 0.577735 -0.800267
+ 1.214e+11Hz 0.577106 -0.800712
+ 1.215e+11Hz 0.576476 -0.801156
+ 1.216e+11Hz 0.575846 -0.8016
+ 1.217e+11Hz 0.575216 -0.802044
+ 1.218e+11Hz 0.574586 -0.802487
+ 1.219e+11Hz 0.573955 -0.802929
+ 1.22e+11Hz 0.573324 -0.803371
+ 1.221e+11Hz 0.572692 -0.803812
+ 1.222e+11Hz 0.57206 -0.804253
+ 1.223e+11Hz 0.571428 -0.804693
+ 1.224e+11Hz 0.570795 -0.805133
+ 1.225e+11Hz 0.570162 -0.805572
+ 1.226e+11Hz 0.569529 -0.806011
+ 1.227e+11Hz 0.568895 -0.806449
+ 1.228e+11Hz 0.568261 -0.806887
+ 1.229e+11Hz 0.567627 -0.807324
+ 1.23e+11Hz 0.566993 -0.807761
+ 1.231e+11Hz 0.566358 -0.808197
+ 1.232e+11Hz 0.565723 -0.808632
+ 1.233e+11Hz 0.565087 -0.809067
+ 1.234e+11Hz 0.564451 -0.809502
+ 1.235e+11Hz 0.563815 -0.809936
+ 1.236e+11Hz 0.563178 -0.810369
+ 1.237e+11Hz 0.562542 -0.810802
+ 1.238e+11Hz 0.561904 -0.811234
+ 1.239e+11Hz 0.561267 -0.811666
+ 1.24e+11Hz 0.560629 -0.812098
+ 1.241e+11Hz 0.559991 -0.812528
+ 1.242e+11Hz 0.559353 -0.812959
+ 1.243e+11Hz 0.558714 -0.813389
+ 1.244e+11Hz 0.558075 -0.813818
+ 1.245e+11Hz 0.557436 -0.814247
+ 1.246e+11Hz 0.556796 -0.814675
+ 1.247e+11Hz 0.556156 -0.815103
+ 1.248e+11Hz 0.555516 -0.81553
+ 1.249e+11Hz 0.554875 -0.815956
+ 1.25e+11Hz 0.554234 -0.816383
+ 1.251e+11Hz 0.553593 -0.816808
+ 1.252e+11Hz 0.552951 -0.817233
+ 1.253e+11Hz 0.552309 -0.817658
+ 1.254e+11Hz 0.551667 -0.818082
+ 1.255e+11Hz 0.551025 -0.818506
+ 1.256e+11Hz 0.550382 -0.818929
+ 1.257e+11Hz 0.549739 -0.819351
+ 1.258e+11Hz 0.549096 -0.819773
+ 1.259e+11Hz 0.548452 -0.820195
+ 1.26e+11Hz 0.547808 -0.820616
+ 1.261e+11Hz 0.547164 -0.821037
+ 1.262e+11Hz 0.546519 -0.821457
+ 1.263e+11Hz 0.545874 -0.821876
+ 1.264e+11Hz 0.545229 -0.822295
+ 1.265e+11Hz 0.544583 -0.822714
+ 1.266e+11Hz 0.543937 -0.823132
+ 1.267e+11Hz 0.543291 -0.823549
+ 1.268e+11Hz 0.542645 -0.823966
+ 1.269e+11Hz 0.541998 -0.824383
+ 1.27e+11Hz 0.541351 -0.824799
+ 1.271e+11Hz 0.540704 -0.825214
+ 1.272e+11Hz 0.540056 -0.825629
+ 1.273e+11Hz 0.539408 -0.826044
+ 1.274e+11Hz 0.53876 -0.826457
+ 1.275e+11Hz 0.538111 -0.826871
+ 1.276e+11Hz 0.537462 -0.827284
+ 1.277e+11Hz 0.536813 -0.827696
+ 1.278e+11Hz 0.536164 -0.828108
+ 1.279e+11Hz 0.535514 -0.82852
+ 1.28e+11Hz 0.534864 -0.828931
+ 1.281e+11Hz 0.534213 -0.829341
+ 1.282e+11Hz 0.533562 -0.829751
+ 1.283e+11Hz 0.532911 -0.830161
+ 1.284e+11Hz 0.53226 -0.83057
+ 1.285e+11Hz 0.531608 -0.830978
+ 1.286e+11Hz 0.530956 -0.831386
+ 1.287e+11Hz 0.530304 -0.831794
+ 1.288e+11Hz 0.529652 -0.832201
+ 1.289e+11Hz 0.528999 -0.832607
+ 1.29e+11Hz 0.528346 -0.833013
+ 1.291e+11Hz 0.527692 -0.833419
+ 1.292e+11Hz 0.527038 -0.833824
+ 1.293e+11Hz 0.526384 -0.834228
+ 1.294e+11Hz 0.52573 -0.834632
+ 1.295e+11Hz 0.525075 -0.835036
+ 1.296e+11Hz 0.52442 -0.835439
+ 1.297e+11Hz 0.523764 -0.835841
+ 1.298e+11Hz 0.523109 -0.836244
+ 1.299e+11Hz 0.522453 -0.836645
+ 1.3e+11Hz 0.521796 -0.837046
+ 1.301e+11Hz 0.52114 -0.837447
+ 1.302e+11Hz 0.520483 -0.837847
+ 1.303e+11Hz 0.519826 -0.838246
+ 1.304e+11Hz 0.519168 -0.838645
+ 1.305e+11Hz 0.51851 -0.839044
+ 1.306e+11Hz 0.517852 -0.839442
+ 1.307e+11Hz 0.517193 -0.83984
+ 1.308e+11Hz 0.516535 -0.840237
+ 1.309e+11Hz 0.515875 -0.840634
+ 1.31e+11Hz 0.515216 -0.84103
+ 1.311e+11Hz 0.514556 -0.841425
+ 1.312e+11Hz 0.513896 -0.84182
+ 1.313e+11Hz 0.513236 -0.842215
+ 1.314e+11Hz 0.512575 -0.842609
+ 1.315e+11Hz 0.511914 -0.843003
+ 1.316e+11Hz 0.511252 -0.843396
+ 1.317e+11Hz 0.510591 -0.843789
+ 1.318e+11Hz 0.509928 -0.844181
+ 1.319e+11Hz 0.509266 -0.844572
+ 1.32e+11Hz 0.508603 -0.844964
+ 1.321e+11Hz 0.50794 -0.845354
+ 1.322e+11Hz 0.507277 -0.845744
+ 1.323e+11Hz 0.506613 -0.846134
+ 1.324e+11Hz 0.505949 -0.846523
+ 1.325e+11Hz 0.505285 -0.846912
+ 1.326e+11Hz 0.50462 -0.8473
+ 1.327e+11Hz 0.503955 -0.847688
+ 1.328e+11Hz 0.50329 -0.848075
+ 1.329e+11Hz 0.502624 -0.848461
+ 1.33e+11Hz 0.501958 -0.848847
+ 1.331e+11Hz 0.501292 -0.849233
+ 1.332e+11Hz 0.500625 -0.849618
+ 1.333e+11Hz 0.499958 -0.850003
+ 1.334e+11Hz 0.499291 -0.850387
+ 1.335e+11Hz 0.498623 -0.85077
+ 1.336e+11Hz 0.497955 -0.851154
+ 1.337e+11Hz 0.497287 -0.851536
+ 1.338e+11Hz 0.496618 -0.851918
+ 1.339e+11Hz 0.495949 -0.8523
+ 1.34e+11Hz 0.49528 -0.852681
+ 1.341e+11Hz 0.49461 -0.853061
+ 1.342e+11Hz 0.49394 -0.853441
+ 1.343e+11Hz 0.49327 -0.853821
+ 1.344e+11Hz 0.492599 -0.8542
+ 1.345e+11Hz 0.491928 -0.854578
+ 1.346e+11Hz 0.491257 -0.854956
+ 1.347e+11Hz 0.490585 -0.855333
+ 1.348e+11Hz 0.489913 -0.85571
+ 1.349e+11Hz 0.489241 -0.856087
+ 1.35e+11Hz 0.488568 -0.856462
+ 1.351e+11Hz 0.487895 -0.856838
+ 1.352e+11Hz 0.487222 -0.857212
+ 1.353e+11Hz 0.486548 -0.857587
+ 1.354e+11Hz 0.485874 -0.85796
+ 1.355e+11Hz 0.4852 -0.858334
+ 1.356e+11Hz 0.484525 -0.858706
+ 1.357e+11Hz 0.48385 -0.859078
+ 1.358e+11Hz 0.483175 -0.85945
+ 1.359e+11Hz 0.482499 -0.859821
+ 1.36e+11Hz 0.481823 -0.860191
+ 1.361e+11Hz 0.481147 -0.860561
+ 1.362e+11Hz 0.48047 -0.860931
+ 1.363e+11Hz 0.479793 -0.8613
+ 1.364e+11Hz 0.479116 -0.861668
+ 1.365e+11Hz 0.478438 -0.862036
+ 1.366e+11Hz 0.47776 -0.862403
+ 1.367e+11Hz 0.477082 -0.86277
+ 1.368e+11Hz 0.476403 -0.863136
+ 1.369e+11Hz 0.475724 -0.863501
+ 1.37e+11Hz 0.475044 -0.863866
+ 1.371e+11Hz 0.474365 -0.864231
+ 1.372e+11Hz 0.473685 -0.864595
+ 1.373e+11Hz 0.473004 -0.864958
+ 1.374e+11Hz 0.472323 -0.865321
+ 1.375e+11Hz 0.471642 -0.865683
+ 1.376e+11Hz 0.470961 -0.866045
+ 1.377e+11Hz 0.470279 -0.866406
+ 1.378e+11Hz 0.469597 -0.866767
+ 1.379e+11Hz 0.468915 -0.867127
+ 1.38e+11Hz 0.468232 -0.867486
+ 1.381e+11Hz 0.467549 -0.867845
+ 1.382e+11Hz 0.466866 -0.868203
+ 1.383e+11Hz 0.466182 -0.868561
+ 1.384e+11Hz 0.465498 -0.868918
+ 1.385e+11Hz 0.464814 -0.869275
+ 1.386e+11Hz 0.464129 -0.869631
+ 1.387e+11Hz 0.463444 -0.869986
+ 1.388e+11Hz 0.462759 -0.870341
+ 1.389e+11Hz 0.462073 -0.870696
+ 1.39e+11Hz 0.461387 -0.871049
+ 1.391e+11Hz 0.460701 -0.871403
+ 1.392e+11Hz 0.460014 -0.871755
+ 1.393e+11Hz 0.459328 -0.872107
+ 1.394e+11Hz 0.45864 -0.872459
+ 1.395e+11Hz 0.457953 -0.872809
+ 1.396e+11Hz 0.457265 -0.87316
+ 1.397e+11Hz 0.456577 -0.873509
+ 1.398e+11Hz 0.455888 -0.873858
+ 1.399e+11Hz 0.4552 -0.874207
+ 1.4e+11Hz 0.45451 -0.874555
+ 1.401e+11Hz 0.453821 -0.874902
+ 1.402e+11Hz 0.453131 -0.875249
+ 1.403e+11Hz 0.452441 -0.875595
+ 1.404e+11Hz 0.451751 -0.87594
+ 1.405e+11Hz 0.45106 -0.876285
+ 1.406e+11Hz 0.450369 -0.87663
+ 1.407e+11Hz 0.449678 -0.876974
+ 1.408e+11Hz 0.448987 -0.877317
+ 1.409e+11Hz 0.448295 -0.877659
+ 1.41e+11Hz 0.447603 -0.878001
+ 1.411e+11Hz 0.44691 -0.878343
+ 1.412e+11Hz 0.446218 -0.878683
+ 1.413e+11Hz 0.445524 -0.879023
+ 1.414e+11Hz 0.444831 -0.879363
+ 1.415e+11Hz 0.444138 -0.879702
+ 1.416e+11Hz 0.443444 -0.88004
+ 1.417e+11Hz 0.44275 -0.880378
+ 1.418e+11Hz 0.442055 -0.880715
+ 1.419e+11Hz 0.44136 -0.881052
+ 1.42e+11Hz 0.440665 -0.881388
+ 1.421e+11Hz 0.43997 -0.881723
+ 1.422e+11Hz 0.439274 -0.882058
+ 1.423e+11Hz 0.438578 -0.882392
+ 1.424e+11Hz 0.437882 -0.882725
+ 1.425e+11Hz 0.437186 -0.883058
+ 1.426e+11Hz 0.436489 -0.883391
+ 1.427e+11Hz 0.435792 -0.883722
+ 1.428e+11Hz 0.435095 -0.884053
+ 1.429e+11Hz 0.434397 -0.884384
+ 1.43e+11Hz 0.433699 -0.884714
+ 1.431e+11Hz 0.433001 -0.885043
+ 1.432e+11Hz 0.432303 -0.885371
+ 1.433e+11Hz 0.431604 -0.885699
+ 1.434e+11Hz 0.430906 -0.886027
+ 1.435e+11Hz 0.430206 -0.886354
+ 1.436e+11Hz 0.429507 -0.88668
+ 1.437e+11Hz 0.428807 -0.887005
+ 1.438e+11Hz 0.428107 -0.88733
+ 1.439e+11Hz 0.427407 -0.887655
+ 1.44e+11Hz 0.426707 -0.887978
+ 1.441e+11Hz 0.426006 -0.888301
+ 1.442e+11Hz 0.425305 -0.888624
+ 1.443e+11Hz 0.424604 -0.888946
+ 1.444e+11Hz 0.423903 -0.889267
+ 1.445e+11Hz 0.423201 -0.889588
+ 1.446e+11Hz 0.422499 -0.889908
+ 1.447e+11Hz 0.421797 -0.890227
+ 1.448e+11Hz 0.421094 -0.890546
+ 1.449e+11Hz 0.420392 -0.890864
+ 1.45e+11Hz 0.419689 -0.891182
+ 1.451e+11Hz 0.418986 -0.891499
+ 1.452e+11Hz 0.418282 -0.891815
+ 1.453e+11Hz 0.417579 -0.892131
+ 1.454e+11Hz 0.416875 -0.892446
+ 1.455e+11Hz 0.416171 -0.89276
+ 1.456e+11Hz 0.415466 -0.893074
+ 1.457e+11Hz 0.414762 -0.893387
+ 1.458e+11Hz 0.414057 -0.8937
+ 1.459e+11Hz 0.413352 -0.894012
+ 1.46e+11Hz 0.412647 -0.894323
+ 1.461e+11Hz 0.411941 -0.894634
+ 1.462e+11Hz 0.411235 -0.894944
+ 1.463e+11Hz 0.410529 -0.895254
+ 1.464e+11Hz 0.409823 -0.895563
+ 1.465e+11Hz 0.409117 -0.895871
+ 1.466e+11Hz 0.40841 -0.896179
+ 1.467e+11Hz 0.407703 -0.896486
+ 1.468e+11Hz 0.406996 -0.896793
+ 1.469e+11Hz 0.406289 -0.897099
+ 1.47e+11Hz 0.405581 -0.897404
+ 1.471e+11Hz 0.404874 -0.897709
+ 1.472e+11Hz 0.404166 -0.898013
+ 1.473e+11Hz 0.403458 -0.898316
+ 1.474e+11Hz 0.402749 -0.898619
+ 1.475e+11Hz 0.402041 -0.898922
+ 1.476e+11Hz 0.401332 -0.899223
+ 1.477e+11Hz 0.400623 -0.899524
+ 1.478e+11Hz 0.399914 -0.899825
+ 1.479e+11Hz 0.399204 -0.900125
+ 1.48e+11Hz 0.398494 -0.900424
+ 1.481e+11Hz 0.397785 -0.900723
+ 1.482e+11Hz 0.397074 -0.901021
+ 1.483e+11Hz 0.396364 -0.901318
+ 1.484e+11Hz 0.395654 -0.901615
+ 1.485e+11Hz 0.394943 -0.901911
+ 1.486e+11Hz 0.394232 -0.902207
+ 1.487e+11Hz 0.393521 -0.902502
+ 1.488e+11Hz 0.39281 -0.902796
+ 1.489e+11Hz 0.392098 -0.90309
+ 1.49e+11Hz 0.391386 -0.903383
+ 1.491e+11Hz 0.390675 -0.903676
+ 1.492e+11Hz 0.389962 -0.903968
+ 1.493e+11Hz 0.38925 -0.904259
+ 1.494e+11Hz 0.388538 -0.90455
+ 1.495e+11Hz 0.387825 -0.90484
+ 1.496e+11Hz 0.387112 -0.90513
+ 1.497e+11Hz 0.386399 -0.905419
+ 1.498e+11Hz 0.385685 -0.905707
+ 1.499e+11Hz 0.384972 -0.905995
+ 1.5e+11Hz 0.384258 -0.906282
+ 1.501e+11Hz 0.383544 -0.906569
+ 1.502e+11Hz 0.38283 -0.906855
+ 1.503e+11Hz 0.382116 -0.907141
+ 1.504e+11Hz 0.381401 -0.907425
+ 1.505e+11Hz 0.380686 -0.90771
+ 1.506e+11Hz 0.379972 -0.907993
+ 1.507e+11Hz 0.379256 -0.908276
+ 1.508e+11Hz 0.378541 -0.908559
+ 1.509e+11Hz 0.377826 -0.908841
+ 1.51e+11Hz 0.37711 -0.909122
+ 1.511e+11Hz 0.376394 -0.909403
+ 1.512e+11Hz 0.375678 -0.909683
+ 1.513e+11Hz 0.374962 -0.909962
+ 1.514e+11Hz 0.374245 -0.910241
+ 1.515e+11Hz 0.373528 -0.91052
+ 1.516e+11Hz 0.372811 -0.910797
+ 1.517e+11Hz 0.372094 -0.911074
+ 1.518e+11Hz 0.371377 -0.911351
+ 1.519e+11Hz 0.37066 -0.911627
+ 1.52e+11Hz 0.369942 -0.911902
+ 1.521e+11Hz 0.369224 -0.912177
+ 1.522e+11Hz 0.368506 -0.912451
+ 1.523e+11Hz 0.367788 -0.912725
+ 1.524e+11Hz 0.367069 -0.912998
+ 1.525e+11Hz 0.366351 -0.91327
+ 1.526e+11Hz 0.365632 -0.913542
+ 1.527e+11Hz 0.364913 -0.913813
+ 1.528e+11Hz 0.364193 -0.914084
+ 1.529e+11Hz 0.363474 -0.914354
+ 1.53e+11Hz 0.362754 -0.914623
+ 1.531e+11Hz 0.362034 -0.914892
+ 1.532e+11Hz 0.361314 -0.915161
+ 1.533e+11Hz 0.360594 -0.915428
+ 1.534e+11Hz 0.359874 -0.915695
+ 1.535e+11Hz 0.359153 -0.915962
+ 1.536e+11Hz 0.358432 -0.916228
+ 1.537e+11Hz 0.357711 -0.916493
+ 1.538e+11Hz 0.35699 -0.916758
+ 1.539e+11Hz 0.356269 -0.917022
+ 1.54e+11Hz 0.355547 -0.917285
+ 1.541e+11Hz 0.354825 -0.917548
+ 1.542e+11Hz 0.354103 -0.91781
+ 1.543e+11Hz 0.353381 -0.918072
+ 1.544e+11Hz 0.352659 -0.918333
+ 1.545e+11Hz 0.351936 -0.918594
+ 1.546e+11Hz 0.351213 -0.918854
+ 1.547e+11Hz 0.35049 -0.919113
+ 1.548e+11Hz 0.349767 -0.919372
+ 1.549e+11Hz 0.349044 -0.91963
+ 1.55e+11Hz 0.34832 -0.919888
+ 1.551e+11Hz 0.347596 -0.920144
+ 1.552e+11Hz 0.346872 -0.920401
+ 1.553e+11Hz 0.346148 -0.920657
+ 1.554e+11Hz 0.345424 -0.920912
+ 1.555e+11Hz 0.344699 -0.921166
+ 1.556e+11Hz 0.343974 -0.92142
+ 1.557e+11Hz 0.343249 -0.921673
+ 1.558e+11Hz 0.342524 -0.921926
+ 1.559e+11Hz 0.341799 -0.922178
+ 1.56e+11Hz 0.341073 -0.92243
+ 1.561e+11Hz 0.340348 -0.922681
+ 1.562e+11Hz 0.339622 -0.922931
+ 1.563e+11Hz 0.338895 -0.923181
+ 1.564e+11Hz 0.338169 -0.92343
+ 1.565e+11Hz 0.337443 -0.923678
+ 1.566e+11Hz 0.336716 -0.923926
+ 1.567e+11Hz 0.335989 -0.924173
+ 1.568e+11Hz 0.335262 -0.92442
+ 1.569e+11Hz 0.334535 -0.924666
+ 1.57e+11Hz 0.333807 -0.924911
+ 1.571e+11Hz 0.333079 -0.925156
+ 1.572e+11Hz 0.332351 -0.9254
+ 1.573e+11Hz 0.331623 -0.925643
+ 1.574e+11Hz 0.330895 -0.925886
+ 1.575e+11Hz 0.330167 -0.926129
+ 1.576e+11Hz 0.329438 -0.92637
+ 1.577e+11Hz 0.328709 -0.926611
+ 1.578e+11Hz 0.32798 -0.926852
+ 1.579e+11Hz 0.327251 -0.927091
+ 1.58e+11Hz 0.326521 -0.927331
+ 1.581e+11Hz 0.325792 -0.927569
+ 1.582e+11Hz 0.325062 -0.927807
+ 1.583e+11Hz 0.324332 -0.928044
+ 1.584e+11Hz 0.323602 -0.928281
+ 1.585e+11Hz 0.322872 -0.928517
+ 1.586e+11Hz 0.322141 -0.928752
+ 1.587e+11Hz 0.32141 -0.928987
+ 1.588e+11Hz 0.320679 -0.929221
+ 1.589e+11Hz 0.319948 -0.929454
+ 1.59e+11Hz 0.319217 -0.929687
+ 1.591e+11Hz 0.318486 -0.929919
+ 1.592e+11Hz 0.317754 -0.930151
+ 1.593e+11Hz 0.317022 -0.930382
+ 1.594e+11Hz 0.31629 -0.930612
+ 1.595e+11Hz 0.315558 -0.930842
+ 1.596e+11Hz 0.314826 -0.931071
+ 1.597e+11Hz 0.314093 -0.931299
+ 1.598e+11Hz 0.313361 -0.931526
+ 1.599e+11Hz 0.312628 -0.931753
+ 1.6e+11Hz 0.311895 -0.93198
+ 1.601e+11Hz 0.311162 -0.932206
+ 1.602e+11Hz 0.310428 -0.932431
+ 1.603e+11Hz 0.309695 -0.932655
+ 1.604e+11Hz 0.308961 -0.932879
+ 1.605e+11Hz 0.308227 -0.933102
+ 1.606e+11Hz 0.307493 -0.933324
+ 1.607e+11Hz 0.306759 -0.933546
+ 1.608e+11Hz 0.306025 -0.933767
+ 1.609e+11Hz 0.305291 -0.933988
+ 1.61e+11Hz 0.304556 -0.934207
+ 1.611e+11Hz 0.303821 -0.934426
+ 1.612e+11Hz 0.303086 -0.934645
+ 1.613e+11Hz 0.302351 -0.934863
+ 1.614e+11Hz 0.301616 -0.93508
+ 1.615e+11Hz 0.300881 -0.935296
+ 1.616e+11Hz 0.300145 -0.935512
+ 1.617e+11Hz 0.299409 -0.935727
+ 1.618e+11Hz 0.298674 -0.935942
+ 1.619e+11Hz 0.297938 -0.936155
+ 1.62e+11Hz 0.297202 -0.936369
+ 1.621e+11Hz 0.296465 -0.936581
+ 1.622e+11Hz 0.295729 -0.936793
+ 1.623e+11Hz 0.294993 -0.937004
+ 1.624e+11Hz 0.294256 -0.937214
+ 1.625e+11Hz 0.293519 -0.937424
+ 1.626e+11Hz 0.292782 -0.937633
+ 1.627e+11Hz 0.292046 -0.937842
+ 1.628e+11Hz 0.291308 -0.938049
+ 1.629e+11Hz 0.290571 -0.938256
+ 1.63e+11Hz 0.289834 -0.938463
+ 1.631e+11Hz 0.289096 -0.938668
+ 1.632e+11Hz 0.288359 -0.938873
+ 1.633e+11Hz 0.287621 -0.939078
+ 1.634e+11Hz 0.286883 -0.939281
+ 1.635e+11Hz 0.286145 -0.939484
+ 1.636e+11Hz 0.285407 -0.939687
+ 1.637e+11Hz 0.284669 -0.939888
+ 1.638e+11Hz 0.283931 -0.940089
+ 1.639e+11Hz 0.283193 -0.940289
+ 1.64e+11Hz 0.282455 -0.940489
+ 1.641e+11Hz 0.281716 -0.940688
+ 1.642e+11Hz 0.280977 -0.940886
+ 1.643e+11Hz 0.280239 -0.941084
+ 1.644e+11Hz 0.2795 -0.941281
+ 1.645e+11Hz 0.278761 -0.941477
+ 1.646e+11Hz 0.278022 -0.941672
+ 1.647e+11Hz 0.277283 -0.941867
+ 1.648e+11Hz 0.276544 -0.942061
+ 1.649e+11Hz 0.275805 -0.942255
+ 1.65e+11Hz 0.275066 -0.942447
+ 1.651e+11Hz 0.274327 -0.94264
+ 1.652e+11Hz 0.273587 -0.942831
+ 1.653e+11Hz 0.272848 -0.943022
+ 1.654e+11Hz 0.272108 -0.943212
+ 1.655e+11Hz 0.271369 -0.943401
+ 1.656e+11Hz 0.270629 -0.94359
+ 1.657e+11Hz 0.269889 -0.943778
+ 1.658e+11Hz 0.26915 -0.943965
+ 1.659e+11Hz 0.26841 -0.944152
+ 1.66e+11Hz 0.26767 -0.944338
+ 1.661e+11Hz 0.26693 -0.944523
+ 1.662e+11Hz 0.26619 -0.944708
+ 1.663e+11Hz 0.26545 -0.944892
+ 1.664e+11Hz 0.26471 -0.945075
+ 1.665e+11Hz 0.26397 -0.945258
+ 1.666e+11Hz 0.26323 -0.94544
+ 1.667e+11Hz 0.26249 -0.945621
+ 1.668e+11Hz 0.26175 -0.945802
+ 1.669e+11Hz 0.26101 -0.945982
+ 1.67e+11Hz 0.26027 -0.946161
+ 1.671e+11Hz 0.259529 -0.946339
+ 1.672e+11Hz 0.258789 -0.946517
+ 1.673e+11Hz 0.258049 -0.946695
+ 1.674e+11Hz 0.257309 -0.946871
+ 1.675e+11Hz 0.256568 -0.947047
+ 1.676e+11Hz 0.255828 -0.947223
+ 1.677e+11Hz 0.255088 -0.947397
+ 1.678e+11Hz 0.254348 -0.947571
+ 1.679e+11Hz 0.253607 -0.947744
+ 1.68e+11Hz 0.252867 -0.947917
+ 1.681e+11Hz 0.252127 -0.948089
+ 1.682e+11Hz 0.251386 -0.94826
+ 1.683e+11Hz 0.250646 -0.948431
+ 1.684e+11Hz 0.249906 -0.948601
+ 1.685e+11Hz 0.249165 -0.948771
+ 1.686e+11Hz 0.248425 -0.948939
+ 1.687e+11Hz 0.247685 -0.949108
+ 1.688e+11Hz 0.246944 -0.949275
+ 1.689e+11Hz 0.246204 -0.949442
+ 1.69e+11Hz 0.245464 -0.949608
+ 1.691e+11Hz 0.244724 -0.949774
+ 1.692e+11Hz 0.243983 -0.949939
+ 1.693e+11Hz 0.243243 -0.950103
+ 1.694e+11Hz 0.242503 -0.950266
+ 1.695e+11Hz 0.241763 -0.950429
+ 1.696e+11Hz 0.241023 -0.950592
+ 1.697e+11Hz 0.240283 -0.950754
+ 1.698e+11Hz 0.239543 -0.950915
+ 1.699e+11Hz 0.238803 -0.951075
+ 1.7e+11Hz 0.238063 -0.951235
+ 1.701e+11Hz 0.237323 -0.951394
+ 1.702e+11Hz 0.236583 -0.951553
+ 1.703e+11Hz 0.235843 -0.951711
+ 1.704e+11Hz 0.235103 -0.951869
+ 1.705e+11Hz 0.234363 -0.952025
+ 1.706e+11Hz 0.233623 -0.952182
+ 1.707e+11Hz 0.232884 -0.952337
+ 1.708e+11Hz 0.232144 -0.952492
+ 1.709e+11Hz 0.231404 -0.952647
+ 1.71e+11Hz 0.230665 -0.952801
+ 1.711e+11Hz 0.229925 -0.952954
+ 1.712e+11Hz 0.229185 -0.953106
+ 1.713e+11Hz 0.228446 -0.953258
+ 1.714e+11Hz 0.227706 -0.95341
+ 1.715e+11Hz 0.226967 -0.953561
+ 1.716e+11Hz 0.226228 -0.953711
+ 1.717e+11Hz 0.225488 -0.953861
+ 1.718e+11Hz 0.224749 -0.95401
+ 1.719e+11Hz 0.22401 -0.954158
+ 1.72e+11Hz 0.223271 -0.954306
+ 1.721e+11Hz 0.222532 -0.954453
+ 1.722e+11Hz 0.221793 -0.9546
+ 1.723e+11Hz 0.221054 -0.954747
+ 1.724e+11Hz 0.220315 -0.954892
+ 1.725e+11Hz 0.219576 -0.955037
+ 1.726e+11Hz 0.218837 -0.955182
+ 1.727e+11Hz 0.218098 -0.955326
+ 1.728e+11Hz 0.21736 -0.955469
+ 1.729e+11Hz 0.216621 -0.955612
+ 1.73e+11Hz 0.215882 -0.955754
+ 1.731e+11Hz 0.215144 -0.955896
+ 1.732e+11Hz 0.214405 -0.956037
+ 1.733e+11Hz 0.213667 -0.956178
+ 1.734e+11Hz 0.212929 -0.956318
+ 1.735e+11Hz 0.21219 -0.956458
+ 1.736e+11Hz 0.211452 -0.956597
+ 1.737e+11Hz 0.210714 -0.956735
+ 1.738e+11Hz 0.209976 -0.956873
+ 1.739e+11Hz 0.209237 -0.95701
+ 1.74e+11Hz 0.208499 -0.957147
+ 1.741e+11Hz 0.207761 -0.957284
+ 1.742e+11Hz 0.207023 -0.957419
+ 1.743e+11Hz 0.206286 -0.957555
+ 1.744e+11Hz 0.205548 -0.957689
+ 1.745e+11Hz 0.20481 -0.957824
+ 1.746e+11Hz 0.204072 -0.957957
+ 1.747e+11Hz 0.203335 -0.958091
+ 1.748e+11Hz 0.202597 -0.958223
+ 1.749e+11Hz 0.201859 -0.958356
+ 1.75e+11Hz 0.201122 -0.958487
+ 1.751e+11Hz 0.200384 -0.958618
+ 1.752e+11Hz 0.199647 -0.958749
+ 1.753e+11Hz 0.19891 -0.958879
+ 1.754e+11Hz 0.198172 -0.959009
+ 1.755e+11Hz 0.197435 -0.959138
+ 1.756e+11Hz 0.196698 -0.959267
+ 1.757e+11Hz 0.195961 -0.959395
+ 1.758e+11Hz 0.195223 -0.959523
+ 1.759e+11Hz 0.194486 -0.95965
+ 1.76e+11Hz 0.193749 -0.959776
+ 1.761e+11Hz 0.193012 -0.959903
+ 1.762e+11Hz 0.192275 -0.960028
+ 1.763e+11Hz 0.191538 -0.960154
+ 1.764e+11Hz 0.190801 -0.960278
+ 1.765e+11Hz 0.190064 -0.960402
+ 1.766e+11Hz 0.189328 -0.960526
+ 1.767e+11Hz 0.188591 -0.96065
+ 1.768e+11Hz 0.187854 -0.960772
+ 1.769e+11Hz 0.187117 -0.960895
+ 1.77e+11Hz 0.186381 -0.961017
+ 1.771e+11Hz 0.185644 -0.961138
+ 1.772e+11Hz 0.184907 -0.961259
+ 1.773e+11Hz 0.184171 -0.961379
+ 1.774e+11Hz 0.183434 -0.961499
+ 1.775e+11Hz 0.182697 -0.961619
+ 1.776e+11Hz 0.181961 -0.961738
+ 1.777e+11Hz 0.181224 -0.961856
+ 1.778e+11Hz 0.180488 -0.961974
+ 1.779e+11Hz 0.179751 -0.962092
+ 1.78e+11Hz 0.179015 -0.962209
+ 1.781e+11Hz 0.178278 -0.962326
+ 1.782e+11Hz 0.177542 -0.962442
+ 1.783e+11Hz 0.176805 -0.962558
+ 1.784e+11Hz 0.176069 -0.962673
+ 1.785e+11Hz 0.175333 -0.962788
+ 1.786e+11Hz 0.174596 -0.962902
+ 1.787e+11Hz 0.17386 -0.963016
+ 1.788e+11Hz 0.173123 -0.96313
+ 1.789e+11Hz 0.172387 -0.963243
+ 1.79e+11Hz 0.171651 -0.963355
+ 1.791e+11Hz 0.170914 -0.963468
+ 1.792e+11Hz 0.170178 -0.963579
+ 1.793e+11Hz 0.169441 -0.96369
+ 1.794e+11Hz 0.168705 -0.963801
+ 1.795e+11Hz 0.167968 -0.963911
+ 1.796e+11Hz 0.167232 -0.964021
+ 1.797e+11Hz 0.166496 -0.964131
+ 1.798e+11Hz 0.165759 -0.96424
+ 1.799e+11Hz 0.165023 -0.964348
+ 1.8e+11Hz 0.164286 -0.964456
+ 1.801e+11Hz 0.16355 -0.964564
+ 1.802e+11Hz 0.162813 -0.964671
+ 1.803e+11Hz 0.162077 -0.964778
+ 1.804e+11Hz 0.16134 -0.964884
+ 1.805e+11Hz 0.160604 -0.96499
+ 1.806e+11Hz 0.159867 -0.965095
+ 1.807e+11Hz 0.15913 -0.9652
+ 1.808e+11Hz 0.158394 -0.965304
+ 1.809e+11Hz 0.157657 -0.965408
+ 1.81e+11Hz 0.15692 -0.965512
+ 1.811e+11Hz 0.156184 -0.965615
+ 1.812e+11Hz 0.155447 -0.965718
+ 1.813e+11Hz 0.15471 -0.96582
+ 1.814e+11Hz 0.153973 -0.965921
+ 1.815e+11Hz 0.153236 -0.966023
+ 1.816e+11Hz 0.152499 -0.966124
+ 1.817e+11Hz 0.151762 -0.966224
+ 1.818e+11Hz 0.151025 -0.966324
+ 1.819e+11Hz 0.150288 -0.966423
+ 1.82e+11Hz 0.149551 -0.966522
+ 1.821e+11Hz 0.148814 -0.966621
+ 1.822e+11Hz 0.148077 -0.966719
+ 1.823e+11Hz 0.14734 -0.966817
+ 1.824e+11Hz 0.146602 -0.966914
+ 1.825e+11Hz 0.145865 -0.967011
+ 1.826e+11Hz 0.145128 -0.967107
+ 1.827e+11Hz 0.14439 -0.967203
+ 1.828e+11Hz 0.143653 -0.967298
+ 1.829e+11Hz 0.142915 -0.967393
+ 1.83e+11Hz 0.142178 -0.967488
+ 1.831e+11Hz 0.14144 -0.967582
+ 1.832e+11Hz 0.140702 -0.967675
+ 1.833e+11Hz 0.139965 -0.967768
+ 1.834e+11Hz 0.139227 -0.967861
+ 1.835e+11Hz 0.138489 -0.967953
+ 1.836e+11Hz 0.137751 -0.968045
+ 1.837e+11Hz 0.137013 -0.968136
+ 1.838e+11Hz 0.136275 -0.968227
+ 1.839e+11Hz 0.135537 -0.968317
+ 1.84e+11Hz 0.134799 -0.968407
+ 1.841e+11Hz 0.13406 -0.968496
+ 1.842e+11Hz 0.133322 -0.968585
+ 1.843e+11Hz 0.132584 -0.968673
+ 1.844e+11Hz 0.131845 -0.968761
+ 1.845e+11Hz 0.131107 -0.968849
+ 1.846e+11Hz 0.130368 -0.968936
+ 1.847e+11Hz 0.129629 -0.969022
+ 1.848e+11Hz 0.128891 -0.969109
+ 1.849e+11Hz 0.128152 -0.969194
+ 1.85e+11Hz 0.127413 -0.969279
+ 1.851e+11Hz 0.126674 -0.969364
+ 1.852e+11Hz 0.125935 -0.969448
+ 1.853e+11Hz 0.125196 -0.969532
+ 1.854e+11Hz 0.124457 -0.969615
+ 1.855e+11Hz 0.123717 -0.969698
+ 1.856e+11Hz 0.122978 -0.96978
+ 1.857e+11Hz 0.122239 -0.969862
+ 1.858e+11Hz 0.121499 -0.969943
+ 1.859e+11Hz 0.120759 -0.970024
+ 1.86e+11Hz 0.12002 -0.970104
+ 1.861e+11Hz 0.11928 -0.970184
+ 1.862e+11Hz 0.11854 -0.970263
+ 1.863e+11Hz 0.1178 -0.970342
+ 1.864e+11Hz 0.11706 -0.97042
+ 1.865e+11Hz 0.11632 -0.970498
+ 1.866e+11Hz 0.11558 -0.970576
+ 1.867e+11Hz 0.11484 -0.970652
+ 1.868e+11Hz 0.1141 -0.970729
+ 1.869e+11Hz 0.113359 -0.970805
+ 1.87e+11Hz 0.112619 -0.97088
+ 1.871e+11Hz 0.111878 -0.970955
+ 1.872e+11Hz 0.111138 -0.971029
+ 1.873e+11Hz 0.110397 -0.971103
+ 1.874e+11Hz 0.109656 -0.971177
+ 1.875e+11Hz 0.108915 -0.971249
+ 1.876e+11Hz 0.108175 -0.971322
+ 1.877e+11Hz 0.107434 -0.971394
+ 1.878e+11Hz 0.106692 -0.971465
+ 1.879e+11Hz 0.105951 -0.971536
+ 1.88e+11Hz 0.10521 -0.971606
+ 1.881e+11Hz 0.104469 -0.971676
+ 1.882e+11Hz 0.103727 -0.971745
+ 1.883e+11Hz 0.102986 -0.971814
+ 1.884e+11Hz 0.102244 -0.971883
+ 1.885e+11Hz 0.101503 -0.97195
+ 1.886e+11Hz 0.100761 -0.972018
+ 1.887e+11Hz 0.100019 -0.972084
+ 1.888e+11Hz 0.0992772 -0.972151
+ 1.889e+11Hz 0.0985352 -0.972216
+ 1.89e+11Hz 0.0977932 -0.972282
+ 1.891e+11Hz 0.0970511 -0.972346
+ 1.892e+11Hz 0.0963089 -0.972411
+ 1.893e+11Hz 0.0955666 -0.972474
+ 1.894e+11Hz 0.0948242 -0.972537
+ 1.895e+11Hz 0.0940818 -0.9726
+ 1.896e+11Hz 0.0933393 -0.972662
+ 1.897e+11Hz 0.0925967 -0.972724
+ 1.898e+11Hz 0.0918541 -0.972785
+ 1.899e+11Hz 0.0911114 -0.972845
+ 1.9e+11Hz 0.0903686 -0.972905
+ 1.901e+11Hz 0.0896257 -0.972965
+ 1.902e+11Hz 0.0888827 -0.973024
+ 1.903e+11Hz 0.0881397 -0.973082
+ 1.904e+11Hz 0.0873966 -0.97314
+ 1.905e+11Hz 0.0866534 -0.973198
+ 1.906e+11Hz 0.0859102 -0.973254
+ 1.907e+11Hz 0.0851669 -0.973311
+ 1.908e+11Hz 0.0844235 -0.973367
+ 1.909e+11Hz 0.08368 -0.973422
+ 1.91e+11Hz 0.0829365 -0.973477
+ 1.911e+11Hz 0.0821929 -0.973531
+ 1.912e+11Hz 0.0814492 -0.973584
+ 1.913e+11Hz 0.0807055 -0.973638
+ 1.914e+11Hz 0.0799617 -0.97369
+ 1.915e+11Hz 0.0792178 -0.973742
+ 1.916e+11Hz 0.0784739 -0.973794
+ 1.917e+11Hz 0.0777299 -0.973845
+ 1.918e+11Hz 0.0769858 -0.973895
+ 1.919e+11Hz 0.0762416 -0.973945
+ 1.92e+11Hz 0.0754974 -0.973995
+ 1.921e+11Hz 0.0747532 -0.974043
+ 1.922e+11Hz 0.0740088 -0.974092
+ 1.923e+11Hz 0.0732644 -0.97414
+ 1.924e+11Hz 0.0725199 -0.974187
+ 1.925e+11Hz 0.0717754 -0.974233
+ 1.926e+11Hz 0.0710308 -0.97428
+ 1.927e+11Hz 0.0702861 -0.974325
+ 1.928e+11Hz 0.0695414 -0.97437
+ 1.929e+11Hz 0.0687966 -0.974415
+ 1.93e+11Hz 0.0680518 -0.974459
+ 1.931e+11Hz 0.0673068 -0.974502
+ 1.932e+11Hz 0.0665619 -0.974545
+ 1.933e+11Hz 0.0658168 -0.974588
+ 1.934e+11Hz 0.0650717 -0.974629
+ 1.935e+11Hz 0.0643266 -0.974671
+ 1.936e+11Hz 0.0635814 -0.974711
+ 1.937e+11Hz 0.0628361 -0.974752
+ 1.938e+11Hz 0.0620907 -0.974791
+ 1.939e+11Hz 0.0613453 -0.97483
+ 1.94e+11Hz 0.0605999 -0.974869
+ 1.941e+11Hz 0.0598544 -0.974907
+ 1.942e+11Hz 0.0591088 -0.974944
+ 1.943e+11Hz 0.0583632 -0.974981
+ 1.944e+11Hz 0.0576175 -0.975018
+ 1.945e+11Hz 0.0568717 -0.975054
+ 1.946e+11Hz 0.0561259 -0.975089
+ 1.947e+11Hz 0.0553801 -0.975123
+ 1.948e+11Hz 0.0546342 -0.975158
+ 1.949e+11Hz 0.0538882 -0.975191
+ 1.95e+11Hz 0.0531422 -0.975224
+ 1.951e+11Hz 0.0523961 -0.975257
+ 1.952e+11Hz 0.05165 -0.975289
+ 1.953e+11Hz 0.0509038 -0.97532
+ 1.954e+11Hz 0.0501575 -0.975351
+ 1.955e+11Hz 0.0494112 -0.975381
+ 1.956e+11Hz 0.0486649 -0.975411
+ 1.957e+11Hz 0.0479185 -0.97544
+ 1.958e+11Hz 0.047172 -0.975469
+ 1.959e+11Hz 0.0464255 -0.975497
+ 1.96e+11Hz 0.045679 -0.975525
+ 1.961e+11Hz 0.0449323 -0.975552
+ 1.962e+11Hz 0.0441857 -0.975578
+ 1.963e+11Hz 0.043439 -0.975604
+ 1.964e+11Hz 0.0426922 -0.975629
+ 1.965e+11Hz 0.0419454 -0.975654
+ 1.966e+11Hz 0.0411985 -0.975678
+ 1.967e+11Hz 0.0404515 -0.975702
+ 1.968e+11Hz 0.0397046 -0.975725
+ 1.969e+11Hz 0.0389575 -0.975748
+ 1.97e+11Hz 0.0382104 -0.97577
+ 1.971e+11Hz 0.0374633 -0.975791
+ 1.972e+11Hz 0.0367161 -0.975812
+ 1.973e+11Hz 0.0359689 -0.975832
+ 1.974e+11Hz 0.0352216 -0.975852
+ 1.975e+11Hz 0.0344743 -0.975871
+ 1.976e+11Hz 0.0337269 -0.97589
+ 1.977e+11Hz 0.0329794 -0.975908
+ 1.978e+11Hz 0.032232 -0.975925
+ 1.979e+11Hz 0.0314844 -0.975942
+ 1.98e+11Hz 0.0307368 -0.975958
+ 1.981e+11Hz 0.0299892 -0.975974
+ 1.982e+11Hz 0.0292415 -0.975989
+ 1.983e+11Hz 0.0284938 -0.976004
+ 1.984e+11Hz 0.027746 -0.976018
+ 1.985e+11Hz 0.0269982 -0.976031
+ 1.986e+11Hz 0.0262503 -0.976044
+ 1.987e+11Hz 0.0255024 -0.976057
+ 1.988e+11Hz 0.0247544 -0.976068
+ 1.989e+11Hz 0.0240064 -0.97608
+ 1.99e+11Hz 0.0232584 -0.97609
+ 1.991e+11Hz 0.0225103 -0.9761
+ 1.992e+11Hz 0.0217621 -0.97611
+ 1.993e+11Hz 0.0210139 -0.976119
+ 1.994e+11Hz 0.0202657 -0.976127
+ 1.995e+11Hz 0.0195174 -0.976135
+ 1.996e+11Hz 0.018769 -0.976142
+ 1.997e+11Hz 0.0180206 -0.976148
+ 1.998e+11Hz 0.0172722 -0.976154
+ 1.999e+11Hz 0.0165238 -0.97616
+ 2e+11Hz 0.0157752 -0.976165
+ 2.001e+11Hz 0.0150267 -0.976169
+ 2.002e+11Hz 0.0142781 -0.976173
+ 2.003e+11Hz 0.0135295 -0.976176
+ 2.004e+11Hz 0.0127808 -0.976178
+ 2.005e+11Hz 0.0120321 -0.97618
+ 2.006e+11Hz 0.0112833 -0.976181
+ 2.007e+11Hz 0.0105345 -0.976182
+ 2.008e+11Hz 0.00978566 -0.976182
+ 2.009e+11Hz 0.00903679 -0.976182
+ 2.01e+11Hz 0.00828787 -0.976181
+ 2.011e+11Hz 0.00753892 -0.976179
+ 2.012e+11Hz 0.00678993 -0.976177
+ 2.013e+11Hz 0.00604091 -0.976174
+ 2.014e+11Hz 0.00529185 -0.97617
+ 2.015e+11Hz 0.00454275 -0.976166
+ 2.016e+11Hz 0.00379363 -0.976162
+ 2.017e+11Hz 0.00304447 -0.976156
+ 2.018e+11Hz 0.00229528 -0.97615
+ 2.019e+11Hz 0.00154605 -0.976144
+ 2.02e+11Hz 0.000796802 -0.976137
+ 2.021e+11Hz 4.7521e-05 -0.976129
+ 2.022e+11Hz -0.000701788 -0.976121
+ 2.023e+11Hz -0.00145112 -0.976112
+ 2.024e+11Hz -0.00220049 -0.976102
+ 2.025e+11Hz -0.00294987 -0.976092
+ 2.026e+11Hz -0.00369929 -0.976081
+ 2.027e+11Hz -0.00444872 -0.97607
+ 2.028e+11Hz -0.00519818 -0.976058
+ 2.029e+11Hz -0.00594765 -0.976045
+ 2.03e+11Hz -0.00669715 -0.976032
+ 2.031e+11Hz -0.00744666 -0.976018
+ 2.032e+11Hz -0.00819619 -0.976004
+ 2.033e+11Hz -0.00894573 -0.975988
+ 2.034e+11Hz -0.00969529 -0.975973
+ 2.035e+11Hz -0.0104449 -0.975956
+ 2.036e+11Hz -0.0111944 -0.975939
+ 2.037e+11Hz -0.011944 -0.975922
+ 2.038e+11Hz -0.0126936 -0.975903
+ 2.039e+11Hz -0.0134432 -0.975884
+ 2.04e+11Hz -0.0141928 -0.975865
+ 2.041e+11Hz -0.0149425 -0.975845
+ 2.042e+11Hz -0.0156921 -0.975824
+ 2.043e+11Hz -0.0164417 -0.975802
+ 2.044e+11Hz -0.0171913 -0.97578
+ 2.045e+11Hz -0.0179409 -0.975758
+ 2.046e+11Hz -0.0186905 -0.975734
+ 2.047e+11Hz -0.0194401 -0.97571
+ 2.048e+11Hz -0.0201897 -0.975686
+ 2.049e+11Hz -0.0209393 -0.97566
+ 2.05e+11Hz -0.0216888 -0.975634
+ 2.051e+11Hz -0.0224384 -0.975608
+ 2.052e+11Hz -0.0231879 -0.975581
+ 2.053e+11Hz -0.0239374 -0.975553
+ 2.054e+11Hz -0.0246869 -0.975524
+ 2.055e+11Hz -0.0254363 -0.975495
+ 2.056e+11Hz -0.0261858 -0.975465
+ 2.057e+11Hz -0.0269352 -0.975435
+ 2.058e+11Hz -0.0276845 -0.975403
+ 2.059e+11Hz -0.0284339 -0.975372
+ 2.06e+11Hz -0.0291832 -0.975339
+ 2.061e+11Hz -0.0299325 -0.975306
+ 2.062e+11Hz -0.0306817 -0.975272
+ 2.063e+11Hz -0.0314309 -0.975238
+ 2.064e+11Hz -0.03218 -0.975203
+ 2.065e+11Hz -0.0329291 -0.975167
+ 2.066e+11Hz -0.0336781 -0.975131
+ 2.067e+11Hz -0.0344271 -0.975094
+ 2.068e+11Hz -0.035176 -0.975056
+ 2.069e+11Hz -0.0359249 -0.975017
+ 2.07e+11Hz -0.0366737 -0.974978
+ 2.071e+11Hz -0.0374225 -0.974939
+ 2.072e+11Hz -0.0381711 -0.974898
+ 2.073e+11Hz -0.0389197 -0.974857
+ 2.074e+11Hz -0.0396683 -0.974816
+ 2.075e+11Hz -0.0404167 -0.974773
+ 2.076e+11Hz -0.0411651 -0.97473
+ 2.077e+11Hz -0.0419134 -0.974686
+ 2.078e+11Hz -0.0426616 -0.974642
+ 2.079e+11Hz -0.0434098 -0.974597
+ 2.08e+11Hz -0.0441578 -0.974551
+ 2.081e+11Hz -0.0449058 -0.974505
+ 2.082e+11Hz -0.0456536 -0.974458
+ 2.083e+11Hz -0.0464014 -0.97441
+ 2.084e+11Hz -0.047149 -0.974362
+ 2.085e+11Hz -0.0478966 -0.974313
+ 2.086e+11Hz -0.048644 -0.974263
+ 2.087e+11Hz -0.0493913 -0.974213
+ 2.088e+11Hz -0.0501385 -0.974162
+ 2.089e+11Hz -0.0508856 -0.974111
+ 2.09e+11Hz -0.0516326 -0.974058
+ 2.091e+11Hz -0.0523794 -0.974005
+ 2.092e+11Hz -0.0531262 -0.973952
+ 2.093e+11Hz -0.0538728 -0.973897
+ 2.094e+11Hz -0.0546192 -0.973843
+ 2.095e+11Hz -0.0553656 -0.973787
+ 2.096e+11Hz -0.0561117 -0.973731
+ 2.097e+11Hz -0.0568578 -0.973674
+ 2.098e+11Hz -0.0576037 -0.973616
+ 2.099e+11Hz -0.0583494 -0.973558
+ 2.1e+11Hz -0.059095 -0.973499
+ 2.101e+11Hz -0.0598405 -0.97344
+ 2.102e+11Hz -0.0605858 -0.97338
+ 2.103e+11Hz -0.0613309 -0.973319
+ 2.104e+11Hz -0.0620758 -0.973257
+ 2.105e+11Hz -0.0628206 -0.973195
+ 2.106e+11Hz -0.0635652 -0.973133
+ 2.107e+11Hz -0.0643097 -0.973069
+ 2.108e+11Hz -0.065054 -0.973005
+ 2.109e+11Hz -0.0657981 -0.972941
+ 2.11e+11Hz -0.066542 -0.972875
+ 2.111e+11Hz -0.0672857 -0.97281
+ 2.112e+11Hz -0.0680292 -0.972743
+ 2.113e+11Hz -0.0687726 -0.972676
+ 2.114e+11Hz -0.0695157 -0.972608
+ 2.115e+11Hz -0.0702587 -0.97254
+ 2.116e+11Hz -0.0710014 -0.972471
+ 2.117e+11Hz -0.071744 -0.972401
+ 2.118e+11Hz -0.0724863 -0.972331
+ 2.119e+11Hz -0.0732284 -0.97226
+ 2.12e+11Hz -0.0739704 -0.972189
+ 2.121e+11Hz -0.0747121 -0.972116
+ 2.122e+11Hz -0.0754535 -0.972044
+ 2.123e+11Hz -0.0761948 -0.97197
+ 2.124e+11Hz -0.0769359 -0.971897
+ 2.125e+11Hz -0.0776767 -0.971822
+ 2.126e+11Hz -0.0784173 -0.971747
+ 2.127e+11Hz -0.0791577 -0.971671
+ 2.128e+11Hz -0.0798978 -0.971595
+ 2.129e+11Hz -0.0806377 -0.971518
+ 2.13e+11Hz -0.0813774 -0.971441
+ 2.131e+11Hz -0.0821168 -0.971363
+ 2.132e+11Hz -0.082856 -0.971284
+ 2.133e+11Hz -0.0835949 -0.971205
+ 2.134e+11Hz -0.0843336 -0.971125
+ 2.135e+11Hz -0.0850721 -0.971045
+ 2.136e+11Hz -0.0858103 -0.970964
+ 2.137e+11Hz -0.0865482 -0.970883
+ 2.138e+11Hz -0.0872859 -0.970801
+ 2.139e+11Hz -0.0880233 -0.970718
+ 2.14e+11Hz -0.0887605 -0.970635
+ 2.141e+11Hz -0.0894975 -0.970552
+ 2.142e+11Hz -0.0902341 -0.970468
+ 2.143e+11Hz -0.0909705 -0.970383
+ 2.144e+11Hz -0.0917067 -0.970298
+ 2.145e+11Hz -0.0924426 -0.970212
+ 2.146e+11Hz -0.0931782 -0.970126
+ 2.147e+11Hz -0.0939135 -0.970039
+ 2.148e+11Hz -0.0946486 -0.969952
+ 2.149e+11Hz -0.0953834 -0.969864
+ 2.15e+11Hz -0.096118 -0.969776
+ 2.151e+11Hz -0.0968523 -0.969687
+ 2.152e+11Hz -0.0975863 -0.969597
+ 2.153e+11Hz -0.09832 -0.969508
+ 2.154e+11Hz -0.0990535 -0.969417
+ 2.155e+11Hz -0.0997867 -0.969327
+ 2.156e+11Hz -0.10052 -0.969235
+ 2.157e+11Hz -0.101252 -0.969144
+ 2.158e+11Hz -0.101985 -0.969051
+ 2.159e+11Hz -0.102717 -0.968959
+ 2.16e+11Hz -0.103449 -0.968866
+ 2.161e+11Hz -0.10418 -0.968772
+ 2.162e+11Hz -0.104911 -0.968678
+ 2.163e+11Hz -0.105642 -0.968583
+ 2.164e+11Hz -0.106373 -0.968488
+ 2.165e+11Hz -0.107104 -0.968393
+ 2.166e+11Hz -0.107834 -0.968297
+ 2.167e+11Hz -0.108564 -0.968201
+ 2.168e+11Hz -0.109293 -0.968104
+ 2.169e+11Hz -0.110023 -0.968007
+ 2.17e+11Hz -0.110752 -0.96791
+ 2.171e+11Hz -0.111481 -0.967812
+ 2.172e+11Hz -0.112209 -0.967713
+ 2.173e+11Hz -0.112937 -0.967615
+ 2.174e+11Hz -0.113666 -0.967515
+ 2.175e+11Hz -0.114393 -0.967416
+ 2.176e+11Hz -0.115121 -0.967316
+ 2.177e+11Hz -0.115848 -0.967216
+ 2.178e+11Hz -0.116575 -0.967115
+ 2.179e+11Hz -0.117302 -0.967014
+ 2.18e+11Hz -0.118028 -0.966912
+ 2.181e+11Hz -0.118754 -0.96681
+ 2.182e+11Hz -0.11948 -0.966708
+ 2.183e+11Hz -0.120206 -0.966606
+ 2.184e+11Hz -0.120932 -0.966503
+ 2.185e+11Hz -0.121657 -0.966399
+ 2.186e+11Hz -0.122382 -0.966296
+ 2.187e+11Hz -0.123106 -0.966192
+ 2.188e+11Hz -0.123831 -0.966087
+ 2.189e+11Hz -0.124555 -0.965983
+ 2.19e+11Hz -0.125279 -0.965878
+ 2.191e+11Hz -0.126003 -0.965772
+ 2.192e+11Hz -0.126727 -0.965667
+ 2.193e+11Hz -0.12745 -0.965561
+ 2.194e+11Hz -0.128173 -0.965454
+ 2.195e+11Hz -0.128896 -0.965348
+ 2.196e+11Hz -0.129619 -0.965241
+ 2.197e+11Hz -0.130341 -0.965134
+ 2.198e+11Hz -0.131063 -0.965026
+ 2.199e+11Hz -0.131786 -0.964918
+ 2.2e+11Hz -0.132507 -0.96481
+ 2.201e+11Hz -0.133229 -0.964702
+ 2.202e+11Hz -0.133951 -0.964593
+ 2.203e+11Hz -0.134672 -0.964484
+ 2.204e+11Hz -0.135393 -0.964375
+ 2.205e+11Hz -0.136114 -0.964265
+ 2.206e+11Hz -0.136835 -0.964155
+ 2.207e+11Hz -0.137555 -0.964045
+ 2.208e+11Hz -0.138275 -0.963935
+ 2.209e+11Hz -0.138996 -0.963824
+ 2.21e+11Hz -0.139716 -0.963713
+ 2.211e+11Hz -0.140436 -0.963602
+ 2.212e+11Hz -0.141155 -0.963491
+ 2.213e+11Hz -0.141875 -0.963379
+ 2.214e+11Hz -0.142594 -0.963267
+ 2.215e+11Hz -0.143314 -0.963155
+ 2.216e+11Hz -0.144033 -0.963042
+ 2.217e+11Hz -0.144752 -0.96293
+ 2.218e+11Hz -0.145471 -0.962817
+ 2.219e+11Hz -0.14619 -0.962703
+ 2.22e+11Hz -0.146908 -0.96259
+ 2.221e+11Hz -0.147627 -0.962476
+ 2.222e+11Hz -0.148346 -0.962362
+ 2.223e+11Hz -0.149064 -0.962248
+ 2.224e+11Hz -0.149782 -0.962134
+ 2.225e+11Hz -0.1505 -0.962019
+ 2.226e+11Hz -0.151219 -0.961904
+ 2.227e+11Hz -0.151937 -0.961789
+ 2.228e+11Hz -0.152655 -0.961673
+ 2.229e+11Hz -0.153372 -0.961558
+ 2.23e+11Hz -0.15409 -0.961442
+ 2.231e+11Hz -0.154808 -0.961326
+ 2.232e+11Hz -0.155526 -0.96121
+ 2.233e+11Hz -0.156243 -0.961093
+ 2.234e+11Hz -0.156961 -0.960976
+ 2.235e+11Hz -0.157679 -0.960859
+ 2.236e+11Hz -0.158396 -0.960742
+ 2.237e+11Hz -0.159114 -0.960625
+ 2.238e+11Hz -0.159831 -0.960507
+ 2.239e+11Hz -0.160549 -0.960389
+ 2.24e+11Hz -0.161266 -0.960271
+ 2.241e+11Hz -0.161984 -0.960152
+ 2.242e+11Hz -0.162701 -0.960034
+ 2.243e+11Hz -0.163419 -0.959915
+ 2.244e+11Hz -0.164136 -0.959796
+ 2.245e+11Hz -0.164854 -0.959677
+ 2.246e+11Hz -0.165571 -0.959557
+ 2.247e+11Hz -0.166289 -0.959437
+ 2.248e+11Hz -0.167006 -0.959317
+ 2.249e+11Hz -0.167724 -0.959197
+ 2.25e+11Hz -0.168442 -0.959076
+ 2.251e+11Hz -0.169159 -0.958955
+ 2.252e+11Hz -0.169877 -0.958834
+ 2.253e+11Hz -0.170595 -0.958713
+ 2.254e+11Hz -0.171313 -0.958592
+ 2.255e+11Hz -0.172031 -0.95847
+ 2.256e+11Hz -0.172749 -0.958348
+ 2.257e+11Hz -0.173467 -0.958225
+ 2.258e+11Hz -0.174185 -0.958103
+ 2.259e+11Hz -0.174904 -0.95798
+ 2.26e+11Hz -0.175622 -0.957857
+ 2.261e+11Hz -0.176341 -0.957734
+ 2.262e+11Hz -0.177059 -0.95761
+ 2.263e+11Hz -0.177778 -0.957486
+ 2.264e+11Hz -0.178497 -0.957362
+ 2.265e+11Hz -0.179216 -0.957238
+ 2.266e+11Hz -0.179935 -0.957113
+ 2.267e+11Hz -0.180654 -0.956988
+ 2.268e+11Hz -0.181374 -0.956862
+ 2.269e+11Hz -0.182093 -0.956737
+ 2.27e+11Hz -0.182813 -0.956611
+ 2.271e+11Hz -0.183533 -0.956485
+ 2.272e+11Hz -0.184252 -0.956358
+ 2.273e+11Hz -0.184973 -0.956231
+ 2.274e+11Hz -0.185693 -0.956104
+ 2.275e+11Hz -0.186413 -0.955977
+ 2.276e+11Hz -0.187134 -0.955849
+ 2.277e+11Hz -0.187855 -0.955721
+ 2.278e+11Hz -0.188576 -0.955592
+ 2.279e+11Hz -0.189297 -0.955464
+ 2.28e+11Hz -0.190018 -0.955335
+ 2.281e+11Hz -0.19074 -0.955205
+ 2.282e+11Hz -0.191461 -0.955075
+ 2.283e+11Hz -0.192183 -0.954945
+ 2.284e+11Hz -0.192905 -0.954815
+ 2.285e+11Hz -0.193627 -0.954684
+ 2.286e+11Hz -0.19435 -0.954552
+ 2.287e+11Hz -0.195073 -0.954421
+ 2.288e+11Hz -0.195796 -0.954289
+ 2.289e+11Hz -0.196519 -0.954156
+ 2.29e+11Hz -0.197242 -0.954023
+ 2.291e+11Hz -0.197965 -0.95389
+ 2.292e+11Hz -0.198689 -0.953757
+ 2.293e+11Hz -0.199413 -0.953623
+ 2.294e+11Hz -0.200137 -0.953488
+ 2.295e+11Hz -0.200862 -0.953353
+ 2.296e+11Hz -0.201587 -0.953218
+ 2.297e+11Hz -0.202311 -0.953082
+ 2.298e+11Hz -0.203037 -0.952946
+ 2.299e+11Hz -0.203762 -0.95281
+ 2.3e+11Hz -0.204487 -0.952673
+ 2.301e+11Hz -0.205213 -0.952535
+ 2.302e+11Hz -0.205939 -0.952397
+ 2.303e+11Hz -0.206666 -0.952259
+ 2.304e+11Hz -0.207392 -0.95212
+ 2.305e+11Hz -0.208119 -0.95198
+ 2.306e+11Hz -0.208846 -0.951841
+ 2.307e+11Hz -0.209573 -0.9517
+ 2.308e+11Hz -0.210301 -0.951559
+ 2.309e+11Hz -0.211029 -0.951418
+ 2.31e+11Hz -0.211757 -0.951276
+ 2.311e+11Hz -0.212485 -0.951134
+ 2.312e+11Hz -0.213213 -0.950991
+ 2.313e+11Hz -0.213942 -0.950848
+ 2.314e+11Hz -0.214671 -0.950704
+ 2.315e+11Hz -0.2154 -0.950559
+ 2.316e+11Hz -0.21613 -0.950414
+ 2.317e+11Hz -0.21686 -0.950268
+ 2.318e+11Hz -0.21759 -0.950122
+ 2.319e+11Hz -0.21832 -0.949976
+ 2.32e+11Hz -0.21905 -0.949828
+ 2.321e+11Hz -0.219781 -0.94968
+ 2.322e+11Hz -0.220512 -0.949532
+ 2.323e+11Hz -0.221243 -0.949383
+ 2.324e+11Hz -0.221974 -0.949233
+ 2.325e+11Hz -0.222706 -0.949083
+ 2.326e+11Hz -0.223438 -0.948932
+ 2.327e+11Hz -0.22417 -0.948781
+ 2.328e+11Hz -0.224902 -0.948629
+ 2.329e+11Hz -0.225635 -0.948476
+ 2.33e+11Hz -0.226368 -0.948323
+ 2.331e+11Hz -0.227101 -0.948169
+ 2.332e+11Hz -0.227834 -0.948014
+ 2.333e+11Hz -0.228568 -0.947859
+ 2.334e+11Hz -0.229301 -0.947703
+ 2.335e+11Hz -0.230035 -0.947546
+ 2.336e+11Hz -0.230769 -0.947389
+ 2.337e+11Hz -0.231504 -0.947231
+ 2.338e+11Hz -0.232238 -0.947073
+ 2.339e+11Hz -0.232973 -0.946913
+ 2.34e+11Hz -0.233708 -0.946753
+ 2.341e+11Hz -0.234443 -0.946593
+ 2.342e+11Hz -0.235178 -0.946431
+ 2.343e+11Hz -0.235914 -0.946269
+ 2.344e+11Hz -0.23665 -0.946107
+ 2.345e+11Hz -0.237385 -0.945943
+ 2.346e+11Hz -0.238122 -0.945779
+ 2.347e+11Hz -0.238858 -0.945614
+ 2.348e+11Hz -0.239594 -0.945448
+ 2.349e+11Hz -0.240331 -0.945282
+ 2.35e+11Hz -0.241068 -0.945115
+ 2.351e+11Hz -0.241805 -0.944947
+ 2.352e+11Hz -0.242542 -0.944778
+ 2.353e+11Hz -0.243279 -0.944609
+ 2.354e+11Hz -0.244016 -0.944439
+ 2.355e+11Hz -0.244754 -0.944268
+ 2.356e+11Hz -0.245491 -0.944096
+ 2.357e+11Hz -0.246229 -0.943924
+ 2.358e+11Hz -0.246967 -0.943751
+ 2.359e+11Hz -0.247705 -0.943577
+ 2.36e+11Hz -0.248443 -0.943402
+ 2.361e+11Hz -0.249182 -0.943227
+ 2.362e+11Hz -0.24992 -0.94305
+ 2.363e+11Hz -0.250659 -0.942873
+ 2.364e+11Hz -0.251397 -0.942695
+ 2.365e+11Hz -0.252136 -0.942517
+ 2.366e+11Hz -0.252875 -0.942337
+ 2.367e+11Hz -0.253614 -0.942157
+ 2.368e+11Hz -0.254353 -0.941976
+ 2.369e+11Hz -0.255092 -0.941794
+ 2.37e+11Hz -0.255831 -0.941611
+ 2.371e+11Hz -0.25657 -0.941427
+ 2.372e+11Hz -0.257309 -0.941243
+ 2.373e+11Hz -0.258049 -0.941058
+ 2.374e+11Hz -0.258788 -0.940872
+ 2.375e+11Hz -0.259527 -0.940685
+ 2.376e+11Hz -0.260267 -0.940497
+ 2.377e+11Hz -0.261006 -0.940309
+ 2.378e+11Hz -0.261746 -0.94012
+ 2.379e+11Hz -0.262485 -0.93993
+ 2.38e+11Hz -0.263225 -0.939739
+ 2.381e+11Hz -0.263964 -0.939547
+ 2.382e+11Hz -0.264704 -0.939354
+ 2.383e+11Hz -0.265443 -0.939161
+ 2.384e+11Hz -0.266183 -0.938966
+ 2.385e+11Hz -0.266923 -0.938771
+ 2.386e+11Hz -0.267662 -0.938575
+ 2.387e+11Hz -0.268402 -0.938378
+ 2.388e+11Hz -0.269141 -0.938181
+ 2.389e+11Hz -0.26988 -0.937982
+ 2.39e+11Hz -0.27062 -0.937783
+ 2.391e+11Hz -0.271359 -0.937582
+ 2.392e+11Hz -0.272098 -0.937381
+ 2.393e+11Hz -0.272838 -0.937179
+ 2.394e+11Hz -0.273577 -0.936976
+ 2.395e+11Hz -0.274316 -0.936773
+ 2.396e+11Hz -0.275055 -0.936568
+ 2.397e+11Hz -0.275794 -0.936363
+ 2.398e+11Hz -0.276533 -0.936157
+ 2.399e+11Hz -0.277272 -0.93595
+ 2.4e+11Hz -0.27801 -0.935742
+ 2.401e+11Hz -0.278749 -0.935533
+ 2.402e+11Hz -0.279487 -0.935324
+ 2.403e+11Hz -0.280226 -0.935113
+ 2.404e+11Hz -0.280964 -0.934902
+ 2.405e+11Hz -0.281702 -0.93469
+ 2.406e+11Hz -0.28244 -0.934477
+ 2.407e+11Hz -0.283178 -0.934263
+ 2.408e+11Hz -0.283916 -0.934048
+ 2.409e+11Hz -0.284653 -0.933833
+ 2.41e+11Hz -0.285391 -0.933617
+ 2.411e+11Hz -0.286128 -0.933399
+ 2.412e+11Hz -0.286865 -0.933181
+ 2.413e+11Hz -0.287602 -0.932963
+ 2.414e+11Hz -0.288339 -0.932743
+ 2.415e+11Hz -0.289076 -0.932522
+ 2.416e+11Hz -0.289812 -0.932301
+ 2.417e+11Hz -0.290549 -0.932079
+ 2.418e+11Hz -0.291285 -0.931856
+ 2.419e+11Hz -0.292021 -0.931632
+ 2.42e+11Hz -0.292756 -0.931407
+ 2.421e+11Hz -0.293492 -0.931182
+ 2.422e+11Hz -0.294227 -0.930956
+ 2.423e+11Hz -0.294962 -0.930728
+ 2.424e+11Hz -0.295697 -0.930501
+ 2.425e+11Hz -0.296432 -0.930272
+ 2.426e+11Hz -0.297166 -0.930042
+ 2.427e+11Hz -0.297901 -0.929812
+ 2.428e+11Hz -0.298635 -0.929581
+ 2.429e+11Hz -0.299368 -0.929349
+ 2.43e+11Hz -0.300102 -0.929116
+ 2.431e+11Hz -0.300835 -0.928882
+ 2.432e+11Hz -0.301568 -0.928648
+ 2.433e+11Hz -0.302301 -0.928413
+ 2.434e+11Hz -0.303034 -0.928177
+ 2.435e+11Hz -0.303766 -0.92794
+ 2.436e+11Hz -0.304498 -0.927703
+ 2.437e+11Hz -0.30523 -0.927464
+ 2.438e+11Hz -0.305962 -0.927225
+ 2.439e+11Hz -0.306693 -0.926985
+ 2.44e+11Hz -0.307424 -0.926745
+ 2.441e+11Hz -0.308155 -0.926503
+ 2.442e+11Hz -0.308885 -0.926261
+ 2.443e+11Hz -0.309616 -0.926018
+ 2.444e+11Hz -0.310345 -0.925774
+ 2.445e+11Hz -0.311075 -0.92553
+ 2.446e+11Hz -0.311805 -0.925285
+ 2.447e+11Hz -0.312534 -0.925039
+ 2.448e+11Hz -0.313262 -0.924792
+ 2.449e+11Hz -0.313991 -0.924545
+ 2.45e+11Hz -0.314719 -0.924296
+ 2.451e+11Hz -0.315447 -0.924047
+ 2.452e+11Hz -0.316175 -0.923798
+ 2.453e+11Hz -0.316902 -0.923547
+ 2.454e+11Hz -0.317629 -0.923296
+ 2.455e+11Hz -0.318356 -0.923044
+ 2.456e+11Hz -0.319082 -0.922791
+ 2.457e+11Hz -0.319808 -0.922538
+ 2.458e+11Hz -0.320534 -0.922284
+ 2.459e+11Hz -0.321259 -0.922029
+ 2.46e+11Hz -0.321985 -0.921774
+ 2.461e+11Hz -0.32271 -0.921517
+ 2.462e+11Hz -0.323434 -0.92126
+ 2.463e+11Hz -0.324158 -0.921003
+ 2.464e+11Hz -0.324882 -0.920744
+ 2.465e+11Hz -0.325606 -0.920485
+ 2.466e+11Hz -0.326329 -0.920225
+ 2.467e+11Hz -0.327052 -0.919965
+ 2.468e+11Hz -0.327775 -0.919704
+ 2.469e+11Hz -0.328497 -0.919442
+ 2.47e+11Hz -0.329219 -0.919179
+ 2.471e+11Hz -0.329941 -0.918916
+ 2.472e+11Hz -0.330662 -0.918652
+ 2.473e+11Hz -0.331383 -0.918388
+ 2.474e+11Hz -0.332103 -0.918122
+ 2.475e+11Hz -0.332824 -0.917856
+ 2.476e+11Hz -0.333544 -0.91759
+ 2.477e+11Hz -0.334264 -0.917322
+ 2.478e+11Hz -0.334983 -0.917054
+ 2.479e+11Hz -0.335702 -0.916786
+ 2.48e+11Hz -0.336421 -0.916516
+ 2.481e+11Hz -0.337139 -0.916247
+ 2.482e+11Hz -0.337857 -0.915976
+ 2.483e+11Hz -0.338575 -0.915705
+ 2.484e+11Hz -0.339292 -0.915433
+ 2.485e+11Hz -0.340009 -0.91516
+ 2.486e+11Hz -0.340726 -0.914887
+ 2.487e+11Hz -0.341442 -0.914613
+ 2.488e+11Hz -0.342158 -0.914338
+ 2.489e+11Hz -0.342874 -0.914063
+ 2.49e+11Hz -0.343589 -0.913787
+ 2.491e+11Hz -0.344304 -0.913511
+ 2.492e+11Hz -0.345019 -0.913234
+ 2.493e+11Hz -0.345733 -0.912956
+ 2.494e+11Hz -0.346447 -0.912678
+ 2.495e+11Hz -0.347161 -0.912399
+ 2.496e+11Hz -0.347874 -0.912119
+ 2.497e+11Hz -0.348587 -0.911839
+ 2.498e+11Hz -0.3493 -0.911558
+ 2.499e+11Hz -0.350012 -0.911276
+ 2.5e+11Hz -0.350724 -0.910994
+ 2.501e+11Hz -0.351436 -0.910712
+ 2.502e+11Hz -0.352147 -0.910428
+ 2.503e+11Hz -0.352858 -0.910144
+ 2.504e+11Hz -0.353569 -0.909859
+ 2.505e+11Hz -0.354279 -0.909574
+ 2.506e+11Hz -0.354989 -0.909288
+ 2.507e+11Hz -0.355699 -0.909002
+ 2.508e+11Hz -0.356408 -0.908715
+ 2.509e+11Hz -0.357117 -0.908427
+ 2.51e+11Hz -0.357826 -0.908139
+ 2.511e+11Hz -0.358534 -0.90785
+ 2.512e+11Hz -0.359242 -0.90756
+ 2.513e+11Hz -0.35995 -0.90727
+ 2.514e+11Hz -0.360657 -0.906979
+ 2.515e+11Hz -0.361364 -0.906688
+ 2.516e+11Hz -0.36207 -0.906396
+ 2.517e+11Hz -0.362777 -0.906103
+ 2.518e+11Hz -0.363483 -0.90581
+ 2.519e+11Hz -0.364188 -0.905516
+ 2.52e+11Hz -0.364894 -0.905221
+ 2.521e+11Hz -0.365598 -0.904926
+ 2.522e+11Hz -0.366303 -0.904631
+ 2.523e+11Hz -0.367007 -0.904334
+ 2.524e+11Hz -0.367711 -0.904038
+ 2.525e+11Hz -0.368415 -0.90374
+ 2.526e+11Hz -0.369118 -0.903442
+ 2.527e+11Hz -0.369821 -0.903143
+ 2.528e+11Hz -0.370523 -0.902844
+ 2.529e+11Hz -0.371226 -0.902544
+ 2.53e+11Hz -0.371928 -0.902244
+ 2.531e+11Hz -0.372629 -0.901943
+ 2.532e+11Hz -0.37333 -0.901641
+ 2.533e+11Hz -0.374031 -0.901339
+ 2.534e+11Hz -0.374732 -0.901036
+ 2.535e+11Hz -0.375432 -0.900732
+ 2.536e+11Hz -0.376131 -0.900428
+ 2.537e+11Hz -0.376831 -0.900123
+ 2.538e+11Hz -0.37753 -0.899818
+ 2.539e+11Hz -0.378229 -0.899512
+ 2.54e+11Hz -0.378927 -0.899206
+ 2.541e+11Hz -0.379625 -0.898899
+ 2.542e+11Hz -0.380323 -0.898591
+ 2.543e+11Hz -0.38102 -0.898283
+ 2.544e+11Hz -0.381717 -0.897974
+ 2.545e+11Hz -0.382414 -0.897664
+ 2.546e+11Hz -0.38311 -0.897354
+ 2.547e+11Hz -0.383806 -0.897044
+ 2.548e+11Hz -0.384502 -0.896732
+ 2.549e+11Hz -0.385197 -0.896421
+ 2.55e+11Hz -0.385892 -0.896108
+ 2.551e+11Hz -0.386586 -0.895795
+ 2.552e+11Hz -0.38728 -0.895481
+ 2.553e+11Hz -0.387974 -0.895167
+ 2.554e+11Hz -0.388667 -0.894852
+ 2.555e+11Hz -0.38936 -0.894537
+ 2.556e+11Hz -0.390053 -0.894221
+ 2.557e+11Hz -0.390745 -0.893904
+ 2.558e+11Hz -0.391437 -0.893587
+ 2.559e+11Hz -0.392128 -0.893269
+ 2.56e+11Hz -0.392819 -0.892951
+ 2.561e+11Hz -0.39351 -0.892632
+ 2.562e+11Hz -0.3942 -0.892312
+ 2.563e+11Hz -0.39489 -0.891992
+ 2.564e+11Hz -0.39558 -0.891672
+ 2.565e+11Hz -0.396269 -0.89135
+ 2.566e+11Hz -0.396958 -0.891028
+ 2.567e+11Hz -0.397646 -0.890706
+ 2.568e+11Hz -0.398334 -0.890383
+ 2.569e+11Hz -0.399022 -0.890059
+ 2.57e+11Hz -0.399709 -0.889735
+ 2.571e+11Hz -0.400396 -0.88941
+ 2.572e+11Hz -0.401082 -0.889085
+ 2.573e+11Hz -0.401768 -0.888759
+ 2.574e+11Hz -0.402454 -0.888432
+ 2.575e+11Hz -0.403139 -0.888105
+ 2.576e+11Hz -0.403824 -0.887778
+ 2.577e+11Hz -0.404508 -0.887449
+ 2.578e+11Hz -0.405192 -0.887121
+ 2.579e+11Hz -0.405875 -0.886791
+ 2.58e+11Hz -0.406558 -0.886461
+ 2.581e+11Hz -0.407241 -0.886131
+ 2.582e+11Hz -0.407923 -0.8858
+ 2.583e+11Hz -0.408605 -0.885468
+ 2.584e+11Hz -0.409286 -0.885136
+ 2.585e+11Hz -0.409967 -0.884803
+ 2.586e+11Hz -0.410648 -0.88447
+ 2.587e+11Hz -0.411328 -0.884136
+ 2.588e+11Hz -0.412007 -0.883802
+ 2.589e+11Hz -0.412686 -0.883467
+ 2.59e+11Hz -0.413365 -0.883131
+ 2.591e+11Hz -0.414043 -0.882795
+ 2.592e+11Hz -0.414721 -0.882458
+ 2.593e+11Hz -0.415398 -0.882121
+ 2.594e+11Hz -0.416075 -0.881784
+ 2.595e+11Hz -0.416752 -0.881446
+ 2.596e+11Hz -0.417428 -0.881107
+ 2.597e+11Hz -0.418103 -0.880768
+ 2.598e+11Hz -0.418778 -0.880428
+ 2.599e+11Hz -0.419453 -0.880088
+ 2.6e+11Hz -0.420127 -0.879747
+ 2.601e+11Hz -0.420801 -0.879405
+ 2.602e+11Hz -0.421474 -0.879064
+ 2.603e+11Hz -0.422146 -0.878721
+ 2.604e+11Hz -0.422819 -0.878379
+ 2.605e+11Hz -0.42349 -0.878035
+ 2.606e+11Hz -0.424162 -0.877691
+ 2.607e+11Hz -0.424832 -0.877347
+ 2.608e+11Hz -0.425503 -0.877002
+ 2.609e+11Hz -0.426173 -0.876657
+ 2.61e+11Hz -0.426842 -0.876311
+ 2.611e+11Hz -0.427511 -0.875965
+ 2.612e+11Hz -0.428179 -0.875618
+ 2.613e+11Hz -0.428847 -0.875271
+ 2.614e+11Hz -0.429514 -0.874923
+ 2.615e+11Hz -0.430181 -0.874575
+ 2.616e+11Hz -0.430847 -0.874227
+ 2.617e+11Hz -0.431513 -0.873878
+ 2.618e+11Hz -0.432179 -0.873528
+ 2.619e+11Hz -0.432843 -0.873178
+ 2.62e+11Hz -0.433508 -0.872828
+ 2.621e+11Hz -0.434172 -0.872477
+ 2.622e+11Hz -0.434835 -0.872126
+ 2.623e+11Hz -0.435498 -0.871774
+ 2.624e+11Hz -0.43616 -0.871422
+ 2.625e+11Hz -0.436822 -0.87107
+ 2.626e+11Hz -0.437484 -0.870717
+ 2.627e+11Hz -0.438144 -0.870364
+ 2.628e+11Hz -0.438805 -0.87001
+ 2.629e+11Hz -0.439465 -0.869656
+ 2.63e+11Hz -0.440124 -0.869301
+ 2.631e+11Hz -0.440783 -0.868947
+ 2.632e+11Hz -0.441441 -0.868591
+ 2.633e+11Hz -0.442099 -0.868236
+ 2.634e+11Hz -0.442756 -0.86788
+ 2.635e+11Hz -0.443413 -0.867523
+ 2.636e+11Hz -0.444069 -0.867167
+ 2.637e+11Hz -0.444725 -0.86681
+ 2.638e+11Hz -0.44538 -0.866452
+ 2.639e+11Hz -0.446035 -0.866094
+ 2.64e+11Hz -0.44669 -0.865736
+ 2.641e+11Hz -0.447343 -0.865378
+ 2.642e+11Hz -0.447997 -0.865019
+ 2.643e+11Hz -0.448649 -0.86466
+ 2.644e+11Hz -0.449302 -0.8643
+ 2.645e+11Hz -0.449954 -0.863941
+ 2.646e+11Hz -0.450605 -0.863581
+ 2.647e+11Hz -0.451256 -0.86322
+ 2.648e+11Hz -0.451906 -0.86286
+ 2.649e+11Hz -0.452556 -0.862499
+ 2.65e+11Hz -0.453205 -0.862137
+ 2.651e+11Hz -0.453854 -0.861776
+ 2.652e+11Hz -0.454503 -0.861414
+ 2.653e+11Hz -0.455151 -0.861052
+ 2.654e+11Hz -0.455798 -0.86069
+ 2.655e+11Hz -0.456445 -0.860327
+ 2.656e+11Hz -0.457092 -0.859964
+ 2.657e+11Hz -0.457738 -0.859601
+ 2.658e+11Hz -0.458384 -0.859238
+ 2.659e+11Hz -0.459029 -0.858874
+ 2.66e+11Hz -0.459673 -0.85851
+ 2.661e+11Hz -0.460318 -0.858146
+ 2.662e+11Hz -0.460962 -0.857782
+ 2.663e+11Hz -0.461605 -0.857418
+ 2.664e+11Hz -0.462248 -0.857053
+ 2.665e+11Hz -0.46289 -0.856688
+ 2.666e+11Hz -0.463532 -0.856323
+ 2.667e+11Hz -0.464174 -0.855957
+ 2.668e+11Hz -0.464815 -0.855592
+ 2.669e+11Hz -0.465456 -0.855226
+ 2.67e+11Hz -0.466097 -0.85486
+ 2.671e+11Hz -0.466737 -0.854494
+ 2.672e+11Hz -0.467376 -0.854128
+ 2.673e+11Hz -0.468015 -0.853761
+ 2.674e+11Hz -0.468654 -0.853395
+ 2.675e+11Hz -0.469293 -0.853028
+ 2.676e+11Hz -0.469931 -0.852661
+ 2.677e+11Hz -0.470568 -0.852293
+ 2.678e+11Hz -0.471205 -0.851926
+ 2.679e+11Hz -0.471842 -0.851559
+ 2.68e+11Hz -0.472479 -0.851191
+ 2.681e+11Hz -0.473115 -0.850823
+ 2.682e+11Hz -0.473751 -0.850455
+ 2.683e+11Hz -0.474386 -0.850087
+ 2.684e+11Hz -0.475022 -0.849719
+ 2.685e+11Hz -0.475656 -0.849351
+ 2.686e+11Hz -0.476291 -0.848982
+ 2.687e+11Hz -0.476925 -0.848613
+ 2.688e+11Hz -0.477559 -0.848245
+ 2.689e+11Hz -0.478193 -0.847876
+ 2.69e+11Hz -0.478826 -0.847507
+ 2.691e+11Hz -0.479459 -0.847138
+ 2.692e+11Hz -0.480091 -0.846768
+ 2.693e+11Hz -0.480724 -0.846399
+ 2.694e+11Hz -0.481356 -0.846029
+ 2.695e+11Hz -0.481988 -0.84566
+ 2.696e+11Hz -0.482619 -0.84529
+ 2.697e+11Hz -0.483251 -0.84492
+ 2.698e+11Hz -0.483882 -0.84455
+ 2.699e+11Hz -0.484513 -0.84418
+ 2.7e+11Hz -0.485143 -0.84381
+ 2.701e+11Hz -0.485774 -0.84344
+ 2.702e+11Hz -0.486404 -0.843069
+ 2.703e+11Hz -0.487034 -0.842699
+ 2.704e+11Hz -0.487664 -0.842328
+ 2.705e+11Hz -0.488293 -0.841957
+ 2.706e+11Hz -0.488923 -0.841586
+ 2.707e+11Hz -0.489552 -0.841215
+ 2.708e+11Hz -0.490181 -0.840844
+ 2.709e+11Hz -0.49081 -0.840473
+ 2.71e+11Hz -0.491439 -0.840102
+ 2.711e+11Hz -0.492067 -0.83973
+ 2.712e+11Hz -0.492696 -0.839359
+ 2.713e+11Hz -0.493324 -0.838987
+ 2.714e+11Hz -0.493952 -0.838615
+ 2.715e+11Hz -0.49458 -0.838243
+ 2.716e+11Hz -0.495208 -0.837871
+ 2.717e+11Hz -0.495836 -0.837499
+ 2.718e+11Hz -0.496464 -0.837127
+ 2.719e+11Hz -0.497092 -0.836754
+ 2.72e+11Hz -0.497719 -0.836382
+ 2.721e+11Hz -0.498347 -0.836009
+ 2.722e+11Hz -0.498974 -0.835636
+ 2.723e+11Hz -0.499601 -0.835263
+ 2.724e+11Hz -0.500229 -0.83489
+ 2.725e+11Hz -0.500856 -0.834517
+ 2.726e+11Hz -0.501483 -0.834144
+ 2.727e+11Hz -0.50211 -0.83377
+ 2.728e+11Hz -0.502738 -0.833396
+ 2.729e+11Hz -0.503365 -0.833022
+ 2.73e+11Hz -0.503992 -0.832648
+ 2.731e+11Hz -0.504619 -0.832274
+ 2.732e+11Hz -0.505246 -0.8319
+ 2.733e+11Hz -0.505873 -0.831525
+ 2.734e+11Hz -0.5065 -0.83115
+ 2.735e+11Hz -0.507127 -0.830775
+ 2.736e+11Hz -0.507755 -0.8304
+ 2.737e+11Hz -0.508382 -0.830025
+ 2.738e+11Hz -0.509009 -0.829649
+ 2.739e+11Hz -0.509636 -0.829273
+ 2.74e+11Hz -0.510264 -0.828897
+ 2.741e+11Hz -0.510891 -0.828521
+ 2.742e+11Hz -0.511519 -0.828145
+ 2.743e+11Hz -0.512146 -0.827768
+ 2.744e+11Hz -0.512774 -0.827391
+ 2.745e+11Hz -0.513401 -0.827014
+ 2.746e+11Hz -0.514029 -0.826636
+ 2.747e+11Hz -0.514657 -0.826259
+ 2.748e+11Hz -0.515285 -0.825881
+ 2.749e+11Hz -0.515913 -0.825502
+ 2.75e+11Hz -0.516541 -0.825124
+ 2.751e+11Hz -0.517169 -0.824745
+ 2.752e+11Hz -0.517798 -0.824366
+ 2.753e+11Hz -0.518426 -0.823987
+ 2.754e+11Hz -0.519055 -0.823607
+ 2.755e+11Hz -0.519683 -0.823227
+ 2.756e+11Hz -0.520312 -0.822846
+ 2.757e+11Hz -0.520941 -0.822466
+ 2.758e+11Hz -0.52157 -0.822084
+ 2.759e+11Hz -0.522199 -0.821703
+ 2.76e+11Hz -0.522829 -0.821321
+ 2.761e+11Hz -0.523458 -0.820939
+ 2.762e+11Hz -0.524088 -0.820556
+ 2.763e+11Hz -0.524718 -0.820174
+ 2.764e+11Hz -0.525348 -0.81979
+ 2.765e+11Hz -0.525978 -0.819406
+ 2.766e+11Hz -0.526608 -0.819022
+ 2.767e+11Hz -0.527238 -0.818638
+ 2.768e+11Hz -0.527869 -0.818253
+ 2.769e+11Hz -0.5285 -0.817867
+ 2.77e+11Hz -0.529131 -0.817481
+ 2.771e+11Hz -0.529762 -0.817095
+ 2.772e+11Hz -0.530393 -0.816708
+ 2.773e+11Hz -0.531024 -0.816321
+ 2.774e+11Hz -0.531656 -0.815933
+ 2.775e+11Hz -0.532287 -0.815545
+ 2.776e+11Hz -0.532919 -0.815156
+ 2.777e+11Hz -0.533551 -0.814767
+ 2.778e+11Hz -0.534184 -0.814377
+ 2.779e+11Hz -0.534816 -0.813987
+ 2.78e+11Hz -0.535448 -0.813596
+ 2.781e+11Hz -0.536081 -0.813205
+ 2.782e+11Hz -0.536714 -0.812813
+ 2.783e+11Hz -0.537347 -0.81242
+ 2.784e+11Hz -0.53798 -0.812027
+ 2.785e+11Hz -0.538613 -0.811633
+ 2.786e+11Hz -0.539247 -0.811239
+ 2.787e+11Hz -0.53988 -0.810844
+ 2.788e+11Hz -0.540514 -0.810449
+ 2.789e+11Hz -0.541148 -0.810053
+ 2.79e+11Hz -0.541782 -0.809656
+ 2.791e+11Hz -0.542416 -0.809258
+ 2.792e+11Hz -0.54305 -0.80886
+ 2.793e+11Hz -0.543685 -0.808462
+ 2.794e+11Hz -0.544319 -0.808062
+ 2.795e+11Hz -0.544954 -0.807662
+ 2.796e+11Hz -0.545589 -0.807262
+ 2.797e+11Hz -0.546224 -0.80686
+ 2.798e+11Hz -0.546859 -0.806458
+ 2.799e+11Hz -0.547494 -0.806055
+ 2.8e+11Hz -0.548129 -0.805652
+ 2.801e+11Hz -0.548765 -0.805248
+ 2.802e+11Hz -0.5494 -0.804843
+ 2.803e+11Hz -0.550036 -0.804437
+ 2.804e+11Hz -0.550671 -0.804031
+ 2.805e+11Hz -0.551307 -0.803623
+ 2.806e+11Hz -0.551943 -0.803215
+ 2.807e+11Hz -0.552579 -0.802807
+ 2.808e+11Hz -0.553215 -0.802397
+ 2.809e+11Hz -0.553851 -0.801987
+ 2.81e+11Hz -0.554487 -0.801576
+ 2.811e+11Hz -0.555123 -0.801164
+ 2.812e+11Hz -0.555759 -0.800751
+ 2.813e+11Hz -0.556395 -0.800338
+ 2.814e+11Hz -0.557031 -0.799923
+ 2.815e+11Hz -0.557667 -0.799508
+ 2.816e+11Hz -0.558303 -0.799092
+ 2.817e+11Hz -0.55894 -0.798675
+ 2.818e+11Hz -0.559576 -0.798258
+ 2.819e+11Hz -0.560212 -0.797839
+ 2.82e+11Hz -0.560848 -0.79742
+ 2.821e+11Hz -0.561484 -0.797
+ 2.822e+11Hz -0.56212 -0.796579
+ 2.823e+11Hz -0.562756 -0.796157
+ 2.824e+11Hz -0.563392 -0.795734
+ 2.825e+11Hz -0.564028 -0.79531
+ 2.826e+11Hz -0.564664 -0.794885
+ 2.827e+11Hz -0.5653 -0.79446
+ 2.828e+11Hz -0.565935 -0.794033
+ 2.829e+11Hz -0.566571 -0.793606
+ 2.83e+11Hz -0.567207 -0.793178
+ 2.831e+11Hz -0.567842 -0.792749
+ 2.832e+11Hz -0.568477 -0.792319
+ 2.833e+11Hz -0.569112 -0.791888
+ 2.834e+11Hz -0.569747 -0.791456
+ 2.835e+11Hz -0.570382 -0.791023
+ 2.836e+11Hz -0.571017 -0.790589
+ 2.837e+11Hz -0.571651 -0.790155
+ 2.838e+11Hz -0.572285 -0.789719
+ 2.839e+11Hz -0.572919 -0.789283
+ 2.84e+11Hz -0.573553 -0.788845
+ 2.841e+11Hz -0.574187 -0.788407
+ 2.842e+11Hz -0.57482 -0.787968
+ 2.843e+11Hz -0.575454 -0.787527
+ 2.844e+11Hz -0.576087 -0.787086
+ 2.845e+11Hz -0.57672 -0.786644
+ 2.846e+11Hz -0.577352 -0.786201
+ 2.847e+11Hz -0.577984 -0.785757
+ 2.848e+11Hz -0.578616 -0.785312
+ 2.849e+11Hz -0.579248 -0.784866
+ 2.85e+11Hz -0.579879 -0.784419
+ 2.851e+11Hz -0.58051 -0.783972
+ 2.852e+11Hz -0.581141 -0.783523
+ 2.853e+11Hz -0.581772 -0.783073
+ 2.854e+11Hz -0.582402 -0.782623
+ 2.855e+11Hz -0.583032 -0.782171
+ 2.856e+11Hz -0.583661 -0.781719
+ 2.857e+11Hz -0.58429 -0.781265
+ 2.858e+11Hz -0.584919 -0.780811
+ 2.859e+11Hz -0.585547 -0.780356
+ 2.86e+11Hz -0.586175 -0.779899
+ 2.861e+11Hz -0.586802 -0.779442
+ 2.862e+11Hz -0.58743 -0.778984
+ 2.863e+11Hz -0.588056 -0.778525
+ 2.864e+11Hz -0.588683 -0.778065
+ 2.865e+11Hz -0.589308 -0.777605
+ 2.866e+11Hz -0.589934 -0.777143
+ 2.867e+11Hz -0.590559 -0.77668
+ 2.868e+11Hz -0.591183 -0.776217
+ 2.869e+11Hz -0.591807 -0.775752
+ 2.87e+11Hz -0.592431 -0.775287
+ 2.871e+11Hz -0.593054 -0.77482
+ 2.872e+11Hz -0.593677 -0.774353
+ 2.873e+11Hz -0.594299 -0.773885
+ 2.874e+11Hz -0.59492 -0.773416
+ 2.875e+11Hz -0.595541 -0.772947
+ 2.876e+11Hz -0.596162 -0.772476
+ 2.877e+11Hz -0.596782 -0.772004
+ 2.878e+11Hz -0.597401 -0.771532
+ 2.879e+11Hz -0.59802 -0.771059
+ 2.88e+11Hz -0.598638 -0.770585
+ 2.881e+11Hz -0.599256 -0.77011
+ 2.882e+11Hz -0.599873 -0.769634
+ 2.883e+11Hz -0.60049 -0.769157
+ 2.884e+11Hz -0.601106 -0.76868
+ 2.885e+11Hz -0.601722 -0.768201
+ 2.886e+11Hz -0.602336 -0.767722
+ 2.887e+11Hz -0.602951 -0.767242
+ 2.888e+11Hz -0.603564 -0.766762
+ 2.889e+11Hz -0.604177 -0.76628
+ 2.89e+11Hz -0.60479 -0.765798
+ 2.891e+11Hz -0.605402 -0.765315
+ 2.892e+11Hz -0.606013 -0.764831
+ 2.893e+11Hz -0.606623 -0.764346
+ 2.894e+11Hz -0.607233 -0.763861
+ 2.895e+11Hz -0.607843 -0.763374
+ 2.896e+11Hz -0.608451 -0.762888
+ 2.897e+11Hz -0.609059 -0.7624
+ 2.898e+11Hz -0.609666 -0.761911
+ 2.899e+11Hz -0.610273 -0.761422
+ 2.9e+11Hz -0.610879 -0.760932
+ 2.901e+11Hz -0.611484 -0.760442
+ 2.902e+11Hz -0.612089 -0.759951
+ 2.903e+11Hz -0.612693 -0.759459
+ 2.904e+11Hz -0.613296 -0.758966
+ 2.905e+11Hz -0.613899 -0.758473
+ 2.906e+11Hz -0.614501 -0.757978
+ 2.907e+11Hz -0.615102 -0.757484
+ 2.908e+11Hz -0.615703 -0.756988
+ 2.909e+11Hz -0.616302 -0.756492
+ 2.91e+11Hz -0.616902 -0.755996
+ 2.911e+11Hz -0.6175 -0.755498
+ 2.912e+11Hz -0.618098 -0.755
+ 2.913e+11Hz -0.618695 -0.754502
+ 2.914e+11Hz -0.619291 -0.754003
+ 2.915e+11Hz -0.619887 -0.753503
+ 2.916e+11Hz -0.620482 -0.753003
+ 2.917e+11Hz -0.621076 -0.752502
+ 2.918e+11Hz -0.62167 -0.752
+ 2.919e+11Hz -0.622262 -0.751498
+ 2.92e+11Hz -0.622855 -0.750995
+ 2.921e+11Hz -0.623446 -0.750492
+ 2.922e+11Hz -0.624037 -0.749988
+ 2.923e+11Hz -0.624627 -0.749484
+ 2.924e+11Hz -0.625216 -0.748979
+ 2.925e+11Hz -0.625805 -0.748473
+ 2.926e+11Hz -0.626392 -0.747967
+ 2.927e+11Hz -0.62698 -0.747461
+ 2.928e+11Hz -0.627566 -0.746954
+ 2.929e+11Hz -0.628152 -0.746446
+ 2.93e+11Hz -0.628737 -0.745938
+ 2.931e+11Hz -0.629322 -0.74543
+ 2.932e+11Hz -0.629905 -0.744921
+ 2.933e+11Hz -0.630488 -0.744411
+ 2.934e+11Hz -0.631071 -0.743901
+ 2.935e+11Hz -0.631652 -0.743391
+ 2.936e+11Hz -0.632233 -0.74288
+ 2.937e+11Hz -0.632813 -0.742369
+ 2.938e+11Hz -0.633393 -0.741857
+ 2.939e+11Hz -0.633972 -0.741345
+ 2.94e+11Hz -0.63455 -0.740832
+ 2.941e+11Hz -0.635128 -0.740319
+ 2.942e+11Hz -0.635705 -0.739805
+ 2.943e+11Hz -0.636281 -0.739291
+ 2.944e+11Hz -0.636856 -0.738777
+ 2.945e+11Hz -0.637431 -0.738262
+ 2.946e+11Hz -0.638005 -0.737747
+ 2.947e+11Hz -0.638579 -0.737231
+ 2.948e+11Hz -0.639152 -0.736716
+ 2.949e+11Hz -0.639724 -0.736199
+ 2.95e+11Hz -0.640296 -0.735682
+ 2.951e+11Hz -0.640867 -0.735165
+ 2.952e+11Hz -0.641437 -0.734648
+ 2.953e+11Hz -0.642007 -0.73413
+ 2.954e+11Hz -0.642576 -0.733612
+ 2.955e+11Hz -0.643144 -0.733093
+ 2.956e+11Hz -0.643712 -0.732574
+ 2.957e+11Hz -0.644279 -0.732055
+ 2.958e+11Hz -0.644846 -0.731535
+ 2.959e+11Hz -0.645412 -0.731015
+ 2.96e+11Hz -0.645978 -0.730494
+ 2.961e+11Hz -0.646542 -0.729974
+ 2.962e+11Hz -0.647107 -0.729452
+ 2.963e+11Hz -0.64767 -0.728931
+ 2.964e+11Hz -0.648233 -0.728409
+ 2.965e+11Hz -0.648796 -0.727887
+ 2.966e+11Hz -0.649358 -0.727364
+ 2.967e+11Hz -0.649919 -0.726842
+ 2.968e+11Hz -0.65048 -0.726318
+ 2.969e+11Hz -0.65104 -0.725795
+ 2.97e+11Hz -0.651599 -0.725271
+ 2.971e+11Hz -0.652158 -0.724747
+ 2.972e+11Hz -0.652717 -0.724222
+ 2.973e+11Hz -0.653275 -0.723698
+ 2.974e+11Hz -0.653832 -0.723172
+ 2.975e+11Hz -0.654389 -0.722647
+ 2.976e+11Hz -0.654946 -0.722121
+ 2.977e+11Hz -0.655501 -0.721595
+ 2.978e+11Hz -0.656057 -0.721069
+ 2.979e+11Hz -0.656612 -0.720542
+ 2.98e+11Hz -0.657166 -0.720015
+ 2.981e+11Hz -0.65772 -0.719487
+ 2.982e+11Hz -0.658273 -0.718959
+ 2.983e+11Hz -0.658826 -0.718431
+ 2.984e+11Hz -0.659378 -0.717903
+ 2.985e+11Hz -0.659929 -0.717374
+ 2.986e+11Hz -0.660481 -0.716845
+ 2.987e+11Hz -0.661031 -0.716316
+ 2.988e+11Hz -0.661582 -0.715786
+ 2.989e+11Hz -0.662131 -0.715256
+ 2.99e+11Hz -0.662681 -0.714725
+ 2.991e+11Hz -0.66323 -0.714194
+ 2.992e+11Hz -0.663778 -0.713663
+ 2.993e+11Hz -0.664326 -0.713132
+ 2.994e+11Hz -0.664873 -0.7126
+ 2.995e+11Hz -0.66542 -0.712068
+ 2.996e+11Hz -0.665967 -0.711535
+ 2.997e+11Hz -0.666513 -0.711002
+ 2.998e+11Hz -0.667058 -0.710469
+ 2.999e+11Hz -0.667603 -0.709936
+ 3e+11Hz -0.668148 -0.709402
+ ]

A22 %vd(20 3) %vd(22, 3) xfer4
.model xfer4 xfer R_I=true table=[
+ 0Hz 0.0047718 0
+ 1e+08Hz 0.00477202 3.3416e-06
+ 2e+08Hz 0.00477265 6.6748e-06
+ 3e+08Hz 0.0047737 9.99121e-06
+ 4e+08Hz 0.00477517 1.32825e-05
+ 5e+08Hz 0.00477706 1.65402e-05
+ 6e+08Hz 0.00477937 1.9756e-05
+ 7e+08Hz 0.0047821 2.29215e-05
+ 8e+08Hz 0.00478524 2.60286e-05
+ 9e+08Hz 0.0047888 2.90688e-05
+ 1e+09Hz 0.00479277 3.20341e-05
+ 1.1e+09Hz 0.00479716 3.49161e-05
+ 1.2e+09Hz 0.00480195 3.77067e-05
+ 1.3e+09Hz 0.00480715 4.03978e-05
+ 1.4e+09Hz 0.00481276 4.29814e-05
+ 1.5e+09Hz 0.00481877 4.54495e-05
+ 1.6e+09Hz 0.00482518 4.77941e-05
+ 1.7e+09Hz 0.00483198 5.00074e-05
+ 1.8e+09Hz 0.00483919 5.20816e-05
+ 1.9e+09Hz 0.00484678 5.40089e-05
+ 2e+09Hz 0.00485476 5.57818e-05
+ 2.1e+09Hz 0.00486313 5.73926e-05
+ 2.2e+09Hz 0.00487188 5.88339e-05
+ 2.3e+09Hz 0.00488101 6.00983e-05
+ 2.4e+09Hz 0.00489051 6.11784e-05
+ 2.5e+09Hz 0.00490038 6.20672e-05
+ 2.6e+09Hz 0.00491061 6.27574e-05
+ 2.7e+09Hz 0.00492121 6.32421e-05
+ 2.8e+09Hz 0.00493216 6.35144e-05
+ 2.9e+09Hz 0.00494347 6.35675e-05
+ 3e+09Hz 0.00495512 6.33948e-05
+ 3.1e+09Hz 0.00496711 6.29896e-05
+ 3.2e+09Hz 0.00497945 6.23456e-05
+ 3.3e+09Hz 0.00499211 6.14564e-05
+ 3.4e+09Hz 0.0050051 6.03159e-05
+ 3.5e+09Hz 0.00501841 5.89179e-05
+ 3.6e+09Hz 0.00503204 5.72566e-05
+ 3.7e+09Hz 0.00504598 5.53262e-05
+ 3.8e+09Hz 0.00506022 5.3121e-05
+ 3.9e+09Hz 0.00507476 5.06354e-05
+ 4e+09Hz 0.00508959 4.78642e-05
+ 4.1e+09Hz 0.00510471 4.48019e-05
+ 4.2e+09Hz 0.00512011 4.14436e-05
+ 4.3e+09Hz 0.00513579 3.77843e-05
+ 4.4e+09Hz 0.00515173 3.38191e-05
+ 4.5e+09Hz 0.00516793 2.95435e-05
+ 4.6e+09Hz 0.00518439 2.49528e-05
+ 4.7e+09Hz 0.0052011 2.00428e-05
+ 4.8e+09Hz 0.00521804 1.48093e-05
+ 4.9e+09Hz 0.00523522 9.24808e-06
+ 5e+09Hz 0.00525263 3.3554e-06
+ 5.1e+09Hz 0.00527026 -2.87253e-06
+ 5.2e+09Hz 0.00528811 -9.43928e-06
+ 5.3e+09Hz 0.00530616 -1.63483e-05
+ 5.4e+09Hz 0.00532441 -2.36027e-05
+ 5.5e+09Hz 0.00534285 -3.12058e-05
+ 5.6e+09Hz 0.00536148 -3.91605e-05
+ 5.7e+09Hz 0.00538029 -4.74694e-05
+ 5.8e+09Hz 0.00539927 -5.61353e-05
+ 5.9e+09Hz 0.00541841 -6.51606e-05
+ 6e+09Hz 0.00543771 -7.45476e-05
+ 6.1e+09Hz 0.00545716 -8.42984e-05
+ 6.2e+09Hz 0.00547675 -9.44149e-05
+ 6.3e+09Hz 0.00549648 -0.000104899
+ 6.4e+09Hz 0.00551633 -0.000115753
+ 6.5e+09Hz 0.0055363 -0.000126977
+ 6.6e+09Hz 0.00555639 -0.000138573
+ 6.7e+09Hz 0.00557658 -0.000150542
+ 6.8e+09Hz 0.00559687 -0.000162886
+ 6.9e+09Hz 0.00561724 -0.000175605
+ 7e+09Hz 0.00563771 -0.0001887
+ 7.1e+09Hz 0.00565825 -0.00020217
+ 7.2e+09Hz 0.00567885 -0.000216018
+ 7.3e+09Hz 0.00569952 -0.000230243
+ 7.4e+09Hz 0.00572024 -0.000244844
+ 7.5e+09Hz 0.00574101 -0.000259822
+ 7.6e+09Hz 0.00576182 -0.000275178
+ 7.7e+09Hz 0.00578266 -0.000290909
+ 7.8e+09Hz 0.00580352 -0.000307016
+ 7.9e+09Hz 0.00582441 -0.000323498
+ 8e+09Hz 0.0058453 -0.000340355
+ 8.1e+09Hz 0.0058662 -0.000357584
+ 8.2e+09Hz 0.00588709 -0.000375186
+ 8.3e+09Hz 0.00590798 -0.000393159
+ 8.4e+09Hz 0.00592884 -0.000411502
+ 8.5e+09Hz 0.00594969 -0.000430212
+ 8.6e+09Hz 0.0059705 -0.000449289
+ 8.7e+09Hz 0.00599128 -0.00046873
+ 8.8e+09Hz 0.00601201 -0.000488534
+ 8.9e+09Hz 0.0060327 -0.000508699
+ 9e+09Hz 0.00605332 -0.000529222
+ 9.1e+09Hz 0.00607388 -0.000550101
+ 9.2e+09Hz 0.00609438 -0.000571334
+ 9.3e+09Hz 0.0061148 -0.000592918
+ 9.4e+09Hz 0.00613513 -0.00061485
+ 9.5e+09Hz 0.00615538 -0.000637128
+ 9.6e+09Hz 0.00617553 -0.000659749
+ 9.7e+09Hz 0.00619559 -0.00068271
+ 9.8e+09Hz 0.00621554 -0.000706007
+ 9.9e+09Hz 0.00623537 -0.000729638
+ 1e+10Hz 0.00625509 -0.0007536
+ 1.01e+10Hz 0.00627469 -0.000777888
+ 1.02e+10Hz 0.00629416 -0.000802499
+ 1.03e+10Hz 0.0063135 -0.00082743
+ 1.04e+10Hz 0.0063327 -0.000852677
+ 1.05e+10Hz 0.00635175 -0.000878236
+ 1.06e+10Hz 0.00637065 -0.000904103
+ 1.07e+10Hz 0.00638941 -0.000930275
+ 1.08e+10Hz 0.006408 -0.000956747
+ 1.09e+10Hz 0.00642643 -0.000983515
+ 1.1e+10Hz 0.00644469 -0.00101058
+ 1.11e+10Hz 0.00646278 -0.00103792
+ 1.12e+10Hz 0.00648069 -0.00106555
+ 1.13e+10Hz 0.00649842 -0.00109346
+ 1.14e+10Hz 0.00651597 -0.00112165
+ 1.15e+10Hz 0.00653332 -0.0011501
+ 1.16e+10Hz 0.00655049 -0.00117882
+ 1.17e+10Hz 0.00656745 -0.0012078
+ 1.18e+10Hz 0.00658422 -0.00123704
+ 1.19e+10Hz 0.00660078 -0.00126653
+ 1.2e+10Hz 0.00661713 -0.00129626
+ 1.21e+10Hz 0.00663328 -0.00132624
+ 1.22e+10Hz 0.0066492 -0.00135645
+ 1.23e+10Hz 0.00666491 -0.0013869
+ 1.24e+10Hz 0.0066804 -0.00141757
+ 1.25e+10Hz 0.00669567 -0.00144846
+ 1.26e+10Hz 0.00671071 -0.00147957
+ 1.27e+10Hz 0.00672552 -0.00151089
+ 1.28e+10Hz 0.0067401 -0.00154242
+ 1.29e+10Hz 0.00675444 -0.00157415
+ 1.3e+10Hz 0.00676855 -0.00160607
+ 1.31e+10Hz 0.00678242 -0.00163819
+ 1.32e+10Hz 0.00679605 -0.00167049
+ 1.33e+10Hz 0.00680944 -0.00170297
+ 1.34e+10Hz 0.00682259 -0.00173563
+ 1.35e+10Hz 0.00683548 -0.00176846
+ 1.36e+10Hz 0.00684813 -0.00180146
+ 1.37e+10Hz 0.00686054 -0.00183461
+ 1.38e+10Hz 0.00687269 -0.00186792
+ 1.39e+10Hz 0.00688459 -0.00190138
+ 1.4e+10Hz 0.00689623 -0.00193498
+ 1.41e+10Hz 0.00690763 -0.00196872
+ 1.42e+10Hz 0.00691877 -0.00200259
+ 1.43e+10Hz 0.00692965 -0.0020366
+ 1.44e+10Hz 0.00694028 -0.00207073
+ 1.45e+10Hz 0.00695065 -0.00210497
+ 1.46e+10Hz 0.00696076 -0.00213933
+ 1.47e+10Hz 0.00697062 -0.0021738
+ 1.48e+10Hz 0.00698022 -0.00220837
+ 1.49e+10Hz 0.00698956 -0.00224303
+ 1.5e+10Hz 0.00699865 -0.00227779
+ 1.51e+10Hz 0.00700747 -0.00231264
+ 1.52e+10Hz 0.00701604 -0.00234757
+ 1.53e+10Hz 0.00702435 -0.00238258
+ 1.54e+10Hz 0.00703241 -0.00241767
+ 1.55e+10Hz 0.00704021 -0.00245282
+ 1.56e+10Hz 0.00704775 -0.00248803
+ 1.57e+10Hz 0.00705504 -0.0025233
+ 1.58e+10Hz 0.00706207 -0.00255863
+ 1.59e+10Hz 0.00706885 -0.00259401
+ 1.6e+10Hz 0.00707538 -0.00262943
+ 1.61e+10Hz 0.00708166 -0.00266489
+ 1.62e+10Hz 0.00708769 -0.00270038
+ 1.63e+10Hz 0.00709347 -0.00273591
+ 1.64e+10Hz 0.007099 -0.00277146
+ 1.65e+10Hz 0.00710429 -0.00280704
+ 1.66e+10Hz 0.00710933 -0.00284263
+ 1.67e+10Hz 0.00711413 -0.00287824
+ 1.68e+10Hz 0.00711869 -0.00291386
+ 1.69e+10Hz 0.007123 -0.00294948
+ 1.7e+10Hz 0.00712709 -0.0029851
+ 1.71e+10Hz 0.00713093 -0.00302072
+ 1.72e+10Hz 0.00713454 -0.00305634
+ 1.73e+10Hz 0.00713792 -0.00309194
+ 1.74e+10Hz 0.00714107 -0.00312753
+ 1.75e+10Hz 0.007144 -0.0031631
+ 1.76e+10Hz 0.0071467 -0.00319865
+ 1.77e+10Hz 0.00714917 -0.00323418
+ 1.78e+10Hz 0.00715143 -0.00326967
+ 1.79e+10Hz 0.00715346 -0.00330514
+ 1.8e+10Hz 0.00715529 -0.00334057
+ 1.81e+10Hz 0.0071569 -0.00337596
+ 1.82e+10Hz 0.0071583 -0.00341131
+ 1.83e+10Hz 0.00715949 -0.00344661
+ 1.84e+10Hz 0.00716048 -0.00348187
+ 1.85e+10Hz 0.00716126 -0.00351707
+ 1.86e+10Hz 0.00716185 -0.00355222
+ 1.87e+10Hz 0.00716224 -0.00358732
+ 1.88e+10Hz 0.00716243 -0.00362236
+ 1.89e+10Hz 0.00716244 -0.00365733
+ 1.9e+10Hz 0.00716225 -0.00369224
+ 1.91e+10Hz 0.00716189 -0.00372709
+ 1.92e+10Hz 0.00716134 -0.00376186
+ 1.93e+10Hz 0.00716061 -0.00379657
+ 1.94e+10Hz 0.00715971 -0.0038312
+ 1.95e+10Hz 0.00715863 -0.00386576
+ 1.96e+10Hz 0.00715739 -0.00390024
+ 1.97e+10Hz 0.00715598 -0.00393464
+ 1.98e+10Hz 0.00715441 -0.00396895
+ 1.99e+10Hz 0.00715267 -0.00400319
+ 2e+10Hz 0.00715079 -0.00403734
+ 2.01e+10Hz 0.00714874 -0.00407141
+ 2.02e+10Hz 0.00714655 -0.00410539
+ 2.03e+10Hz 0.00714421 -0.00413928
+ 2.04e+10Hz 0.00714173 -0.00417308
+ 2.05e+10Hz 0.0071391 -0.00420679
+ 2.06e+10Hz 0.00713634 -0.0042404
+ 2.07e+10Hz 0.00713345 -0.00427393
+ 2.08e+10Hz 0.00713043 -0.00430736
+ 2.09e+10Hz 0.00712727 -0.00434069
+ 2.1e+10Hz 0.007124 -0.00437393
+ 2.11e+10Hz 0.0071206 -0.00440707
+ 2.12e+10Hz 0.00711709 -0.00444012
+ 2.13e+10Hz 0.00711346 -0.00447306
+ 2.14e+10Hz 0.00710972 -0.00450591
+ 2.15e+10Hz 0.00710587 -0.00453866
+ 2.16e+10Hz 0.00710192 -0.00457131
+ 2.17e+10Hz 0.00709786 -0.00460386
+ 2.18e+10Hz 0.00709371 -0.00463632
+ 2.19e+10Hz 0.00708946 -0.00466867
+ 2.2e+10Hz 0.00708512 -0.00470093
+ 2.21e+10Hz 0.00708069 -0.00473308
+ 2.22e+10Hz 0.00707617 -0.00476514
+ 2.23e+10Hz 0.00707157 -0.0047971
+ 2.24e+10Hz 0.00706689 -0.00482896
+ 2.25e+10Hz 0.00706213 -0.00486072
+ 2.26e+10Hz 0.0070573 -0.00489238
+ 2.27e+10Hz 0.00705239 -0.00492395
+ 2.28e+10Hz 0.00704742 -0.00495542
+ 2.29e+10Hz 0.00704238 -0.0049868
+ 2.3e+10Hz 0.00703728 -0.00501808
+ 2.31e+10Hz 0.00703211 -0.00504927
+ 2.32e+10Hz 0.00702689 -0.00508036
+ 2.33e+10Hz 0.00702161 -0.00511136
+ 2.34e+10Hz 0.00701628 -0.00514227
+ 2.35e+10Hz 0.0070109 -0.00517309
+ 2.36e+10Hz 0.00700547 -0.00520382
+ 2.37e+10Hz 0.00699999 -0.00523446
+ 2.38e+10Hz 0.00699447 -0.00526501
+ 2.39e+10Hz 0.00698891 -0.00529548
+ 2.4e+10Hz 0.00698331 -0.00532587
+ 2.41e+10Hz 0.00697767 -0.00535617
+ 2.42e+10Hz 0.006972 -0.00538639
+ 2.43e+10Hz 0.0069663 -0.00541653
+ 2.44e+10Hz 0.00696057 -0.00544659
+ 2.45e+10Hz 0.0069548 -0.00547657
+ 2.46e+10Hz 0.00694902 -0.00550648
+ 2.47e+10Hz 0.0069432 -0.00553631
+ 2.48e+10Hz 0.00693737 -0.00556607
+ 2.49e+10Hz 0.00693151 -0.00559576
+ 2.5e+10Hz 0.00692563 -0.00562538
+ 2.51e+10Hz 0.00691974 -0.00565493
+ 2.52e+10Hz 0.00691383 -0.00568442
+ 2.53e+10Hz 0.0069079 -0.00571384
+ 2.54e+10Hz 0.00690196 -0.0057432
+ 2.55e+10Hz 0.00689601 -0.0057725
+ 2.56e+10Hz 0.00689004 -0.00580175
+ 2.57e+10Hz 0.00688407 -0.00583093
+ 2.58e+10Hz 0.00687809 -0.00586006
+ 2.59e+10Hz 0.0068721 -0.00588914
+ 2.6e+10Hz 0.00686611 -0.00591816
+ 2.61e+10Hz 0.00686011 -0.00594714
+ 2.62e+10Hz 0.0068541 -0.00597607
+ 2.63e+10Hz 0.0068481 -0.00600495
+ 2.64e+10Hz 0.00684208 -0.00603379
+ 2.65e+10Hz 0.00683607 -0.00606259
+ 2.66e+10Hz 0.00683006 -0.00609135
+ 2.67e+10Hz 0.00682404 -0.00612007
+ 2.68e+10Hz 0.00681803 -0.00614876
+ 2.69e+10Hz 0.00681201 -0.00617741
+ 2.7e+10Hz 0.006806 -0.00620604
+ 2.71e+10Hz 0.00679998 -0.00623463
+ 2.72e+10Hz 0.00679397 -0.00626319
+ 2.73e+10Hz 0.00678796 -0.00629173
+ 2.74e+10Hz 0.00678195 -0.00632025
+ 2.75e+10Hz 0.00677594 -0.00634874
+ 2.76e+10Hz 0.00676994 -0.00637721
+ 2.77e+10Hz 0.00676394 -0.00640566
+ 2.78e+10Hz 0.00675793 -0.0064341
+ 2.79e+10Hz 0.00675193 -0.00646252
+ 2.8e+10Hz 0.00674593 -0.00649093
+ 2.81e+10Hz 0.00673994 -0.00651933
+ 2.82e+10Hz 0.00673394 -0.00654773
+ 2.83e+10Hz 0.00672795 -0.00657611
+ 2.84e+10Hz 0.00672195 -0.00660449
+ 2.85e+10Hz 0.00671596 -0.00663286
+ 2.86e+10Hz 0.00670996 -0.00666123
+ 2.87e+10Hz 0.00670396 -0.0066896
+ 2.88e+10Hz 0.00669797 -0.00671798
+ 2.89e+10Hz 0.00669197 -0.00674635
+ 2.9e+10Hz 0.00668596 -0.00677473
+ 2.91e+10Hz 0.00667996 -0.00680312
+ 2.92e+10Hz 0.00667394 -0.00683151
+ 2.93e+10Hz 0.00666793 -0.00685991
+ 2.94e+10Hz 0.00666191 -0.00688833
+ 2.95e+10Hz 0.00665588 -0.00691675
+ 2.96e+10Hz 0.00664984 -0.00694519
+ 2.97e+10Hz 0.00664379 -0.00697364
+ 2.98e+10Hz 0.00663774 -0.00700211
+ 2.99e+10Hz 0.00663167 -0.00703059
+ 3e+10Hz 0.00662559 -0.0070591
+ 3.01e+10Hz 0.0066195 -0.00708762
+ 3.02e+10Hz 0.0066134 -0.00711617
+ 3.03e+10Hz 0.00660728 -0.00714473
+ 3.04e+10Hz 0.00660115 -0.00717332
+ 3.05e+10Hz 0.00659499 -0.00720193
+ 3.06e+10Hz 0.00658882 -0.00723057
+ 3.07e+10Hz 0.00658263 -0.00725924
+ 3.08e+10Hz 0.00657642 -0.00728793
+ 3.09e+10Hz 0.00657018 -0.00731664
+ 3.1e+10Hz 0.00656392 -0.00734539
+ 3.11e+10Hz 0.00655764 -0.00737417
+ 3.12e+10Hz 0.00655133 -0.00740297
+ 3.13e+10Hz 0.00654499 -0.00743181
+ 3.14e+10Hz 0.00653862 -0.00746067
+ 3.15e+10Hz 0.00653223 -0.00748957
+ 3.16e+10Hz 0.0065258 -0.00751851
+ 3.17e+10Hz 0.00651933 -0.00754747
+ 3.18e+10Hz 0.00651284 -0.00757647
+ 3.19e+10Hz 0.0065063 -0.0076055
+ 3.2e+10Hz 0.00649973 -0.00763456
+ 3.21e+10Hz 0.00649312 -0.00766366
+ 3.22e+10Hz 0.00648647 -0.0076928
+ 3.23e+10Hz 0.00647977 -0.00772197
+ 3.24e+10Hz 0.00647304 -0.00775117
+ 3.25e+10Hz 0.00646626 -0.00778041
+ 3.26e+10Hz 0.00645943 -0.00780968
+ 3.27e+10Hz 0.00645255 -0.00783899
+ 3.28e+10Hz 0.00644563 -0.00786834
+ 3.29e+10Hz 0.00643865 -0.00789772
+ 3.3e+10Hz 0.00643162 -0.00792713
+ 3.31e+10Hz 0.00642454 -0.00795658
+ 3.32e+10Hz 0.00641741 -0.00798607
+ 3.33e+10Hz 0.00641021 -0.00801559
+ 3.34e+10Hz 0.00640296 -0.00804514
+ 3.35e+10Hz 0.00639565 -0.00807473
+ 3.36e+10Hz 0.00638828 -0.00810435
+ 3.37e+10Hz 0.00638085 -0.00813401
+ 3.38e+10Hz 0.00637336 -0.0081637
+ 3.39e+10Hz 0.00636579 -0.00819342
+ 3.4e+10Hz 0.00635817 -0.00822317
+ 3.41e+10Hz 0.00635047 -0.00825296
+ 3.42e+10Hz 0.00634271 -0.00828277
+ 3.43e+10Hz 0.00633488 -0.00831262
+ 3.44e+10Hz 0.00632698 -0.00834249
+ 3.45e+10Hz 0.006319 -0.00837239
+ 3.46e+10Hz 0.00631095 -0.00840233
+ 3.47e+10Hz 0.00630283 -0.00843229
+ 3.48e+10Hz 0.00629463 -0.00846227
+ 3.49e+10Hz 0.00628635 -0.00849228
+ 3.5e+10Hz 0.006278 -0.00852232
+ 3.51e+10Hz 0.00626956 -0.00855238
+ 3.52e+10Hz 0.00626105 -0.00858247
+ 3.53e+10Hz 0.00625245 -0.00861258
+ 3.54e+10Hz 0.00624377 -0.0086427
+ 3.55e+10Hz 0.00623501 -0.00867285
+ 3.56e+10Hz 0.00622617 -0.00870302
+ 3.57e+10Hz 0.00621724 -0.00873321
+ 3.58e+10Hz 0.00620822 -0.00876341
+ 3.59e+10Hz 0.00619912 -0.00879363
+ 3.6e+10Hz 0.00618992 -0.00882387
+ 3.61e+10Hz 0.00618064 -0.00885412
+ 3.62e+10Hz 0.00617128 -0.00888438
+ 3.63e+10Hz 0.00616182 -0.00891465
+ 3.64e+10Hz 0.00615227 -0.00894494
+ 3.65e+10Hz 0.00614262 -0.00897523
+ 3.66e+10Hz 0.00613289 -0.00900553
+ 3.67e+10Hz 0.00612307 -0.00903584
+ 3.68e+10Hz 0.00611315 -0.00906616
+ 3.69e+10Hz 0.00610313 -0.00909648
+ 3.7e+10Hz 0.00609303 -0.0091268
+ 3.71e+10Hz 0.00608282 -0.00915712
+ 3.72e+10Hz 0.00607253 -0.00918745
+ 3.73e+10Hz 0.00606213 -0.00921777
+ 3.74e+10Hz 0.00605165 -0.00924809
+ 3.75e+10Hz 0.00604106 -0.00927841
+ 3.76e+10Hz 0.00603038 -0.00930872
+ 3.77e+10Hz 0.0060196 -0.00933903
+ 3.78e+10Hz 0.00600873 -0.00936933
+ 3.79e+10Hz 0.00599776 -0.00939962
+ 3.8e+10Hz 0.00598669 -0.0094299
+ 3.81e+10Hz 0.00597552 -0.00946017
+ 3.82e+10Hz 0.00596426 -0.00949043
+ 3.83e+10Hz 0.0059529 -0.00952067
+ 3.84e+10Hz 0.00594144 -0.0095509
+ 3.85e+10Hz 0.00592989 -0.00958111
+ 3.86e+10Hz 0.00591823 -0.00961131
+ 3.87e+10Hz 0.00590648 -0.00964148
+ 3.88e+10Hz 0.00589464 -0.00967163
+ 3.89e+10Hz 0.00588269 -0.00970177
+ 3.9e+10Hz 0.00587065 -0.00973187
+ 3.91e+10Hz 0.00585851 -0.00976196
+ 3.92e+10Hz 0.00584628 -0.00979201
+ 3.93e+10Hz 0.00583395 -0.00982204
+ 3.94e+10Hz 0.00582152 -0.00985205
+ 3.95e+10Hz 0.005809 -0.00988202
+ 3.96e+10Hz 0.00579639 -0.00991196
+ 3.97e+10Hz 0.00578368 -0.00994187
+ 3.98e+10Hz 0.00577088 -0.00997175
+ 3.99e+10Hz 0.00575798 -0.0100016
+ 4e+10Hz 0.00574499 -0.0100314
+ 4.01e+10Hz 0.00573191 -0.0100612
+ 4.02e+10Hz 0.00571873 -0.0100909
+ 4.03e+10Hz 0.00570547 -0.0101206
+ 4.04e+10Hz 0.00569211 -0.0101502
+ 4.05e+10Hz 0.00567866 -0.0101798
+ 4.06e+10Hz 0.00566513 -0.0102094
+ 4.07e+10Hz 0.0056515 -0.0102389
+ 4.08e+10Hz 0.00563779 -0.0102684
+ 4.09e+10Hz 0.00562399 -0.0102979
+ 4.1e+10Hz 0.00561011 -0.0103272
+ 4.11e+10Hz 0.00559614 -0.0103566
+ 4.12e+10Hz 0.00558208 -0.0103859
+ 4.13e+10Hz 0.00556794 -0.0104151
+ 4.14e+10Hz 0.00555372 -0.0104443
+ 4.15e+10Hz 0.00553941 -0.0104734
+ 4.16e+10Hz 0.00552503 -0.0105025
+ 4.17e+10Hz 0.00551056 -0.0105316
+ 4.18e+10Hz 0.00549601 -0.0105605
+ 4.19e+10Hz 0.00548139 -0.0105895
+ 4.2e+10Hz 0.00546669 -0.0106183
+ 4.21e+10Hz 0.00545191 -0.0106472
+ 4.22e+10Hz 0.00543705 -0.0106759
+ 4.23e+10Hz 0.00542212 -0.0107046
+ 4.24e+10Hz 0.00540712 -0.0107333
+ 4.25e+10Hz 0.00539205 -0.0107619
+ 4.26e+10Hz 0.0053769 -0.0107904
+ 4.27e+10Hz 0.00536168 -0.0108189
+ 4.28e+10Hz 0.0053464 -0.0108473
+ 4.29e+10Hz 0.00533104 -0.0108756
+ 4.3e+10Hz 0.00531562 -0.0109039
+ 4.31e+10Hz 0.00530013 -0.0109321
+ 4.32e+10Hz 0.00528458 -0.0109603
+ 4.33e+10Hz 0.00526896 -0.0109884
+ 4.34e+10Hz 0.00525328 -0.0110164
+ 4.35e+10Hz 0.00523754 -0.0110444
+ 4.36e+10Hz 0.00522174 -0.0110723
+ 4.37e+10Hz 0.00520587 -0.0111001
+ 4.38e+10Hz 0.00518995 -0.0111279
+ 4.39e+10Hz 0.00517397 -0.0111556
+ 4.4e+10Hz 0.00515794 -0.0111833
+ 4.41e+10Hz 0.00514185 -0.0112109
+ 4.42e+10Hz 0.0051257 -0.0112384
+ 4.43e+10Hz 0.00510951 -0.0112659
+ 4.44e+10Hz 0.00509326 -0.0112933
+ 4.45e+10Hz 0.00507696 -0.0113206
+ 4.46e+10Hz 0.00506061 -0.0113479
+ 4.47e+10Hz 0.00504421 -0.0113751
+ 4.48e+10Hz 0.00502776 -0.0114022
+ 4.49e+10Hz 0.00501127 -0.0114293
+ 4.5e+10Hz 0.00499473 -0.0114563
+ 4.51e+10Hz 0.00497815 -0.0114833
+ 4.52e+10Hz 0.00496152 -0.0115102
+ 4.53e+10Hz 0.00494485 -0.011537
+ 4.54e+10Hz 0.00492814 -0.0115637
+ 4.55e+10Hz 0.00491139 -0.0115904
+ 4.56e+10Hz 0.0048946 -0.0116171
+ 4.57e+10Hz 0.00487777 -0.0116436
+ 4.58e+10Hz 0.00486091 -0.0116701
+ 4.59e+10Hz 0.004844 -0.0116966
+ 4.6e+10Hz 0.00482706 -0.0117229
+ 4.61e+10Hz 0.00481009 -0.0117493
+ 4.62e+10Hz 0.00479308 -0.0117755
+ 4.63e+10Hz 0.00477604 -0.0118017
+ 4.64e+10Hz 0.00475897 -0.0118279
+ 4.65e+10Hz 0.00474187 -0.0118539
+ 4.66e+10Hz 0.00472473 -0.01188
+ 4.67e+10Hz 0.00470757 -0.0119059
+ 4.68e+10Hz 0.00469037 -0.0119318
+ 4.69e+10Hz 0.00467315 -0.0119577
+ 4.7e+10Hz 0.0046559 -0.0119834
+ 4.71e+10Hz 0.00463863 -0.0120092
+ 4.72e+10Hz 0.00462133 -0.0120349
+ 4.73e+10Hz 0.004604 -0.0120605
+ 4.74e+10Hz 0.00458665 -0.012086
+ 4.75e+10Hz 0.00456928 -0.0121115
+ 4.76e+10Hz 0.00455188 -0.012137
+ 4.77e+10Hz 0.00453446 -0.0121624
+ 4.78e+10Hz 0.00451701 -0.0121878
+ 4.79e+10Hz 0.00449955 -0.0122131
+ 4.8e+10Hz 0.00448206 -0.0122383
+ 4.81e+10Hz 0.00446456 -0.0122635
+ 4.82e+10Hz 0.00444703 -0.0122887
+ 4.83e+10Hz 0.00442948 -0.0123138
+ 4.84e+10Hz 0.00441192 -0.0123388
+ 4.85e+10Hz 0.00439433 -0.0123638
+ 4.86e+10Hz 0.00437673 -0.0123888
+ 4.87e+10Hz 0.00435911 -0.0124137
+ 4.88e+10Hz 0.00434147 -0.0124386
+ 4.89e+10Hz 0.00432381 -0.0124634
+ 4.9e+10Hz 0.00430614 -0.0124882
+ 4.91e+10Hz 0.00428845 -0.0125129
+ 4.92e+10Hz 0.00427074 -0.0125376
+ 4.93e+10Hz 0.00425302 -0.0125623
+ 4.94e+10Hz 0.00423528 -0.0125869
+ 4.95e+10Hz 0.00421752 -0.0126114
+ 4.96e+10Hz 0.00419975 -0.012636
+ 4.97e+10Hz 0.00418197 -0.0126605
+ 4.98e+10Hz 0.00416416 -0.0126849
+ 4.99e+10Hz 0.00414634 -0.0127094
+ 5e+10Hz 0.00412851 -0.0127337
+ 5.01e+10Hz 0.00411066 -0.0127581
+ 5.02e+10Hz 0.00409279 -0.0127824
+ 5.03e+10Hz 0.00407491 -0.0128067
+ 5.04e+10Hz 0.00405702 -0.0128309
+ 5.05e+10Hz 0.00403911 -0.0128552
+ 5.06e+10Hz 0.00402118 -0.0128793
+ 5.07e+10Hz 0.00400323 -0.0129035
+ 5.08e+10Hz 0.00398527 -0.0129276
+ 5.09e+10Hz 0.0039673 -0.0129517
+ 5.1e+10Hz 0.0039493 -0.0129758
+ 5.11e+10Hz 0.00393129 -0.0129998
+ 5.12e+10Hz 0.00391327 -0.0130238
+ 5.13e+10Hz 0.00389523 -0.0130478
+ 5.14e+10Hz 0.00387717 -0.0130718
+ 5.15e+10Hz 0.00385909 -0.0130957
+ 5.16e+10Hz 0.00384099 -0.0131196
+ 5.17e+10Hz 0.00382288 -0.0131435
+ 5.18e+10Hz 0.00380475 -0.0131673
+ 5.19e+10Hz 0.00378659 -0.0131912
+ 5.2e+10Hz 0.00376842 -0.013215
+ 5.21e+10Hz 0.00375023 -0.0132388
+ 5.22e+10Hz 0.00373202 -0.0132625
+ 5.23e+10Hz 0.00371379 -0.0132863
+ 5.24e+10Hz 0.00369554 -0.01331
+ 5.25e+10Hz 0.00367727 -0.0133337
+ 5.26e+10Hz 0.00365898 -0.0133574
+ 5.27e+10Hz 0.00364066 -0.013381
+ 5.28e+10Hz 0.00362232 -0.0134047
+ 5.29e+10Hz 0.00360396 -0.0134283
+ 5.3e+10Hz 0.00358558 -0.0134519
+ 5.31e+10Hz 0.00356717 -0.0134755
+ 5.32e+10Hz 0.00354873 -0.0134991
+ 5.33e+10Hz 0.00353027 -0.0135226
+ 5.34e+10Hz 0.00351179 -0.0135462
+ 5.35e+10Hz 0.00349328 -0.0135697
+ 5.36e+10Hz 0.00347474 -0.0135932
+ 5.37e+10Hz 0.00345617 -0.0136167
+ 5.38e+10Hz 0.00343758 -0.0136402
+ 5.39e+10Hz 0.00341896 -0.0136636
+ 5.4e+10Hz 0.00340031 -0.0136871
+ 5.41e+10Hz 0.00338162 -0.0137105
+ 5.42e+10Hz 0.00336291 -0.0137339
+ 5.43e+10Hz 0.00334417 -0.0137573
+ 5.44e+10Hz 0.0033254 -0.0137807
+ 5.45e+10Hz 0.00330659 -0.0138041
+ 5.46e+10Hz 0.00328775 -0.0138274
+ 5.47e+10Hz 0.00326888 -0.0138507
+ 5.48e+10Hz 0.00324997 -0.0138741
+ 5.49e+10Hz 0.00323103 -0.0138974
+ 5.5e+10Hz 0.00321206 -0.0139207
+ 5.51e+10Hz 0.00319305 -0.013944
+ 5.52e+10Hz 0.003174 -0.0139672
+ 5.53e+10Hz 0.00315491 -0.0139905
+ 5.54e+10Hz 0.00313579 -0.0140137
+ 5.55e+10Hz 0.00311663 -0.0140369
+ 5.56e+10Hz 0.00309743 -0.0140601
+ 5.57e+10Hz 0.00307819 -0.0140833
+ 5.58e+10Hz 0.00305891 -0.0141065
+ 5.59e+10Hz 0.00303959 -0.0141296
+ 5.6e+10Hz 0.00302023 -0.0141528
+ 5.61e+10Hz 0.00300083 -0.0141759
+ 5.62e+10Hz 0.00298138 -0.014199
+ 5.63e+10Hz 0.0029619 -0.0142221
+ 5.64e+10Hz 0.00294236 -0.0142452
+ 5.65e+10Hz 0.00292279 -0.0142682
+ 5.66e+10Hz 0.00290317 -0.0142913
+ 5.67e+10Hz 0.0028835 -0.0143143
+ 5.68e+10Hz 0.00286379 -0.0143373
+ 5.69e+10Hz 0.00284404 -0.0143603
+ 5.7e+10Hz 0.00282424 -0.0143832
+ 5.71e+10Hz 0.00280439 -0.0144062
+ 5.72e+10Hz 0.00278449 -0.0144291
+ 5.73e+10Hz 0.00276454 -0.014452
+ 5.74e+10Hz 0.00274455 -0.0144749
+ 5.75e+10Hz 0.00272451 -0.0144978
+ 5.76e+10Hz 0.00270442 -0.0145206
+ 5.77e+10Hz 0.00268427 -0.0145434
+ 5.78e+10Hz 0.00266408 -0.0145662
+ 5.79e+10Hz 0.00264384 -0.014589
+ 5.8e+10Hz 0.00262355 -0.0146117
+ 5.81e+10Hz 0.0026032 -0.0146345
+ 5.82e+10Hz 0.00258281 -0.0146571
+ 5.83e+10Hz 0.00256236 -0.0146798
+ 5.84e+10Hz 0.00254186 -0.0147025
+ 5.85e+10Hz 0.00252131 -0.0147251
+ 5.86e+10Hz 0.00250071 -0.0147477
+ 5.87e+10Hz 0.00248005 -0.0147702
+ 5.88e+10Hz 0.00245934 -0.0147928
+ 5.89e+10Hz 0.00243858 -0.0148153
+ 5.9e+10Hz 0.00241776 -0.0148378
+ 5.91e+10Hz 0.00239689 -0.0148602
+ 5.92e+10Hz 0.00237597 -0.0148826
+ 5.93e+10Hz 0.00235499 -0.014905
+ 5.94e+10Hz 0.00233395 -0.0149274
+ 5.95e+10Hz 0.00231287 -0.0149497
+ 5.96e+10Hz 0.00229172 -0.014972
+ 5.97e+10Hz 0.00227053 -0.0149942
+ 5.98e+10Hz 0.00224928 -0.0150164
+ 5.99e+10Hz 0.00222797 -0.0150386
+ 6e+10Hz 0.00220661 -0.0150607
+ 6.01e+10Hz 0.0021852 -0.0150829
+ 6.02e+10Hz 0.00216373 -0.0151049
+ 6.03e+10Hz 0.0021422 -0.015127
+ 6.04e+10Hz 0.00212063 -0.0151489
+ 6.05e+10Hz 0.00209899 -0.0151709
+ 6.06e+10Hz 0.00207731 -0.0151928
+ 6.07e+10Hz 0.00205556 -0.0152147
+ 6.08e+10Hz 0.00203377 -0.0152365
+ 6.09e+10Hz 0.00201192 -0.0152583
+ 6.1e+10Hz 0.00199002 -0.01528
+ 6.11e+10Hz 0.00196806 -0.0153017
+ 6.12e+10Hz 0.00194605 -0.0153234
+ 6.13e+10Hz 0.00192398 -0.015345
+ 6.14e+10Hz 0.00190187 -0.0153665
+ 6.15e+10Hz 0.0018797 -0.015388
+ 6.16e+10Hz 0.00185747 -0.0154095
+ 6.17e+10Hz 0.0018352 -0.0154309
+ 6.18e+10Hz 0.00181287 -0.0154523
+ 6.19e+10Hz 0.00179049 -0.0154736
+ 6.2e+10Hz 0.00176806 -0.0154949
+ 6.21e+10Hz 0.00174558 -0.0155161
+ 6.22e+10Hz 0.00172305 -0.0155373
+ 6.23e+10Hz 0.00170047 -0.0155584
+ 6.24e+10Hz 0.00167783 -0.0155795
+ 6.25e+10Hz 0.00165515 -0.0156005
+ 6.26e+10Hz 0.00163242 -0.0156214
+ 6.27e+10Hz 0.00160964 -0.0156423
+ 6.28e+10Hz 0.00158682 -0.0156632
+ 6.29e+10Hz 0.00156394 -0.015684
+ 6.3e+10Hz 0.00154102 -0.0157047
+ 6.31e+10Hz 0.00151805 -0.0157254
+ 6.32e+10Hz 0.00149503 -0.015746
+ 6.33e+10Hz 0.00147197 -0.0157666
+ 6.34e+10Hz 0.00144886 -0.0157871
+ 6.35e+10Hz 0.00142571 -0.0158076
+ 6.36e+10Hz 0.00140252 -0.015828
+ 6.37e+10Hz 0.00137928 -0.0158483
+ 6.38e+10Hz 0.001356 -0.0158686
+ 6.39e+10Hz 0.00133267 -0.0158888
+ 6.4e+10Hz 0.0013093 -0.015909
+ 6.41e+10Hz 0.0012859 -0.0159291
+ 6.42e+10Hz 0.00126245 -0.0159491
+ 6.43e+10Hz 0.00123896 -0.0159691
+ 6.44e+10Hz 0.00121543 -0.015989
+ 6.45e+10Hz 0.00119186 -0.0160089
+ 6.46e+10Hz 0.00116826 -0.0160287
+ 6.47e+10Hz 0.00114461 -0.0160484
+ 6.48e+10Hz 0.00112093 -0.016068
+ 6.49e+10Hz 0.00109722 -0.0160876
+ 6.5e+10Hz 0.00107346 -0.0161072
+ 6.51e+10Hz 0.00104968 -0.0161267
+ 6.52e+10Hz 0.00102586 -0.0161461
+ 6.53e+10Hz 0.001002 -0.0161654
+ 6.54e+10Hz 0.000978114 -0.0161847
+ 6.55e+10Hz 0.000954194 -0.0162039
+ 6.56e+10Hz 0.000930242 -0.0162231
+ 6.57e+10Hz 0.000906259 -0.0162422
+ 6.58e+10Hz 0.000882246 -0.0162612
+ 6.59e+10Hz 0.000858204 -0.0162802
+ 6.6e+10Hz 0.000834133 -0.0162991
+ 6.61e+10Hz 0.000810033 -0.0163179
+ 6.62e+10Hz 0.000785906 -0.0163367
+ 6.63e+10Hz 0.000761752 -0.0163554
+ 6.64e+10Hz 0.000737572 -0.016374
+ 6.65e+10Hz 0.000713366 -0.0163926
+ 6.66e+10Hz 0.000689136 -0.0164111
+ 6.67e+10Hz 0.000664881 -0.0164295
+ 6.68e+10Hz 0.000640603 -0.0164479
+ 6.69e+10Hz 0.000616302 -0.0164662
+ 6.7e+10Hz 0.000591979 -0.0164845
+ 6.71e+10Hz 0.000567634 -0.0165026
+ 6.72e+10Hz 0.000543269 -0.0165208
+ 6.73e+10Hz 0.000518883 -0.0165388
+ 6.74e+10Hz 0.000494478 -0.0165568
+ 6.75e+10Hz 0.000470054 -0.0165747
+ 6.76e+10Hz 0.000445611 -0.0165926
+ 6.77e+10Hz 0.000421151 -0.0166104
+ 6.78e+10Hz 0.000396674 -0.0166281
+ 6.79e+10Hz 0.00037218 -0.0166458
+ 6.8e+10Hz 0.00034767 -0.0166634
+ 6.81e+10Hz 0.000323145 -0.016681
+ 6.82e+10Hz 0.000298606 -0.0166985
+ 6.83e+10Hz 0.000274052 -0.0167159
+ 6.84e+10Hz 0.000249484 -0.0167332
+ 6.85e+10Hz 0.000224904 -0.0167505
+ 6.86e+10Hz 0.00020031 -0.0167678
+ 6.87e+10Hz 0.000175705 -0.016785
+ 6.88e+10Hz 0.000151089 -0.0168021
+ 6.89e+10Hz 0.000126461 -0.0168191
+ 6.9e+10Hz 0.000101823 -0.0168361
+ 6.91e+10Hz 7.71752e-05 -0.0168531
+ 6.92e+10Hz 5.25176e-05 -0.01687
+ 6.93e+10Hz 2.7851e-05 -0.0168868
+ 6.94e+10Hz 3.17567e-06 -0.0169035
+ 6.95e+10Hz -2.15078e-05 -0.0169202
+ 6.96e+10Hz -4.61991e-05 -0.0169369
+ 6.97e+10Hz -7.08978e-05 -0.0169535
+ 6.98e+10Hz -9.56035e-05 -0.01697
+ 6.99e+10Hz -0.000120316 -0.0169865
+ 7e+10Hz -0.000145034 -0.0170029
+ 7.01e+10Hz -0.000169759 -0.0170193
+ 7.02e+10Hz -0.000194489 -0.0170356
+ 7.03e+10Hz -0.000219224 -0.0170519
+ 7.04e+10Hz -0.000243964 -0.0170681
+ 7.05e+10Hz -0.000268709 -0.0170842
+ 7.06e+10Hz -0.000293458 -0.0171003
+ 7.07e+10Hz -0.000318212 -0.0171163
+ 7.08e+10Hz -0.000342969 -0.0171323
+ 7.09e+10Hz -0.00036773 -0.0171483
+ 7.1e+10Hz -0.000392494 -0.0171642
+ 7.11e+10Hz -0.000417262 -0.01718
+ 7.12e+10Hz -0.000442032 -0.0171958
+ 7.13e+10Hz -0.000466806 -0.0172116
+ 7.14e+10Hz -0.000491582 -0.0172272
+ 7.15e+10Hz -0.000516361 -0.0172429
+ 7.16e+10Hz -0.000541142 -0.0172585
+ 7.17e+10Hz -0.000565925 -0.017274
+ 7.18e+10Hz -0.000590711 -0.0172895
+ 7.19e+10Hz -0.000615499 -0.017305
+ 7.2e+10Hz -0.000640289 -0.0173204
+ 7.21e+10Hz -0.000665081 -0.0173358
+ 7.22e+10Hz -0.000689875 -0.0173511
+ 7.23e+10Hz -0.000714671 -0.0173664
+ 7.24e+10Hz -0.000739469 -0.0173816
+ 7.25e+10Hz -0.000764269 -0.0173968
+ 7.26e+10Hz -0.000789071 -0.0174119
+ 7.27e+10Hz -0.000813875 -0.017427
+ 7.28e+10Hz -0.000838681 -0.0174421
+ 7.29e+10Hz -0.00086349 -0.0174571
+ 7.3e+10Hz -0.0008883 -0.0174721
+ 7.31e+10Hz -0.000913113 -0.017487
+ 7.32e+10Hz -0.000937929 -0.0175019
+ 7.33e+10Hz -0.000962747 -0.0175168
+ 7.34e+10Hz -0.000987567 -0.0175316
+ 7.35e+10Hz -0.00101239 -0.0175464
+ 7.36e+10Hz -0.00103722 -0.0175611
+ 7.37e+10Hz -0.00106205 -0.0175758
+ 7.38e+10Hz -0.00108688 -0.0175905
+ 7.39e+10Hz -0.00111172 -0.0176051
+ 7.4e+10Hz -0.00113656 -0.0176197
+ 7.41e+10Hz -0.0011614 -0.0176343
+ 7.42e+10Hz -0.00118625 -0.0176488
+ 7.43e+10Hz -0.0012111 -0.0176633
+ 7.44e+10Hz -0.00123596 -0.0176778
+ 7.45e+10Hz -0.00126082 -0.0176922
+ 7.46e+10Hz -0.00128569 -0.0177066
+ 7.47e+10Hz -0.00131056 -0.0177209
+ 7.48e+10Hz -0.00133544 -0.0177352
+ 7.49e+10Hz -0.00136033 -0.0177495
+ 7.5e+10Hz -0.00138522 -0.0177638
+ 7.51e+10Hz -0.00141012 -0.017778
+ 7.52e+10Hz -0.00143503 -0.0177921
+ 7.53e+10Hz -0.00145994 -0.0178063
+ 7.54e+10Hz -0.00148486 -0.0178204
+ 7.55e+10Hz -0.00150979 -0.0178345
+ 7.56e+10Hz -0.00153472 -0.0178486
+ 7.57e+10Hz -0.00155967 -0.0178626
+ 7.58e+10Hz -0.00158463 -0.0178766
+ 7.59e+10Hz -0.00160959 -0.0178905
+ 7.6e+10Hz -0.00163456 -0.0179045
+ 7.61e+10Hz -0.00165955 -0.0179184
+ 7.62e+10Hz -0.00168454 -0.0179322
+ 7.63e+10Hz -0.00170955 -0.0179461
+ 7.64e+10Hz -0.00173457 -0.0179599
+ 7.65e+10Hz -0.0017596 -0.0179737
+ 7.66e+10Hz -0.00178464 -0.0179874
+ 7.67e+10Hz -0.00180969 -0.0180011
+ 7.68e+10Hz -0.00183476 -0.0180148
+ 7.69e+10Hz -0.00185984 -0.0180285
+ 7.7e+10Hz -0.00188493 -0.0180421
+ 7.71e+10Hz -0.00191004 -0.0180557
+ 7.72e+10Hz -0.00193516 -0.0180693
+ 7.73e+10Hz -0.0019603 -0.0180828
+ 7.74e+10Hz -0.00198546 -0.0180963
+ 7.75e+10Hz -0.00201062 -0.0181098
+ 7.76e+10Hz -0.00203581 -0.0181232
+ 7.77e+10Hz -0.00206101 -0.0181366
+ 7.78e+10Hz -0.00208623 -0.01815
+ 7.79e+10Hz -0.00211147 -0.0181634
+ 7.8e+10Hz -0.00213672 -0.0181767
+ 7.81e+10Hz -0.00216199 -0.01819
+ 7.82e+10Hz -0.00218728 -0.0182033
+ 7.83e+10Hz -0.00221259 -0.0182165
+ 7.84e+10Hz -0.00223792 -0.0182297
+ 7.85e+10Hz -0.00226327 -0.0182429
+ 7.86e+10Hz -0.00228864 -0.018256
+ 7.87e+10Hz -0.00231403 -0.0182691
+ 7.88e+10Hz -0.00233944 -0.0182822
+ 7.89e+10Hz -0.00236487 -0.0182952
+ 7.9e+10Hz -0.00239032 -0.0183083
+ 7.91e+10Hz -0.0024158 -0.0183212
+ 7.92e+10Hz -0.00244129 -0.0183342
+ 7.93e+10Hz -0.00246681 -0.0183471
+ 7.94e+10Hz -0.00249235 -0.01836
+ 7.95e+10Hz -0.00251792 -0.0183728
+ 7.96e+10Hz -0.00254351 -0.0183856
+ 7.97e+10Hz -0.00256912 -0.0183984
+ 7.98e+10Hz -0.00259475 -0.0184112
+ 7.99e+10Hz -0.00262041 -0.0184239
+ 8e+10Hz -0.0026461 -0.0184366
+ 8.01e+10Hz -0.00267181 -0.0184492
+ 8.02e+10Hz -0.00269754 -0.0184618
+ 8.03e+10Hz -0.0027233 -0.0184744
+ 8.04e+10Hz -0.00274908 -0.0184869
+ 8.05e+10Hz -0.00277489 -0.0184994
+ 8.06e+10Hz -0.00280073 -0.0185119
+ 8.07e+10Hz -0.00282659 -0.0185243
+ 8.08e+10Hz -0.00285248 -0.0185367
+ 8.09e+10Hz -0.0028784 -0.018549
+ 8.1e+10Hz -0.00290434 -0.0185613
+ 8.11e+10Hz -0.00293031 -0.0185736
+ 8.12e+10Hz -0.0029563 -0.0185858
+ 8.13e+10Hz -0.00298233 -0.018598
+ 8.14e+10Hz -0.00300838 -0.0186101
+ 8.15e+10Hz -0.00303445 -0.0186222
+ 8.16e+10Hz -0.00306056 -0.0186343
+ 8.17e+10Hz -0.00308669 -0.0186463
+ 8.18e+10Hz -0.00311285 -0.0186583
+ 8.19e+10Hz -0.00313904 -0.0186702
+ 8.2e+10Hz -0.00316525 -0.0186821
+ 8.21e+10Hz -0.00319149 -0.018694
+ 8.22e+10Hz -0.00321776 -0.0187058
+ 8.23e+10Hz -0.00324406 -0.0187175
+ 8.24e+10Hz -0.00327039 -0.0187293
+ 8.25e+10Hz -0.00329674 -0.0187409
+ 8.26e+10Hz -0.00332312 -0.0187525
+ 8.27e+10Hz -0.00334953 -0.0187641
+ 8.28e+10Hz -0.00337596 -0.0187756
+ 8.29e+10Hz -0.00340242 -0.0187871
+ 8.3e+10Hz -0.00342892 -0.0187986
+ 8.31e+10Hz -0.00345543 -0.0188099
+ 8.32e+10Hz -0.00348198 -0.0188213
+ 8.33e+10Hz -0.00350855 -0.0188326
+ 8.34e+10Hz -0.00353515 -0.0188438
+ 8.35e+10Hz -0.00356177 -0.018855
+ 8.36e+10Hz -0.00358843 -0.0188661
+ 8.37e+10Hz -0.0036151 -0.0188772
+ 8.38e+10Hz -0.00364181 -0.0188882
+ 8.39e+10Hz -0.00366854 -0.0188992
+ 8.4e+10Hz -0.0036953 -0.0189101
+ 8.41e+10Hz -0.00372208 -0.018921
+ 8.42e+10Hz -0.00374888 -0.0189318
+ 8.43e+10Hz -0.00377572 -0.0189426
+ 8.44e+10Hz -0.00380258 -0.0189533
+ 8.45e+10Hz -0.00382946 -0.0189639
+ 8.46e+10Hz -0.00385636 -0.0189745
+ 8.47e+10Hz -0.00388329 -0.0189851
+ 8.48e+10Hz -0.00391025 -0.0189956
+ 8.49e+10Hz -0.00393723 -0.019006
+ 8.5e+10Hz -0.00396423 -0.0190164
+ 8.51e+10Hz -0.00399125 -0.0190267
+ 8.52e+10Hz -0.0040183 -0.0190369
+ 8.53e+10Hz -0.00404537 -0.0190471
+ 8.54e+10Hz -0.00407246 -0.0190573
+ 8.55e+10Hz -0.00409957 -0.0190674
+ 8.56e+10Hz -0.0041267 -0.0190774
+ 8.57e+10Hz -0.00415385 -0.0190873
+ 8.58e+10Hz -0.00418103 -0.0190972
+ 8.59e+10Hz -0.00420822 -0.0191071
+ 8.6e+10Hz -0.00423543 -0.0191168
+ 8.61e+10Hz -0.00426266 -0.0191266
+ 8.62e+10Hz -0.00428991 -0.0191362
+ 8.63e+10Hz -0.00431718 -0.0191458
+ 8.64e+10Hz -0.00434447 -0.0191554
+ 8.65e+10Hz -0.00437177 -0.0191648
+ 8.66e+10Hz -0.00439909 -0.0191742
+ 8.67e+10Hz -0.00442643 -0.0191836
+ 8.68e+10Hz -0.00445378 -0.0191929
+ 8.69e+10Hz -0.00448115 -0.0192021
+ 8.7e+10Hz -0.00450853 -0.0192112
+ 8.71e+10Hz -0.00453593 -0.0192203
+ 8.72e+10Hz -0.00456334 -0.0192293
+ 8.73e+10Hz -0.00459076 -0.0192383
+ 8.74e+10Hz -0.0046182 -0.0192472
+ 8.75e+10Hz -0.00464565 -0.019256
+ 8.76e+10Hz -0.00467311 -0.0192648
+ 8.77e+10Hz -0.00470059 -0.0192735
+ 8.78e+10Hz -0.00472807 -0.0192822
+ 8.79e+10Hz -0.00475556 -0.0192907
+ 8.8e+10Hz -0.00478307 -0.0192992
+ 8.81e+10Hz -0.00481058 -0.0193077
+ 8.82e+10Hz -0.00483811 -0.0193161
+ 8.83e+10Hz -0.00486564 -0.0193244
+ 8.84e+10Hz -0.00489318 -0.0193326
+ 8.85e+10Hz -0.00492072 -0.0193408
+ 8.86e+10Hz -0.00494828 -0.0193489
+ 8.87e+10Hz -0.00497583 -0.019357
+ 8.88e+10Hz -0.0050034 -0.0193649
+ 8.89e+10Hz -0.00503097 -0.0193729
+ 8.9e+10Hz -0.00505855 -0.0193807
+ 8.91e+10Hz -0.00508613 -0.0193885
+ 8.92e+10Hz -0.00511371 -0.0193962
+ 8.93e+10Hz -0.0051413 -0.0194039
+ 8.94e+10Hz -0.00516888 -0.0194115
+ 8.95e+10Hz -0.00519648 -0.019419
+ 8.96e+10Hz -0.00522407 -0.0194265
+ 8.97e+10Hz -0.00525166 -0.0194338
+ 8.98e+10Hz -0.00527926 -0.0194412
+ 8.99e+10Hz -0.00530685 -0.0194484
+ 9e+10Hz -0.00533445 -0.0194556
+ 9.01e+10Hz -0.00536204 -0.0194628
+ 9.02e+10Hz -0.00538963 -0.0194698
+ 9.03e+10Hz -0.00541723 -0.0194768
+ 9.04e+10Hz -0.00544481 -0.0194838
+ 9.05e+10Hz -0.0054724 -0.0194907
+ 9.06e+10Hz -0.00549998 -0.0194975
+ 9.07e+10Hz -0.00552756 -0.0195042
+ 9.08e+10Hz -0.00555514 -0.0195109
+ 9.09e+10Hz -0.00558271 -0.0195175
+ 9.1e+10Hz -0.00561028 -0.0195241
+ 9.11e+10Hz -0.00563784 -0.0195306
+ 9.12e+10Hz -0.00566539 -0.019537
+ 9.13e+10Hz -0.00569294 -0.0195433
+ 9.14e+10Hz -0.00572048 -0.0195497
+ 9.15e+10Hz -0.00574802 -0.0195559
+ 9.16e+10Hz -0.00577554 -0.0195621
+ 9.17e+10Hz -0.00580306 -0.0195682
+ 9.18e+10Hz -0.00583058 -0.0195742
+ 9.19e+10Hz -0.00585808 -0.0195802
+ 9.2e+10Hz -0.00588557 -0.0195862
+ 9.21e+10Hz -0.00591306 -0.019592
+ 9.22e+10Hz -0.00594053 -0.0195979
+ 9.23e+10Hz -0.005968 -0.0196036
+ 9.24e+10Hz -0.00599545 -0.0196093
+ 9.25e+10Hz -0.0060229 -0.0196149
+ 9.26e+10Hz -0.00605033 -0.0196205
+ 9.27e+10Hz -0.00607776 -0.019626
+ 9.28e+10Hz -0.00610517 -0.0196315
+ 9.29e+10Hz -0.00613257 -0.0196369
+ 9.3e+10Hz -0.00615996 -0.0196422
+ 9.31e+10Hz -0.00618733 -0.0196475
+ 9.32e+10Hz -0.0062147 -0.0196527
+ 9.33e+10Hz -0.00624205 -0.0196579
+ 9.34e+10Hz -0.00626938 -0.019663
+ 9.35e+10Hz -0.00629671 -0.0196681
+ 9.36e+10Hz -0.00632402 -0.0196731
+ 9.37e+10Hz -0.00635132 -0.019678
+ 9.38e+10Hz -0.0063786 -0.0196829
+ 9.39e+10Hz -0.00640587 -0.0196877
+ 9.4e+10Hz -0.00643313 -0.0196925
+ 9.41e+10Hz -0.00646037 -0.0196972
+ 9.42e+10Hz -0.0064876 -0.0197019
+ 9.43e+10Hz -0.00651481 -0.0197065
+ 9.44e+10Hz -0.00654201 -0.0197111
+ 9.45e+10Hz -0.00656919 -0.0197156
+ 9.46e+10Hz -0.00659636 -0.0197201
+ 9.47e+10Hz -0.00662351 -0.0197245
+ 9.48e+10Hz -0.00665065 -0.0197288
+ 9.49e+10Hz -0.00667778 -0.0197331
+ 9.5e+10Hz -0.00670488 -0.0197374
+ 9.51e+10Hz -0.00673198 -0.0197416
+ 9.52e+10Hz -0.00675905 -0.0197457
+ 9.53e+10Hz -0.00678612 -0.0197499
+ 9.54e+10Hz -0.00681316 -0.0197539
+ 9.55e+10Hz -0.0068402 -0.0197579
+ 9.56e+10Hz -0.00686721 -0.0197619
+ 9.57e+10Hz -0.00689421 -0.0197658
+ 9.58e+10Hz -0.0069212 -0.0197696
+ 9.59e+10Hz -0.00694817 -0.0197734
+ 9.6e+10Hz -0.00697512 -0.0197772
+ 9.61e+10Hz -0.00700206 -0.0197809
+ 9.62e+10Hz -0.00702899 -0.0197846
+ 9.63e+10Hz -0.00705589 -0.0197882
+ 9.64e+10Hz -0.00708279 -0.0197918
+ 9.65e+10Hz -0.00710967 -0.0197953
+ 9.66e+10Hz -0.00713653 -0.0197988
+ 9.67e+10Hz -0.00716338 -0.0198023
+ 9.68e+10Hz -0.00719021 -0.0198056
+ 9.69e+10Hz -0.00721703 -0.019809
+ 9.7e+10Hz -0.00724383 -0.0198123
+ 9.71e+10Hz -0.00727062 -0.0198156
+ 9.72e+10Hz -0.0072974 -0.0198188
+ 9.73e+10Hz -0.00732416 -0.0198219
+ 9.74e+10Hz -0.0073509 -0.0198251
+ 9.75e+10Hz -0.00737763 -0.0198281
+ 9.76e+10Hz -0.00740435 -0.0198312
+ 9.77e+10Hz -0.00743105 -0.0198342
+ 9.78e+10Hz -0.00745774 -0.0198371
+ 9.79e+10Hz -0.00748442 -0.01984
+ 9.8e+10Hz -0.00751108 -0.0198429
+ 9.81e+10Hz -0.00753773 -0.0198457
+ 9.82e+10Hz -0.00756437 -0.0198485
+ 9.83e+10Hz -0.00759099 -0.0198513
+ 9.84e+10Hz -0.0076176 -0.0198539
+ 9.85e+10Hz -0.0076442 -0.0198566
+ 9.86e+10Hz -0.00767078 -0.0198592
+ 9.87e+10Hz -0.00769736 -0.0198618
+ 9.88e+10Hz -0.00772392 -0.0198643
+ 9.89e+10Hz -0.00775047 -0.0198668
+ 9.9e+10Hz -0.007777 -0.0198693
+ 9.91e+10Hz -0.00780353 -0.0198717
+ 9.92e+10Hz -0.00783004 -0.019874
+ 9.93e+10Hz -0.00785654 -0.0198763
+ 9.94e+10Hz -0.00788303 -0.0198786
+ 9.95e+10Hz -0.00790951 -0.0198809
+ 9.96e+10Hz -0.00793598 -0.0198831
+ 9.97e+10Hz -0.00796244 -0.0198852
+ 9.98e+10Hz -0.00798889 -0.0198873
+ 9.99e+10Hz -0.00801533 -0.0198894
+ 1e+11Hz -0.00804175 -0.0198914
+ 1.001e+11Hz -0.00806817 -0.0198934
+ 1.002e+11Hz -0.00809458 -0.0198954
+ 1.003e+11Hz -0.00812098 -0.0198973
+ 1.004e+11Hz -0.00814737 -0.0198992
+ 1.005e+11Hz -0.00817375 -0.019901
+ 1.006e+11Hz -0.00820012 -0.0199028
+ 1.007e+11Hz -0.00822648 -0.0199045
+ 1.008e+11Hz -0.00825283 -0.0199063
+ 1.009e+11Hz -0.00827917 -0.0199079
+ 1.01e+11Hz -0.00830551 -0.0199095
+ 1.011e+11Hz -0.00833184 -0.0199111
+ 1.012e+11Hz -0.00835816 -0.0199127
+ 1.013e+11Hz -0.00838447 -0.0199142
+ 1.014e+11Hz -0.00841077 -0.0199156
+ 1.015e+11Hz -0.00843707 -0.019917
+ 1.016e+11Hz -0.00846336 -0.0199184
+ 1.017e+11Hz -0.00848964 -0.0199197
+ 1.018e+11Hz -0.00851591 -0.019921
+ 1.019e+11Hz -0.00854217 -0.0199223
+ 1.02e+11Hz -0.00856843 -0.0199235
+ 1.021e+11Hz -0.00859468 -0.0199246
+ 1.022e+11Hz -0.00862093 -0.0199257
+ 1.023e+11Hz -0.00864717 -0.0199268
+ 1.024e+11Hz -0.0086734 -0.0199278
+ 1.025e+11Hz -0.00869962 -0.0199288
+ 1.026e+11Hz -0.00872584 -0.0199298
+ 1.027e+11Hz -0.00875205 -0.0199307
+ 1.028e+11Hz -0.00877825 -0.0199315
+ 1.029e+11Hz -0.00880445 -0.0199323
+ 1.03e+11Hz -0.00883064 -0.0199331
+ 1.031e+11Hz -0.00885682 -0.0199338
+ 1.032e+11Hz -0.008883 -0.0199345
+ 1.033e+11Hz -0.00890917 -0.0199351
+ 1.034e+11Hz -0.00893534 -0.0199357
+ 1.035e+11Hz -0.00896149 -0.0199363
+ 1.036e+11Hz -0.00898764 -0.0199368
+ 1.037e+11Hz -0.00901379 -0.0199372
+ 1.038e+11Hz -0.00903993 -0.0199376
+ 1.039e+11Hz -0.00906606 -0.019938
+ 1.04e+11Hz -0.00909218 -0.0199383
+ 1.041e+11Hz -0.0091183 -0.0199385
+ 1.042e+11Hz -0.00914441 -0.0199388
+ 1.043e+11Hz -0.00917052 -0.0199389
+ 1.044e+11Hz -0.00919662 -0.019939
+ 1.045e+11Hz -0.00922271 -0.0199391
+ 1.046e+11Hz -0.00924879 -0.0199391
+ 1.047e+11Hz -0.00927487 -0.0199391
+ 1.048e+11Hz -0.00930094 -0.019939
+ 1.049e+11Hz -0.009327 -0.0199389
+ 1.05e+11Hz -0.00935305 -0.0199388
+ 1.051e+11Hz -0.0093791 -0.0199385
+ 1.052e+11Hz -0.00940514 -0.0199383
+ 1.053e+11Hz -0.00943117 -0.019938
+ 1.054e+11Hz -0.00945719 -0.0199376
+ 1.055e+11Hz -0.00948321 -0.0199372
+ 1.056e+11Hz -0.00950921 -0.0199367
+ 1.057e+11Hz -0.00953521 -0.0199362
+ 1.058e+11Hz -0.0095612 -0.0199356
+ 1.059e+11Hz -0.00958718 -0.019935
+ 1.06e+11Hz -0.00961315 -0.0199343
+ 1.061e+11Hz -0.00963911 -0.0199336
+ 1.062e+11Hz -0.00966506 -0.0199328
+ 1.063e+11Hz -0.009691 -0.019932
+ 1.064e+11Hz -0.00971693 -0.0199311
+ 1.065e+11Hz -0.00974285 -0.0199302
+ 1.066e+11Hz -0.00976876 -0.0199292
+ 1.067e+11Hz -0.00979465 -0.0199281
+ 1.068e+11Hz -0.00982054 -0.019927
+ 1.069e+11Hz -0.00984641 -0.0199259
+ 1.07e+11Hz -0.00987228 -0.0199247
+ 1.071e+11Hz -0.00989813 -0.0199234
+ 1.072e+11Hz -0.00992397 -0.0199221
+ 1.073e+11Hz -0.00994979 -0.0199208
+ 1.074e+11Hz -0.0099756 -0.0199194
+ 1.075e+11Hz -0.0100014 -0.0199179
+ 1.076e+11Hz -0.0100272 -0.0199164
+ 1.077e+11Hz -0.010053 -0.0199148
+ 1.078e+11Hz -0.0100787 -0.0199132
+ 1.079e+11Hz -0.0101045 -0.0199115
+ 1.08e+11Hz -0.0101302 -0.0199097
+ 1.081e+11Hz -0.0101559 -0.0199079
+ 1.082e+11Hz -0.0101816 -0.0199061
+ 1.083e+11Hz -0.0102073 -0.0199042
+ 1.084e+11Hz -0.0102329 -0.0199022
+ 1.085e+11Hz -0.0102586 -0.0199002
+ 1.086e+11Hz -0.0102842 -0.0198981
+ 1.087e+11Hz -0.0103098 -0.019896
+ 1.088e+11Hz -0.0103354 -0.0198938
+ 1.089e+11Hz -0.010361 -0.0198916
+ 1.09e+11Hz -0.0103865 -0.0198893
+ 1.091e+11Hz -0.0104121 -0.0198869
+ 1.092e+11Hz -0.0104376 -0.0198845
+ 1.093e+11Hz -0.0104631 -0.0198821
+ 1.094e+11Hz -0.0104886 -0.0198796
+ 1.095e+11Hz -0.010514 -0.019877
+ 1.096e+11Hz -0.0105394 -0.0198744
+ 1.097e+11Hz -0.0105648 -0.0198717
+ 1.098e+11Hz -0.0105902 -0.0198689
+ 1.099e+11Hz -0.0106156 -0.0198661
+ 1.1e+11Hz -0.0106409 -0.0198633
+ 1.101e+11Hz -0.0106663 -0.0198604
+ 1.102e+11Hz -0.0106916 -0.0198574
+ 1.103e+11Hz -0.0107168 -0.0198544
+ 1.104e+11Hz -0.0107421 -0.0198513
+ 1.105e+11Hz -0.0107673 -0.0198482
+ 1.106e+11Hz -0.0107925 -0.019845
+ 1.107e+11Hz -0.0108177 -0.0198418
+ 1.108e+11Hz -0.0108428 -0.0198385
+ 1.109e+11Hz -0.0108679 -0.0198351
+ 1.11e+11Hz -0.010893 -0.0198317
+ 1.111e+11Hz -0.0109181 -0.0198283
+ 1.112e+11Hz -0.0109431 -0.0198248
+ 1.113e+11Hz -0.0109681 -0.0198212
+ 1.114e+11Hz -0.0109931 -0.0198176
+ 1.115e+11Hz -0.0110181 -0.0198139
+ 1.116e+11Hz -0.011043 -0.0198102
+ 1.117e+11Hz -0.0110679 -0.0198064
+ 1.118e+11Hz -0.0110927 -0.0198026
+ 1.119e+11Hz -0.0111176 -0.0197987
+ 1.12e+11Hz -0.0111424 -0.0197947
+ 1.121e+11Hz -0.0111671 -0.0197908
+ 1.122e+11Hz -0.0111919 -0.0197867
+ 1.123e+11Hz -0.0112166 -0.0197826
+ 1.124e+11Hz -0.0112412 -0.0197785
+ 1.125e+11Hz -0.0112659 -0.0197743
+ 1.126e+11Hz -0.0112905 -0.01977
+ 1.127e+11Hz -0.011315 -0.0197657
+ 1.128e+11Hz -0.0113396 -0.0197614
+ 1.129e+11Hz -0.0113641 -0.019757
+ 1.13e+11Hz -0.0113886 -0.0197525
+ 1.131e+11Hz -0.011413 -0.019748
+ 1.132e+11Hz -0.0114374 -0.0197435
+ 1.133e+11Hz -0.0114618 -0.0197389
+ 1.134e+11Hz -0.0114861 -0.0197342
+ 1.135e+11Hz -0.0115104 -0.0197295
+ 1.136e+11Hz -0.0115346 -0.0197248
+ 1.137e+11Hz -0.0115588 -0.01972
+ 1.138e+11Hz -0.011583 -0.0197151
+ 1.139e+11Hz -0.0116072 -0.0197102
+ 1.14e+11Hz -0.0116313 -0.0197053
+ 1.141e+11Hz -0.0116553 -0.0197003
+ 1.142e+11Hz -0.0116794 -0.0196953
+ 1.143e+11Hz -0.0117034 -0.0196902
+ 1.144e+11Hz -0.0117273 -0.0196851
+ 1.145e+11Hz -0.0117512 -0.0196799
+ 1.146e+11Hz -0.0117751 -0.0196747
+ 1.147e+11Hz -0.011799 -0.0196695
+ 1.148e+11Hz -0.0118228 -0.0196642
+ 1.149e+11Hz -0.0118465 -0.0196588
+ 1.15e+11Hz -0.0118702 -0.0196534
+ 1.151e+11Hz -0.0118939 -0.019648
+ 1.152e+11Hz -0.0119176 -0.0196425
+ 1.153e+11Hz -0.0119412 -0.019637
+ 1.154e+11Hz -0.0119647 -0.0196315
+ 1.155e+11Hz -0.0119883 -0.0196259
+ 1.156e+11Hz -0.0120117 -0.0196202
+ 1.157e+11Hz -0.0120352 -0.0196146
+ 1.158e+11Hz -0.0120586 -0.0196088
+ 1.159e+11Hz -0.0120819 -0.0196031
+ 1.16e+11Hz -0.0121053 -0.0195973
+ 1.161e+11Hz -0.0121285 -0.0195914
+ 1.162e+11Hz -0.0121518 -0.0195856
+ 1.163e+11Hz -0.012175 -0.0195797
+ 1.164e+11Hz -0.0121981 -0.0195737
+ 1.165e+11Hz -0.0122212 -0.0195677
+ 1.166e+11Hz -0.0122443 -0.0195617
+ 1.167e+11Hz -0.0122673 -0.0195556
+ 1.168e+11Hz -0.0122903 -0.0195495
+ 1.169e+11Hz -0.0123133 -0.0195434
+ 1.17e+11Hz -0.0123362 -0.0195372
+ 1.171e+11Hz -0.012359 -0.019531
+ 1.172e+11Hz -0.0123819 -0.0195248
+ 1.173e+11Hz -0.0124047 -0.0195185
+ 1.174e+11Hz -0.0124274 -0.0195122
+ 1.175e+11Hz -0.0124501 -0.0195059
+ 1.176e+11Hz -0.0124728 -0.0194995
+ 1.177e+11Hz -0.0124954 -0.0194931
+ 1.178e+11Hz -0.012518 -0.0194866
+ 1.179e+11Hz -0.0125405 -0.0194802
+ 1.18e+11Hz -0.012563 -0.0194737
+ 1.181e+11Hz -0.0125854 -0.0194671
+ 1.182e+11Hz -0.0126079 -0.0194606
+ 1.183e+11Hz -0.0126302 -0.019454
+ 1.184e+11Hz -0.0126526 -0.0194473
+ 1.185e+11Hz -0.0126749 -0.0194407
+ 1.186e+11Hz -0.0126971 -0.019434
+ 1.187e+11Hz -0.0127193 -0.0194273
+ 1.188e+11Hz -0.0127415 -0.0194205
+ 1.189e+11Hz -0.0127636 -0.0194137
+ 1.19e+11Hz -0.0127857 -0.0194069
+ 1.191e+11Hz -0.0128078 -0.0194001
+ 1.192e+11Hz -0.0128298 -0.0193932
+ 1.193e+11Hz -0.0128518 -0.0193863
+ 1.194e+11Hz -0.0128737 -0.0193794
+ 1.195e+11Hz -0.0128956 -0.0193725
+ 1.196e+11Hz -0.0129175 -0.0193655
+ 1.197e+11Hz -0.0129393 -0.0193585
+ 1.198e+11Hz -0.0129611 -0.0193515
+ 1.199e+11Hz -0.0129828 -0.0193444
+ 1.2e+11Hz -0.0130045 -0.0193373
+ 1.201e+11Hz -0.0130262 -0.0193302
+ 1.202e+11Hz -0.0130478 -0.0193231
+ 1.203e+11Hz -0.0130694 -0.0193159
+ 1.204e+11Hz -0.0130909 -0.0193088
+ 1.205e+11Hz -0.0131125 -0.0193016
+ 1.206e+11Hz -0.0131339 -0.0192943
+ 1.207e+11Hz -0.0131554 -0.0192871
+ 1.208e+11Hz -0.0131768 -0.0192798
+ 1.209e+11Hz -0.0131982 -0.0192725
+ 1.21e+11Hz -0.0132195 -0.0192651
+ 1.211e+11Hz -0.0132408 -0.0192578
+ 1.212e+11Hz -0.013262 -0.0192504
+ 1.213e+11Hz -0.0132833 -0.019243
+ 1.214e+11Hz -0.0133045 -0.0192356
+ 1.215e+11Hz -0.0133256 -0.0192281
+ 1.216e+11Hz -0.0133467 -0.0192206
+ 1.217e+11Hz -0.0133678 -0.0192131
+ 1.218e+11Hz -0.0133889 -0.0192056
+ 1.219e+11Hz -0.0134099 -0.0191981
+ 1.22e+11Hz -0.0134309 -0.0191905
+ 1.221e+11Hz -0.0134518 -0.0191829
+ 1.222e+11Hz -0.0134727 -0.0191753
+ 1.223e+11Hz -0.0134936 -0.0191676
+ 1.224e+11Hz -0.0135144 -0.01916
+ 1.225e+11Hz -0.0135353 -0.0191523
+ 1.226e+11Hz -0.013556 -0.0191446
+ 1.227e+11Hz -0.0135768 -0.0191369
+ 1.228e+11Hz -0.0135975 -0.0191291
+ 1.229e+11Hz -0.0136182 -0.0191213
+ 1.23e+11Hz -0.0136388 -0.0191135
+ 1.231e+11Hz -0.0136594 -0.0191057
+ 1.232e+11Hz -0.01368 -0.0190978
+ 1.233e+11Hz -0.0137006 -0.0190899
+ 1.234e+11Hz -0.0137211 -0.0190821
+ 1.235e+11Hz -0.0137416 -0.0190741
+ 1.236e+11Hz -0.013762 -0.0190662
+ 1.237e+11Hz -0.0137825 -0.0190582
+ 1.238e+11Hz -0.0138028 -0.0190502
+ 1.239e+11Hz -0.0138232 -0.0190422
+ 1.24e+11Hz -0.0138435 -0.0190342
+ 1.241e+11Hz -0.0138638 -0.0190261
+ 1.242e+11Hz -0.0138841 -0.019018
+ 1.243e+11Hz -0.0139043 -0.0190099
+ 1.244e+11Hz -0.0139246 -0.0190018
+ 1.245e+11Hz -0.0139447 -0.0189936
+ 1.246e+11Hz -0.0139649 -0.0189854
+ 1.247e+11Hz -0.013985 -0.0189772
+ 1.248e+11Hz -0.0140051 -0.018969
+ 1.249e+11Hz -0.0140251 -0.0189607
+ 1.25e+11Hz -0.0140452 -0.0189524
+ 1.251e+11Hz -0.0140652 -0.0189441
+ 1.252e+11Hz -0.0140851 -0.0189358
+ 1.253e+11Hz -0.0141051 -0.0189274
+ 1.254e+11Hz -0.014125 -0.018919
+ 1.255e+11Hz -0.0141448 -0.0189106
+ 1.256e+11Hz -0.0141647 -0.0189022
+ 1.257e+11Hz -0.0141845 -0.0188937
+ 1.258e+11Hz -0.0142043 -0.0188852
+ 1.259e+11Hz -0.0142241 -0.0188767
+ 1.26e+11Hz -0.0142438 -0.0188681
+ 1.261e+11Hz -0.0142635 -0.0188596
+ 1.262e+11Hz -0.0142831 -0.018851
+ 1.263e+11Hz -0.0143028 -0.0188423
+ 1.264e+11Hz -0.0143224 -0.0188337
+ 1.265e+11Hz -0.014342 -0.018825
+ 1.266e+11Hz -0.0143615 -0.0188163
+ 1.267e+11Hz -0.014381 -0.0188076
+ 1.268e+11Hz -0.0144005 -0.0187988
+ 1.269e+11Hz -0.01442 -0.01879
+ 1.27e+11Hz -0.0144394 -0.0187812
+ 1.271e+11Hz -0.0144588 -0.0187724
+ 1.272e+11Hz -0.0144781 -0.0187635
+ 1.273e+11Hz -0.0144975 -0.0187546
+ 1.274e+11Hz -0.0145168 -0.0187456
+ 1.275e+11Hz -0.014536 -0.0187367
+ 1.276e+11Hz -0.0145553 -0.0187277
+ 1.277e+11Hz -0.0145745 -0.0187187
+ 1.278e+11Hz -0.0145937 -0.0187096
+ 1.279e+11Hz -0.0146128 -0.0187005
+ 1.28e+11Hz -0.0146319 -0.0186914
+ 1.281e+11Hz -0.014651 -0.0186823
+ 1.282e+11Hz -0.01467 -0.0186731
+ 1.283e+11Hz -0.014689 -0.0186639
+ 1.284e+11Hz -0.014708 -0.0186547
+ 1.285e+11Hz -0.014727 -0.0186454
+ 1.286e+11Hz -0.0147459 -0.0186362
+ 1.287e+11Hz -0.0147648 -0.0186268
+ 1.288e+11Hz -0.0147836 -0.0186175
+ 1.289e+11Hz -0.0148024 -0.0186081
+ 1.29e+11Hz -0.0148212 -0.0185987
+ 1.291e+11Hz -0.0148399 -0.0185892
+ 1.292e+11Hz -0.0148587 -0.0185798
+ 1.293e+11Hz -0.0148773 -0.0185703
+ 1.294e+11Hz -0.014896 -0.0185607
+ 1.295e+11Hz -0.0149146 -0.0185512
+ 1.296e+11Hz -0.0149331 -0.0185416
+ 1.297e+11Hz -0.0149517 -0.0185319
+ 1.298e+11Hz -0.0149701 -0.0185223
+ 1.299e+11Hz -0.0149886 -0.0185126
+ 1.3e+11Hz -0.015007 -0.0185028
+ 1.301e+11Hz -0.0150254 -0.0184931
+ 1.302e+11Hz -0.0150437 -0.0184833
+ 1.303e+11Hz -0.015062 -0.0184735
+ 1.304e+11Hz -0.0150803 -0.0184636
+ 1.305e+11Hz -0.0150985 -0.0184537
+ 1.306e+11Hz -0.0151167 -0.0184438
+ 1.307e+11Hz -0.0151349 -0.0184339
+ 1.308e+11Hz -0.015153 -0.0184239
+ 1.309e+11Hz -0.015171 -0.0184139
+ 1.31e+11Hz -0.0151891 -0.0184039
+ 1.311e+11Hz -0.0152071 -0.0183938
+ 1.312e+11Hz -0.015225 -0.0183837
+ 1.313e+11Hz -0.0152429 -0.0183735
+ 1.314e+11Hz -0.0152608 -0.0183634
+ 1.315e+11Hz -0.0152786 -0.0183532
+ 1.316e+11Hz -0.0152963 -0.0183429
+ 1.317e+11Hz -0.0153141 -0.0183327
+ 1.318e+11Hz -0.0153318 -0.0183224
+ 1.319e+11Hz -0.0153494 -0.0183121
+ 1.32e+11Hz -0.015367 -0.0183017
+ 1.321e+11Hz -0.0153846 -0.0182913
+ 1.322e+11Hz -0.0154021 -0.0182809
+ 1.323e+11Hz -0.0154195 -0.0182705
+ 1.324e+11Hz -0.0154369 -0.01826
+ 1.325e+11Hz -0.0154543 -0.0182495
+ 1.326e+11Hz -0.0154716 -0.018239
+ 1.327e+11Hz -0.0154889 -0.0182284
+ 1.328e+11Hz -0.0155061 -0.0182178
+ 1.329e+11Hz -0.0155233 -0.0182072
+ 1.33e+11Hz -0.0155404 -0.0181966
+ 1.331e+11Hz -0.0155575 -0.0181859
+ 1.332e+11Hz -0.0155745 -0.0181752
+ 1.333e+11Hz -0.0155915 -0.0181645
+ 1.334e+11Hz -0.0156085 -0.0181537
+ 1.335e+11Hz -0.0156253 -0.0181429
+ 1.336e+11Hz -0.0156422 -0.0181321
+ 1.337e+11Hz -0.0156589 -0.0181212
+ 1.338e+11Hz -0.0156757 -0.0181104
+ 1.339e+11Hz -0.0156923 -0.0180995
+ 1.34e+11Hz -0.015709 -0.0180886
+ 1.341e+11Hz -0.0157255 -0.0180776
+ 1.342e+11Hz -0.0157421 -0.0180666
+ 1.343e+11Hz -0.0157585 -0.0180556
+ 1.344e+11Hz -0.0157749 -0.0180446
+ 1.345e+11Hz -0.0157913 -0.0180336
+ 1.346e+11Hz -0.0158076 -0.0180225
+ 1.347e+11Hz -0.0158238 -0.0180114
+ 1.348e+11Hz -0.01584 -0.0180003
+ 1.349e+11Hz -0.0158562 -0.0179892
+ 1.35e+11Hz -0.0158723 -0.017978
+ 1.351e+11Hz -0.0158883 -0.0179668
+ 1.352e+11Hz -0.0159043 -0.0179556
+ 1.353e+11Hz -0.0159202 -0.0179444
+ 1.354e+11Hz -0.015936 -0.0179332
+ 1.355e+11Hz -0.0159518 -0.0179219
+ 1.356e+11Hz -0.0159676 -0.0179106
+ 1.357e+11Hz -0.0159833 -0.0178993
+ 1.358e+11Hz -0.0159989 -0.017888
+ 1.359e+11Hz -0.0160145 -0.0178766
+ 1.36e+11Hz -0.01603 -0.0178653
+ 1.361e+11Hz -0.0160454 -0.0178539
+ 1.362e+11Hz -0.0160608 -0.0178425
+ 1.363e+11Hz -0.0160761 -0.0178311
+ 1.364e+11Hz -0.0160914 -0.0178197
+ 1.365e+11Hz -0.0161066 -0.0178082
+ 1.366e+11Hz -0.0161218 -0.0177968
+ 1.367e+11Hz -0.0161369 -0.0177853
+ 1.368e+11Hz -0.0161519 -0.0177738
+ 1.369e+11Hz -0.0161669 -0.0177623
+ 1.37e+11Hz -0.0161818 -0.0177508
+ 1.371e+11Hz -0.0161967 -0.0177393
+ 1.372e+11Hz -0.0162115 -0.0177278
+ 1.373e+11Hz -0.0162262 -0.0177162
+ 1.374e+11Hz -0.0162409 -0.0177047
+ 1.375e+11Hz -0.0162555 -0.0176931
+ 1.376e+11Hz -0.0162701 -0.0176816
+ 1.377e+11Hz -0.0162845 -0.01767
+ 1.378e+11Hz -0.016299 -0.0176584
+ 1.379e+11Hz -0.0163133 -0.0176468
+ 1.38e+11Hz -0.0163277 -0.0176352
+ 1.381e+11Hz -0.0163419 -0.0176236
+ 1.382e+11Hz -0.0163561 -0.0176119
+ 1.383e+11Hz -0.0163702 -0.0176003
+ 1.384e+11Hz -0.0163843 -0.0175887
+ 1.385e+11Hz -0.0163983 -0.0175771
+ 1.386e+11Hz -0.0164122 -0.0175654
+ 1.387e+11Hz -0.0164261 -0.0175538
+ 1.388e+11Hz -0.0164399 -0.0175421
+ 1.389e+11Hz -0.0164537 -0.0175305
+ 1.39e+11Hz -0.0164674 -0.0175188
+ 1.391e+11Hz -0.016481 -0.0175072
+ 1.392e+11Hz -0.0164946 -0.0174955
+ 1.393e+11Hz -0.0165081 -0.0174839
+ 1.394e+11Hz -0.0165215 -0.0174722
+ 1.395e+11Hz -0.0165349 -0.0174606
+ 1.396e+11Hz -0.0165482 -0.0174489
+ 1.397e+11Hz -0.0165615 -0.0174373
+ 1.398e+11Hz -0.0165747 -0.0174256
+ 1.399e+11Hz -0.0165879 -0.017414
+ 1.4e+11Hz -0.0166009 -0.0174024
+ 1.401e+11Hz -0.016614 -0.0173907
+ 1.402e+11Hz -0.0166269 -0.0173791
+ 1.403e+11Hz -0.0166398 -0.0173675
+ 1.404e+11Hz -0.0166527 -0.0173559
+ 1.405e+11Hz -0.0166655 -0.0173443
+ 1.406e+11Hz -0.0166782 -0.0173327
+ 1.407e+11Hz -0.0166908 -0.0173211
+ 1.408e+11Hz -0.0167035 -0.0173095
+ 1.409e+11Hz -0.016716 -0.0172979
+ 1.41e+11Hz -0.0167285 -0.0172863
+ 1.411e+11Hz -0.0167409 -0.0172748
+ 1.412e+11Hz -0.0167533 -0.0172632
+ 1.413e+11Hz -0.0167656 -0.0172517
+ 1.414e+11Hz -0.0167779 -0.0172402
+ 1.415e+11Hz -0.01679 -0.0172286
+ 1.416e+11Hz -0.0168022 -0.0172171
+ 1.417e+11Hz -0.0168143 -0.0172056
+ 1.418e+11Hz -0.0168263 -0.0171942
+ 1.419e+11Hz -0.0168383 -0.0171827
+ 1.42e+11Hz -0.0168502 -0.0171712
+ 1.421e+11Hz -0.016862 -0.0171598
+ 1.422e+11Hz -0.0168738 -0.0171484
+ 1.423e+11Hz -0.0168856 -0.017137
+ 1.424e+11Hz -0.0168973 -0.0171256
+ 1.425e+11Hz -0.0169089 -0.0171142
+ 1.426e+11Hz -0.0169205 -0.0171028
+ 1.427e+11Hz -0.016932 -0.0170915
+ 1.428e+11Hz -0.0169435 -0.0170801
+ 1.429e+11Hz -0.0169549 -0.0170688
+ 1.43e+11Hz -0.0169662 -0.0170575
+ 1.431e+11Hz -0.0169775 -0.0170463
+ 1.432e+11Hz -0.0169888 -0.017035
+ 1.433e+11Hz -0.017 -0.0170238
+ 1.434e+11Hz -0.0170112 -0.0170125
+ 1.435e+11Hz -0.0170223 -0.0170013
+ 1.436e+11Hz -0.0170333 -0.0169902
+ 1.437e+11Hz -0.0170443 -0.016979
+ 1.438e+11Hz -0.0170553 -0.0169679
+ 1.439e+11Hz -0.0170661 -0.0169567
+ 1.44e+11Hz -0.017077 -0.0169456
+ 1.441e+11Hz -0.0170878 -0.0169346
+ 1.442e+11Hz -0.0170985 -0.0169235
+ 1.443e+11Hz -0.0171092 -0.0169125
+ 1.444e+11Hz -0.0171199 -0.0169015
+ 1.445e+11Hz -0.0171305 -0.0168905
+ 1.446e+11Hz -0.017141 -0.0168795
+ 1.447e+11Hz -0.0171515 -0.0168686
+ 1.448e+11Hz -0.017162 -0.0168576
+ 1.449e+11Hz -0.0171724 -0.0168468
+ 1.45e+11Hz -0.0171828 -0.0168359
+ 1.451e+11Hz -0.0171931 -0.016825
+ 1.452e+11Hz -0.0172033 -0.0168142
+ 1.453e+11Hz -0.0172136 -0.0168034
+ 1.454e+11Hz -0.0172238 -0.0167926
+ 1.455e+11Hz -0.0172339 -0.0167819
+ 1.456e+11Hz -0.017244 -0.0167712
+ 1.457e+11Hz -0.017254 -0.0167605
+ 1.458e+11Hz -0.017264 -0.0167498
+ 1.459e+11Hz -0.017274 -0.0167391
+ 1.46e+11Hz -0.0172839 -0.0167285
+ 1.461e+11Hz -0.0172938 -0.0167179
+ 1.462e+11Hz -0.0173036 -0.0167073
+ 1.463e+11Hz -0.0173134 -0.0166968
+ 1.464e+11Hz -0.0173231 -0.0166863
+ 1.465e+11Hz -0.0173328 -0.0166758
+ 1.466e+11Hz -0.0173425 -0.0166653
+ 1.467e+11Hz -0.0173521 -0.0166549
+ 1.468e+11Hz -0.0173617 -0.0166445
+ 1.469e+11Hz -0.0173712 -0.0166341
+ 1.47e+11Hz -0.0173807 -0.0166237
+ 1.471e+11Hz -0.0173902 -0.0166134
+ 1.472e+11Hz -0.0173996 -0.0166031
+ 1.473e+11Hz -0.017409 -0.0165928
+ 1.474e+11Hz -0.0174183 -0.0165826
+ 1.475e+11Hz -0.0174276 -0.0165723
+ 1.476e+11Hz -0.0174369 -0.0165622
+ 1.477e+11Hz -0.0174461 -0.016552
+ 1.478e+11Hz -0.0174553 -0.0165419
+ 1.479e+11Hz -0.0174644 -0.0165317
+ 1.48e+11Hz -0.0174736 -0.0165217
+ 1.481e+11Hz -0.0174826 -0.0165116
+ 1.482e+11Hz -0.0174917 -0.0165016
+ 1.483e+11Hz -0.0175007 -0.0164916
+ 1.484e+11Hz -0.0175096 -0.0164816
+ 1.485e+11Hz -0.0175186 -0.0164717
+ 1.486e+11Hz -0.0175275 -0.0164618
+ 1.487e+11Hz -0.0175363 -0.0164519
+ 1.488e+11Hz -0.0175451 -0.0164421
+ 1.489e+11Hz -0.0175539 -0.0164322
+ 1.49e+11Hz -0.0175627 -0.0164224
+ 1.491e+11Hz -0.0175714 -0.0164127
+ 1.492e+11Hz -0.0175801 -0.016403
+ 1.493e+11Hz -0.0175887 -0.0163932
+ 1.494e+11Hz -0.0175973 -0.0163836
+ 1.495e+11Hz -0.0176059 -0.0163739
+ 1.496e+11Hz -0.0176144 -0.0163643
+ 1.497e+11Hz -0.0176229 -0.0163547
+ 1.498e+11Hz -0.0176314 -0.0163452
+ 1.499e+11Hz -0.0176399 -0.0163356
+ 1.5e+11Hz -0.0176483 -0.0163261
+ 1.501e+11Hz -0.0176566 -0.0163167
+ 1.502e+11Hz -0.017665 -0.0163072
+ 1.503e+11Hz -0.0176733 -0.0162978
+ 1.504e+11Hz -0.0176816 -0.0162885
+ 1.505e+11Hz -0.0176898 -0.0162791
+ 1.506e+11Hz -0.017698 -0.0162698
+ 1.507e+11Hz -0.0177062 -0.0162605
+ 1.508e+11Hz -0.0177144 -0.0162513
+ 1.509e+11Hz -0.0177225 -0.016242
+ 1.51e+11Hz -0.0177305 -0.0162329
+ 1.511e+11Hz -0.0177386 -0.0162237
+ 1.512e+11Hz -0.0177466 -0.0162146
+ 1.513e+11Hz -0.0177546 -0.0162055
+ 1.514e+11Hz -0.0177626 -0.0161964
+ 1.515e+11Hz -0.0177705 -0.0161874
+ 1.516e+11Hz -0.0177784 -0.0161784
+ 1.517e+11Hz -0.0177862 -0.0161694
+ 1.518e+11Hz -0.0177941 -0.0161605
+ 1.519e+11Hz -0.0178019 -0.0161516
+ 1.52e+11Hz -0.0178096 -0.0161427
+ 1.521e+11Hz -0.0178174 -0.0161338
+ 1.522e+11Hz -0.0178251 -0.016125
+ 1.523e+11Hz -0.0178327 -0.0161163
+ 1.524e+11Hz -0.0178404 -0.0161075
+ 1.525e+11Hz -0.017848 -0.0160988
+ 1.526e+11Hz -0.0178556 -0.0160901
+ 1.527e+11Hz -0.0178631 -0.0160815
+ 1.528e+11Hz -0.0178707 -0.0160729
+ 1.529e+11Hz -0.0178781 -0.0160643
+ 1.53e+11Hz -0.0178856 -0.0160558
+ 1.531e+11Hz -0.017893 -0.0160473
+ 1.532e+11Hz -0.0179004 -0.0160388
+ 1.533e+11Hz -0.0179078 -0.0160304
+ 1.534e+11Hz -0.0179152 -0.016022
+ 1.535e+11Hz -0.0179225 -0.0160137
+ 1.536e+11Hz -0.0179298 -0.0160053
+ 1.537e+11Hz -0.017937 -0.0159971
+ 1.538e+11Hz -0.0179442 -0.0159888
+ 1.539e+11Hz -0.0179514 -0.0159806
+ 1.54e+11Hz -0.0179586 -0.0159724
+ 1.541e+11Hz -0.0179657 -0.0159643
+ 1.542e+11Hz -0.0179728 -0.0159562
+ 1.543e+11Hz -0.0179799 -0.0159481
+ 1.544e+11Hz -0.017987 -0.0159401
+ 1.545e+11Hz -0.017994 -0.0159321
+ 1.546e+11Hz -0.018001 -0.0159242
+ 1.547e+11Hz -0.018008 -0.0159163
+ 1.548e+11Hz -0.0180149 -0.0159084
+ 1.549e+11Hz -0.0180218 -0.0159006
+ 1.55e+11Hz -0.0180287 -0.0158928
+ 1.551e+11Hz -0.0180355 -0.0158851
+ 1.552e+11Hz -0.0180424 -0.0158774
+ 1.553e+11Hz -0.0180492 -0.0158697
+ 1.554e+11Hz -0.0180559 -0.0158621
+ 1.555e+11Hz -0.0180627 -0.0158546
+ 1.556e+11Hz -0.0180694 -0.015847
+ 1.557e+11Hz -0.0180761 -0.0158396
+ 1.558e+11Hz -0.0180828 -0.0158321
+ 1.559e+11Hz -0.0180894 -0.0158247
+ 1.56e+11Hz -0.018096 -0.0158174
+ 1.561e+11Hz -0.0181026 -0.0158101
+ 1.562e+11Hz -0.0181092 -0.0158028
+ 1.563e+11Hz -0.0181157 -0.0157956
+ 1.564e+11Hz -0.0181222 -0.0157885
+ 1.565e+11Hz -0.0181287 -0.0157814
+ 1.566e+11Hz -0.0181352 -0.0157743
+ 1.567e+11Hz -0.0181416 -0.0157673
+ 1.568e+11Hz -0.018148 -0.0157603
+ 1.569e+11Hz -0.0181544 -0.0157534
+ 1.57e+11Hz -0.0181608 -0.0157465
+ 1.571e+11Hz -0.0181672 -0.0157397
+ 1.572e+11Hz -0.0181735 -0.0157329
+ 1.573e+11Hz -0.0181798 -0.0157262
+ 1.574e+11Hz -0.0181861 -0.0157196
+ 1.575e+11Hz -0.0181924 -0.0157129
+ 1.576e+11Hz -0.0181986 -0.0157064
+ 1.577e+11Hz -0.0182048 -0.0156999
+ 1.578e+11Hz -0.018211 -0.0156934
+ 1.579e+11Hz -0.0182172 -0.015687
+ 1.58e+11Hz -0.0182234 -0.0156807
+ 1.581e+11Hz -0.0182295 -0.0156744
+ 1.582e+11Hz -0.0182357 -0.0156682
+ 1.583e+11Hz -0.0182418 -0.015662
+ 1.584e+11Hz -0.0182479 -0.0156559
+ 1.585e+11Hz -0.018254 -0.0156498
+ 1.586e+11Hz -0.01826 -0.0156438
+ 1.587e+11Hz -0.0182661 -0.0156379
+ 1.588e+11Hz -0.0182721 -0.015632
+ 1.589e+11Hz -0.0182781 -0.0156262
+ 1.59e+11Hz -0.0182842 -0.0156204
+ 1.591e+11Hz -0.0182901 -0.0156147
+ 1.592e+11Hz -0.0182961 -0.0156091
+ 1.593e+11Hz -0.0183021 -0.0156035
+ 1.594e+11Hz -0.0183081 -0.015598
+ 1.595e+11Hz -0.018314 -0.0155925
+ 1.596e+11Hz -0.01832 -0.0155871
+ 1.597e+11Hz -0.0183259 -0.0155818
+ 1.598e+11Hz -0.0183318 -0.0155765
+ 1.599e+11Hz -0.0183378 -0.0155713
+ 1.6e+11Hz -0.0183437 -0.0155662
+ 1.601e+11Hz -0.0183496 -0.0155611
+ 1.602e+11Hz -0.0183555 -0.0155561
+ 1.603e+11Hz -0.0183614 -0.0155512
+ 1.604e+11Hz -0.0183673 -0.0155463
+ 1.605e+11Hz -0.0183732 -0.0155415
+ 1.606e+11Hz -0.0183791 -0.0155368
+ 1.607e+11Hz -0.018385 -0.0155321
+ 1.608e+11Hz -0.0183909 -0.0155275
+ 1.609e+11Hz -0.0183967 -0.0155229
+ 1.61e+11Hz -0.0184026 -0.0155185
+ 1.611e+11Hz -0.0184085 -0.0155141
+ 1.612e+11Hz -0.0184144 -0.0155098
+ 1.613e+11Hz -0.0184204 -0.0155055
+ 1.614e+11Hz -0.0184263 -0.0155013
+ 1.615e+11Hz -0.0184322 -0.0154972
+ 1.616e+11Hz -0.0184381 -0.0154932
+ 1.617e+11Hz -0.0184441 -0.0154892
+ 1.618e+11Hz -0.01845 -0.0154853
+ 1.619e+11Hz -0.018456 -0.0154814
+ 1.62e+11Hz -0.0184619 -0.0154777
+ 1.621e+11Hz -0.0184679 -0.015474
+ 1.622e+11Hz -0.0184739 -0.0154704
+ 1.623e+11Hz -0.0184799 -0.0154668
+ 1.624e+11Hz -0.0184859 -0.0154634
+ 1.625e+11Hz -0.018492 -0.01546
+ 1.626e+11Hz -0.018498 -0.0154567
+ 1.627e+11Hz -0.0185041 -0.0154534
+ 1.628e+11Hz -0.0185102 -0.0154502
+ 1.629e+11Hz -0.0185164 -0.0154471
+ 1.63e+11Hz -0.0185225 -0.0154441
+ 1.631e+11Hz -0.0185287 -0.0154411
+ 1.632e+11Hz -0.0185349 -0.0154383
+ 1.633e+11Hz -0.0185411 -0.0154354
+ 1.634e+11Hz -0.0185473 -0.0154327
+ 1.635e+11Hz -0.0185536 -0.01543
+ 1.636e+11Hz -0.0185599 -0.0154275
+ 1.637e+11Hz -0.0185663 -0.0154249
+ 1.638e+11Hz -0.0185726 -0.0154225
+ 1.639e+11Hz -0.018579 -0.0154201
+ 1.64e+11Hz -0.0185855 -0.0154178
+ 1.641e+11Hz -0.018592 -0.0154156
+ 1.642e+11Hz -0.0185985 -0.0154135
+ 1.643e+11Hz -0.018605 -0.0154114
+ 1.644e+11Hz -0.0186116 -0.0154094
+ 1.645e+11Hz -0.0186183 -0.0154075
+ 1.646e+11Hz -0.0186249 -0.0154056
+ 1.647e+11Hz -0.0186316 -0.0154038
+ 1.648e+11Hz -0.0186384 -0.0154021
+ 1.649e+11Hz -0.0186452 -0.0154005
+ 1.65e+11Hz -0.0186521 -0.0153989
+ 1.651e+11Hz -0.018659 -0.0153974
+ 1.652e+11Hz -0.0186659 -0.0153959
+ 1.653e+11Hz -0.0186729 -0.0153946
+ 1.654e+11Hz -0.01868 -0.0153933
+ 1.655e+11Hz -0.0186871 -0.0153921
+ 1.656e+11Hz -0.0186943 -0.0153909
+ 1.657e+11Hz -0.0187015 -0.0153898
+ 1.658e+11Hz -0.0187088 -0.0153888
+ 1.659e+11Hz -0.0187161 -0.0153878
+ 1.66e+11Hz -0.0187235 -0.015387
+ 1.661e+11Hz -0.018731 -0.0153861
+ 1.662e+11Hz -0.0187385 -0.0153854
+ 1.663e+11Hz -0.0187461 -0.0153847
+ 1.664e+11Hz -0.0187538 -0.0153841
+ 1.665e+11Hz -0.0187615 -0.0153835
+ 1.666e+11Hz -0.0187693 -0.015383
+ 1.667e+11Hz -0.0187771 -0.0153826
+ 1.668e+11Hz -0.0187851 -0.0153822
+ 1.669e+11Hz -0.0187931 -0.0153819
+ 1.67e+11Hz -0.0188011 -0.0153816
+ 1.671e+11Hz -0.0188093 -0.0153814
+ 1.672e+11Hz -0.0188175 -0.0153813
+ 1.673e+11Hz -0.0188258 -0.0153812
+ 1.674e+11Hz -0.0188342 -0.0153812
+ 1.675e+11Hz -0.0188426 -0.0153812
+ 1.676e+11Hz -0.0188512 -0.0153813
+ 1.677e+11Hz -0.0188598 -0.0153814
+ 1.678e+11Hz -0.0188685 -0.0153816
+ 1.679e+11Hz -0.0188773 -0.0153818
+ 1.68e+11Hz -0.0188861 -0.0153821
+ 1.681e+11Hz -0.0188951 -0.0153825
+ 1.682e+11Hz -0.0189041 -0.0153828
+ 1.683e+11Hz -0.0189132 -0.0153833
+ 1.684e+11Hz -0.0189225 -0.0153837
+ 1.685e+11Hz -0.0189318 -0.0153843
+ 1.686e+11Hz -0.0189412 -0.0153848
+ 1.687e+11Hz -0.0189506 -0.0153854
+ 1.688e+11Hz -0.0189602 -0.0153861
+ 1.689e+11Hz -0.0189699 -0.0153868
+ 1.69e+11Hz -0.0189797 -0.0153875
+ 1.691e+11Hz -0.0189895 -0.0153883
+ 1.692e+11Hz -0.0189995 -0.0153891
+ 1.693e+11Hz -0.0190095 -0.0153899
+ 1.694e+11Hz -0.0190197 -0.0153908
+ 1.695e+11Hz -0.01903 -0.0153917
+ 1.696e+11Hz -0.0190403 -0.0153926
+ 1.697e+11Hz -0.0190508 -0.0153936
+ 1.698e+11Hz -0.0190613 -0.0153946
+ 1.699e+11Hz -0.019072 -0.0153956
+ 1.7e+11Hz -0.0190828 -0.0153966
+ 1.701e+11Hz -0.0190936 -0.0153977
+ 1.702e+11Hz -0.0191046 -0.0153988
+ 1.703e+11Hz -0.0191157 -0.0153999
+ 1.704e+11Hz -0.0191269 -0.015401
+ 1.705e+11Hz -0.0191382 -0.0154022
+ 1.706e+11Hz -0.0191496 -0.0154034
+ 1.707e+11Hz -0.0191611 -0.0154045
+ 1.708e+11Hz -0.0191727 -0.0154057
+ 1.709e+11Hz -0.0191844 -0.0154069
+ 1.71e+11Hz -0.0191963 -0.0154081
+ 1.711e+11Hz -0.0192082 -0.0154094
+ 1.712e+11Hz -0.0192203 -0.0154106
+ 1.713e+11Hz -0.0192325 -0.0154118
+ 1.714e+11Hz -0.0192447 -0.0154131
+ 1.715e+11Hz -0.0192571 -0.0154143
+ 1.716e+11Hz -0.0192696 -0.0154155
+ 1.717e+11Hz -0.0192823 -0.0154168
+ 1.718e+11Hz -0.019295 -0.015418
+ 1.719e+11Hz -0.0193079 -0.0154192
+ 1.72e+11Hz -0.0193208 -0.0154205
+ 1.721e+11Hz -0.0193339 -0.0154217
+ 1.722e+11Hz -0.0193471 -0.0154229
+ 1.723e+11Hz -0.0193604 -0.0154241
+ 1.724e+11Hz -0.0193738 -0.0154252
+ 1.725e+11Hz -0.0193874 -0.0154264
+ 1.726e+11Hz -0.019401 -0.0154276
+ 1.727e+11Hz -0.0194148 -0.0154287
+ 1.728e+11Hz -0.0194287 -0.0154298
+ 1.729e+11Hz -0.0194427 -0.0154309
+ 1.73e+11Hz -0.0194568 -0.0154319
+ 1.731e+11Hz -0.019471 -0.015433
+ 1.732e+11Hz -0.0194854 -0.015434
+ 1.733e+11Hz -0.0194999 -0.015435
+ 1.734e+11Hz -0.0195144 -0.0154359
+ 1.735e+11Hz -0.0195291 -0.0154368
+ 1.736e+11Hz -0.0195439 -0.0154377
+ 1.737e+11Hz -0.0195589 -0.0154386
+ 1.738e+11Hz -0.0195739 -0.0154394
+ 1.739e+11Hz -0.019589 -0.0154402
+ 1.74e+11Hz -0.0196043 -0.0154409
+ 1.741e+11Hz -0.0196197 -0.0154416
+ 1.742e+11Hz -0.0196352 -0.0154422
+ 1.743e+11Hz -0.0196508 -0.0154428
+ 1.744e+11Hz -0.0196665 -0.0154434
+ 1.745e+11Hz -0.0196823 -0.0154439
+ 1.746e+11Hz -0.0196983 -0.0154443
+ 1.747e+11Hz -0.0197143 -0.0154447
+ 1.748e+11Hz -0.0197305 -0.015445
+ 1.749e+11Hz -0.0197468 -0.0154453
+ 1.75e+11Hz -0.0197632 -0.0154455
+ 1.751e+11Hz -0.0197797 -0.0154457
+ 1.752e+11Hz -0.0197963 -0.0154458
+ 1.753e+11Hz -0.019813 -0.0154459
+ 1.754e+11Hz -0.0198298 -0.0154458
+ 1.755e+11Hz -0.0198467 -0.0154457
+ 1.756e+11Hz -0.0198637 -0.0154456
+ 1.757e+11Hz -0.0198809 -0.0154453
+ 1.758e+11Hz -0.0198981 -0.015445
+ 1.759e+11Hz -0.0199154 -0.0154447
+ 1.76e+11Hz -0.0199329 -0.0154442
+ 1.761e+11Hz -0.0199504 -0.0154437
+ 1.762e+11Hz -0.0199681 -0.0154431
+ 1.763e+11Hz -0.0199858 -0.0154424
+ 1.764e+11Hz -0.0200037 -0.0154416
+ 1.765e+11Hz -0.0200216 -0.0154408
+ 1.766e+11Hz -0.0200397 -0.0154399
+ 1.767e+11Hz -0.0200578 -0.0154389
+ 1.768e+11Hz -0.020076 -0.0154378
+ 1.769e+11Hz -0.0200943 -0.0154366
+ 1.77e+11Hz -0.0201128 -0.0154353
+ 1.771e+11Hz -0.0201313 -0.0154339
+ 1.772e+11Hz -0.0201499 -0.0154325
+ 1.773e+11Hz -0.0201685 -0.0154309
+ 1.774e+11Hz -0.0201873 -0.0154293
+ 1.775e+11Hz -0.0202062 -0.0154275
+ 1.776e+11Hz -0.0202251 -0.0154257
+ 1.777e+11Hz -0.0202442 -0.0154237
+ 1.778e+11Hz -0.0202633 -0.0154217
+ 1.779e+11Hz -0.0202825 -0.0154196
+ 1.78e+11Hz -0.0203018 -0.0154173
+ 1.781e+11Hz -0.0203211 -0.015415
+ 1.782e+11Hz -0.0203406 -0.0154125
+ 1.783e+11Hz -0.0203601 -0.01541
+ 1.784e+11Hz -0.0203797 -0.0154073
+ 1.785e+11Hz -0.0203993 -0.0154045
+ 1.786e+11Hz -0.0204191 -0.0154016
+ 1.787e+11Hz -0.0204389 -0.0153986
+ 1.788e+11Hz -0.0204588 -0.0153955
+ 1.789e+11Hz -0.0204787 -0.0153923
+ 1.79e+11Hz -0.0204987 -0.015389
+ 1.791e+11Hz -0.0205188 -0.0153855
+ 1.792e+11Hz -0.0205389 -0.015382
+ 1.793e+11Hz -0.0205592 -0.0153783
+ 1.794e+11Hz -0.0205794 -0.0153745
+ 1.795e+11Hz -0.0205997 -0.0153706
+ 1.796e+11Hz -0.0206201 -0.0153666
+ 1.797e+11Hz -0.0206406 -0.0153624
+ 1.798e+11Hz -0.0206611 -0.0153581
+ 1.799e+11Hz -0.0206816 -0.0153538
+ 1.8e+11Hz -0.0207022 -0.0153492
+ 1.801e+11Hz -0.0207229 -0.0153446
+ 1.802e+11Hz -0.0207436 -0.0153399
+ 1.803e+11Hz -0.0207643 -0.015335
+ 1.804e+11Hz -0.0207851 -0.01533
+ 1.805e+11Hz -0.020806 -0.0153248
+ 1.806e+11Hz -0.0208269 -0.0153196
+ 1.807e+11Hz -0.0208478 -0.0153142
+ 1.808e+11Hz -0.0208688 -0.0153087
+ 1.809e+11Hz -0.0208898 -0.015303
+ 1.81e+11Hz -0.0209108 -0.0152973
+ 1.811e+11Hz -0.0209319 -0.0152914
+ 1.812e+11Hz -0.020953 -0.0152854
+ 1.813e+11Hz -0.0209741 -0.0152792
+ 1.814e+11Hz -0.0209953 -0.0152729
+ 1.815e+11Hz -0.0210165 -0.0152665
+ 1.816e+11Hz -0.0210377 -0.01526
+ 1.817e+11Hz -0.0210589 -0.0152533
+ 1.818e+11Hz -0.0210802 -0.0152465
+ 1.819e+11Hz -0.0211015 -0.0152396
+ 1.82e+11Hz -0.0211228 -0.0152325
+ 1.821e+11Hz -0.0211441 -0.0152253
+ 1.822e+11Hz -0.0211655 -0.015218
+ 1.823e+11Hz -0.0211868 -0.0152105
+ 1.824e+11Hz -0.0212082 -0.0152029
+ 1.825e+11Hz -0.0212296 -0.0151952
+ 1.826e+11Hz -0.021251 -0.0151874
+ 1.827e+11Hz -0.0212724 -0.0151794
+ 1.828e+11Hz -0.0212938 -0.0151713
+ 1.829e+11Hz -0.0213152 -0.015163
+ 1.83e+11Hz -0.0213367 -0.0151546
+ 1.831e+11Hz -0.0213581 -0.0151461
+ 1.832e+11Hz -0.0213795 -0.0151375
+ 1.833e+11Hz -0.0214009 -0.0151287
+ 1.834e+11Hz -0.0214223 -0.0151198
+ 1.835e+11Hz -0.0214438 -0.0151107
+ 1.836e+11Hz -0.0214652 -0.0151016
+ 1.837e+11Hz -0.0214866 -0.0150923
+ 1.838e+11Hz -0.021508 -0.0150828
+ 1.839e+11Hz -0.0215293 -0.0150733
+ 1.84e+11Hz -0.0215507 -0.0150636
+ 1.841e+11Hz -0.0215721 -0.0150538
+ 1.842e+11Hz -0.0215934 -0.0150438
+ 1.843e+11Hz -0.0216147 -0.0150337
+ 1.844e+11Hz -0.021636 -0.0150235
+ 1.845e+11Hz -0.0216573 -0.0150132
+ 1.846e+11Hz -0.0216786 -0.0150027
+ 1.847e+11Hz -0.0216998 -0.0149921
+ 1.848e+11Hz -0.021721 -0.0149814
+ 1.849e+11Hz -0.0217422 -0.0149705
+ 1.85e+11Hz -0.0217634 -0.0149595
+ 1.851e+11Hz -0.0217845 -0.0149484
+ 1.852e+11Hz -0.0218057 -0.0149372
+ 1.853e+11Hz -0.0218267 -0.0149258
+ 1.854e+11Hz -0.0218478 -0.0149144
+ 1.855e+11Hz -0.0218688 -0.0149028
+ 1.856e+11Hz -0.0218898 -0.014891
+ 1.857e+11Hz -0.0219107 -0.0148792
+ 1.858e+11Hz -0.0219316 -0.0148672
+ 1.859e+11Hz -0.0219525 -0.0148551
+ 1.86e+11Hz -0.0219733 -0.0148429
+ 1.861e+11Hz -0.0219941 -0.0148306
+ 1.862e+11Hz -0.0220148 -0.0148181
+ 1.863e+11Hz -0.0220355 -0.0148055
+ 1.864e+11Hz -0.0220561 -0.0147928
+ 1.865e+11Hz -0.0220767 -0.01478
+ 1.866e+11Hz -0.0220973 -0.0147671
+ 1.867e+11Hz -0.0221178 -0.014754
+ 1.868e+11Hz -0.0221382 -0.0147409
+ 1.869e+11Hz -0.0221586 -0.0147276
+ 1.87e+11Hz -0.022179 -0.0147142
+ 1.871e+11Hz -0.0221993 -0.0147007
+ 1.872e+11Hz -0.0222195 -0.0146871
+ 1.873e+11Hz -0.0222397 -0.0146734
+ 1.874e+11Hz -0.0222598 -0.0146595
+ 1.875e+11Hz -0.0222799 -0.0146456
+ 1.876e+11Hz -0.0222999 -0.0146315
+ 1.877e+11Hz -0.0223198 -0.0146174
+ 1.878e+11Hz -0.0223397 -0.0146031
+ 1.879e+11Hz -0.0223595 -0.0145887
+ 1.88e+11Hz -0.0223793 -0.0145742
+ 1.881e+11Hz -0.022399 -0.0145597
+ 1.882e+11Hz -0.0224186 -0.014545
+ 1.883e+11Hz -0.0224381 -0.0145302
+ 1.884e+11Hz -0.0224576 -0.0145153
+ 1.885e+11Hz -0.022477 -0.0145003
+ 1.886e+11Hz -0.0224964 -0.0144852
+ 1.887e+11Hz -0.0225157 -0.01447
+ 1.888e+11Hz -0.0225349 -0.0144547
+ 1.889e+11Hz -0.022554 -0.0144393
+ 1.89e+11Hz -0.0225731 -0.0144238
+ 1.891e+11Hz -0.0225921 -0.0144082
+ 1.892e+11Hz -0.022611 -0.0143926
+ 1.893e+11Hz -0.0226298 -0.0143768
+ 1.894e+11Hz -0.0226486 -0.0143609
+ 1.895e+11Hz -0.0226673 -0.014345
+ 1.896e+11Hz -0.0226859 -0.0143289
+ 1.897e+11Hz -0.0227044 -0.0143128
+ 1.898e+11Hz -0.0227228 -0.0142966
+ 1.899e+11Hz -0.0227412 -0.0142803
+ 1.9e+11Hz -0.0227595 -0.0142639
+ 1.901e+11Hz -0.0227777 -0.0142474
+ 1.902e+11Hz -0.0227958 -0.0142308
+ 1.903e+11Hz -0.0228138 -0.0142142
+ 1.904e+11Hz -0.0228318 -0.0141975
+ 1.905e+11Hz -0.0228496 -0.0141807
+ 1.906e+11Hz -0.0228674 -0.0141638
+ 1.907e+11Hz -0.0228851 -0.0141468
+ 1.908e+11Hz -0.0229027 -0.0141298
+ 1.909e+11Hz -0.0229203 -0.0141127
+ 1.91e+11Hz -0.0229377 -0.0140955
+ 1.911e+11Hz -0.022955 -0.0140782
+ 1.912e+11Hz -0.0229723 -0.0140609
+ 1.913e+11Hz -0.0229894 -0.0140434
+ 1.914e+11Hz -0.0230065 -0.014026
+ 1.915e+11Hz -0.0230235 -0.0140084
+ 1.916e+11Hz -0.0230404 -0.0139908
+ 1.917e+11Hz -0.0230572 -0.0139731
+ 1.918e+11Hz -0.0230739 -0.0139553
+ 1.919e+11Hz -0.0230905 -0.0139375
+ 1.92e+11Hz -0.0231071 -0.0139196
+ 1.921e+11Hz -0.0231235 -0.0139017
+ 1.922e+11Hz -0.0231398 -0.0138837
+ 1.923e+11Hz -0.0231561 -0.0138656
+ 1.924e+11Hz -0.0231722 -0.0138475
+ 1.925e+11Hz -0.0231883 -0.0138293
+ 1.926e+11Hz -0.0232042 -0.013811
+ 1.927e+11Hz -0.0232201 -0.0137927
+ 1.928e+11Hz -0.0232359 -0.0137744
+ 1.929e+11Hz -0.0232516 -0.013756
+ 1.93e+11Hz -0.0232671 -0.0137375
+ 1.931e+11Hz -0.0232826 -0.013719
+ 1.932e+11Hz -0.023298 -0.0137004
+ 1.933e+11Hz -0.0233133 -0.0136818
+ 1.934e+11Hz -0.0233285 -0.0136631
+ 1.935e+11Hz -0.0233435 -0.0136444
+ 1.936e+11Hz -0.0233585 -0.0136257
+ 1.937e+11Hz -0.0233734 -0.0136069
+ 1.938e+11Hz -0.0233882 -0.013588
+ 1.939e+11Hz -0.0234029 -0.0135691
+ 1.94e+11Hz -0.0234175 -0.0135502
+ 1.941e+11Hz -0.023432 -0.0135312
+ 1.942e+11Hz -0.0234464 -0.0135122
+ 1.943e+11Hz -0.0234607 -0.0134932
+ 1.944e+11Hz -0.0234749 -0.0134741
+ 1.945e+11Hz -0.023489 -0.013455
+ 1.946e+11Hz -0.023503 -0.0134358
+ 1.947e+11Hz -0.0235169 -0.0134167
+ 1.948e+11Hz -0.0235307 -0.0133974
+ 1.949e+11Hz -0.0235444 -0.0133782
+ 1.95e+11Hz -0.023558 -0.0133589
+ 1.951e+11Hz -0.0235714 -0.0133396
+ 1.952e+11Hz -0.0235848 -0.0133203
+ 1.953e+11Hz -0.0235981 -0.0133009
+ 1.954e+11Hz -0.0236113 -0.0132815
+ 1.955e+11Hz -0.0236244 -0.0132621
+ 1.956e+11Hz -0.0236374 -0.0132427
+ 1.957e+11Hz -0.0236503 -0.0132232
+ 1.958e+11Hz -0.0236631 -0.0132038
+ 1.959e+11Hz -0.0236758 -0.0131843
+ 1.96e+11Hz -0.0236884 -0.0131648
+ 1.961e+11Hz -0.0237009 -0.0131453
+ 1.962e+11Hz -0.0237132 -0.0131257
+ 1.963e+11Hz -0.0237255 -0.0131062
+ 1.964e+11Hz -0.0237377 -0.0130866
+ 1.965e+11Hz -0.0237498 -0.013067
+ 1.966e+11Hz -0.0237618 -0.0130474
+ 1.967e+11Hz -0.0237737 -0.0130278
+ 1.968e+11Hz -0.0237855 -0.0130082
+ 1.969e+11Hz -0.0237972 -0.0129886
+ 1.97e+11Hz -0.0238088 -0.012969
+ 1.971e+11Hz -0.0238202 -0.0129494
+ 1.972e+11Hz -0.0238316 -0.0129297
+ 1.973e+11Hz -0.0238429 -0.0129101
+ 1.974e+11Hz -0.0238541 -0.0128905
+ 1.975e+11Hz -0.0238652 -0.0128709
+ 1.976e+11Hz -0.0238762 -0.0128512
+ 1.977e+11Hz -0.0238871 -0.0128316
+ 1.978e+11Hz -0.0238979 -0.012812
+ 1.979e+11Hz -0.0239087 -0.0127924
+ 1.98e+11Hz -0.0239193 -0.0127728
+ 1.981e+11Hz -0.0239298 -0.0127532
+ 1.982e+11Hz -0.0239402 -0.0127336
+ 1.983e+11Hz -0.0239505 -0.012714
+ 1.984e+11Hz -0.0239608 -0.0126944
+ 1.985e+11Hz -0.0239709 -0.0126749
+ 1.986e+11Hz -0.023981 -0.0126553
+ 1.987e+11Hz -0.0239909 -0.0126358
+ 1.988e+11Hz -0.0240008 -0.0126163
+ 1.989e+11Hz -0.0240105 -0.0125968
+ 1.99e+11Hz -0.0240202 -0.0125773
+ 1.991e+11Hz -0.0240298 -0.0125579
+ 1.992e+11Hz -0.0240393 -0.0125385
+ 1.993e+11Hz -0.0240487 -0.012519
+ 1.994e+11Hz -0.024058 -0.0124997
+ 1.995e+11Hz -0.0240672 -0.0124803
+ 1.996e+11Hz -0.0240764 -0.0124609
+ 1.997e+11Hz -0.0240854 -0.0124416
+ 1.998e+11Hz -0.0240944 -0.0124224
+ 1.999e+11Hz -0.0241033 -0.0124031
+ 2e+11Hz -0.0241121 -0.0123839
+ 2.001e+11Hz -0.0241208 -0.0123647
+ 2.002e+11Hz -0.0241294 -0.0123455
+ 2.003e+11Hz -0.0241379 -0.0123264
+ 2.004e+11Hz -0.0241464 -0.0123073
+ 2.005e+11Hz -0.0241548 -0.0122883
+ 2.006e+11Hz -0.0241631 -0.0122693
+ 2.007e+11Hz -0.0241713 -0.0122503
+ 2.008e+11Hz -0.0241794 -0.0122313
+ 2.009e+11Hz -0.0241875 -0.0122124
+ 2.01e+11Hz -0.0241955 -0.0121936
+ 2.011e+11Hz -0.0242034 -0.0121748
+ 2.012e+11Hz -0.0242112 -0.012156
+ 2.013e+11Hz -0.024219 -0.0121373
+ 2.014e+11Hz -0.0242267 -0.0121186
+ 2.015e+11Hz -0.0242343 -0.0121
+ 2.016e+11Hz -0.0242418 -0.0120814
+ 2.017e+11Hz -0.0242493 -0.0120629
+ 2.018e+11Hz -0.0242567 -0.0120444
+ 2.019e+11Hz -0.024264 -0.012026
+ 2.02e+11Hz -0.0242713 -0.0120076
+ 2.021e+11Hz -0.0242785 -0.0119893
+ 2.022e+11Hz -0.0242856 -0.011971
+ 2.023e+11Hz -0.0242927 -0.0119528
+ 2.024e+11Hz -0.0242997 -0.0119347
+ 2.025e+11Hz -0.0243067 -0.0119166
+ 2.026e+11Hz -0.0243136 -0.0118985
+ 2.027e+11Hz -0.0243204 -0.0118805
+ 2.028e+11Hz -0.0243272 -0.0118626
+ 2.029e+11Hz -0.0243339 -0.0118448
+ 2.03e+11Hz -0.0243406 -0.011827
+ 2.031e+11Hz -0.0243472 -0.0118093
+ 2.032e+11Hz -0.0243538 -0.0117916
+ 2.033e+11Hz -0.0243603 -0.011774
+ 2.034e+11Hz -0.0243668 -0.0117564
+ 2.035e+11Hz -0.0243732 -0.011739
+ 2.036e+11Hz -0.0243796 -0.0117216
+ 2.037e+11Hz -0.0243859 -0.0117042
+ 2.038e+11Hz -0.0243922 -0.011687
+ 2.039e+11Hz -0.0243984 -0.0116698
+ 2.04e+11Hz -0.0244046 -0.0116526
+ 2.041e+11Hz -0.0244108 -0.0116356
+ 2.042e+11Hz -0.024417 -0.0116186
+ 2.043e+11Hz -0.0244231 -0.0116017
+ 2.044e+11Hz -0.0244291 -0.0115848
+ 2.045e+11Hz -0.0244352 -0.0115681
+ 2.046e+11Hz -0.0244412 -0.0115514
+ 2.047e+11Hz -0.0244472 -0.0115348
+ 2.048e+11Hz -0.0244531 -0.0115182
+ 2.049e+11Hz -0.0244591 -0.0115017
+ 2.05e+11Hz -0.024465 -0.0114853
+ 2.051e+11Hz -0.0244709 -0.011469
+ 2.052e+11Hz -0.0244767 -0.0114528
+ 2.053e+11Hz -0.0244826 -0.0114366
+ 2.054e+11Hz -0.0244884 -0.0114205
+ 2.055e+11Hz -0.0244943 -0.0114045
+ 2.056e+11Hz -0.0245001 -0.0113886
+ 2.057e+11Hz -0.0245059 -0.0113727
+ 2.058e+11Hz -0.0245117 -0.0113569
+ 2.059e+11Hz -0.0245175 -0.0113412
+ 2.06e+11Hz -0.0245233 -0.0113256
+ 2.061e+11Hz -0.0245291 -0.0113101
+ 2.062e+11Hz -0.0245349 -0.0112946
+ 2.063e+11Hz -0.0245407 -0.0112792
+ 2.064e+11Hz -0.0245465 -0.0112639
+ 2.065e+11Hz -0.0245523 -0.0112487
+ 2.066e+11Hz -0.0245581 -0.0112335
+ 2.067e+11Hz -0.0245639 -0.0112184
+ 2.068e+11Hz -0.0245698 -0.0112034
+ 2.069e+11Hz -0.0245756 -0.0111885
+ 2.07e+11Hz -0.0245815 -0.0111737
+ 2.071e+11Hz -0.0245874 -0.0111589
+ 2.072e+11Hz -0.0245933 -0.0111442
+ 2.073e+11Hz -0.0245993 -0.0111296
+ 2.074e+11Hz -0.0246052 -0.0111151
+ 2.075e+11Hz -0.0246112 -0.0111006
+ 2.076e+11Hz -0.0246172 -0.0110862
+ 2.077e+11Hz -0.0246233 -0.0110719
+ 2.078e+11Hz -0.0246294 -0.0110577
+ 2.079e+11Hz -0.0246355 -0.0110435
+ 2.08e+11Hz -0.0246417 -0.0110294
+ 2.081e+11Hz -0.0246479 -0.0110154
+ 2.082e+11Hz -0.0246541 -0.0110014
+ 2.083e+11Hz -0.0246604 -0.0109876
+ 2.084e+11Hz -0.0246667 -0.0109738
+ 2.085e+11Hz -0.0246731 -0.01096
+ 2.086e+11Hz -0.0246795 -0.0109464
+ 2.087e+11Hz -0.024686 -0.0109328
+ 2.088e+11Hz -0.0246926 -0.0109192
+ 2.089e+11Hz -0.0246992 -0.0109058
+ 2.09e+11Hz -0.0247058 -0.0108923
+ 2.091e+11Hz -0.0247125 -0.010879
+ 2.092e+11Hz -0.0247193 -0.0108657
+ 2.093e+11Hz -0.0247262 -0.0108525
+ 2.094e+11Hz -0.0247331 -0.0108393
+ 2.095e+11Hz -0.0247401 -0.0108262
+ 2.096e+11Hz -0.0247471 -0.0108132
+ 2.097e+11Hz -0.0247543 -0.0108002
+ 2.098e+11Hz -0.0247615 -0.0107873
+ 2.099e+11Hz -0.0247688 -0.0107744
+ 2.1e+11Hz -0.0247761 -0.0107615
+ 2.101e+11Hz -0.0247836 -0.0107488
+ 2.102e+11Hz -0.0247911 -0.010736
+ 2.103e+11Hz -0.0247988 -0.0107233
+ 2.104e+11Hz -0.0248065 -0.0107107
+ 2.105e+11Hz -0.0248143 -0.0106981
+ 2.106e+11Hz -0.0248222 -0.0106855
+ 2.107e+11Hz -0.0248301 -0.010673
+ 2.108e+11Hz -0.0248382 -0.0106605
+ 2.109e+11Hz -0.0248464 -0.010648
+ 2.11e+11Hz -0.0248547 -0.0106356
+ 2.111e+11Hz -0.0248631 -0.0106232
+ 2.112e+11Hz -0.0248715 -0.0106109
+ 2.113e+11Hz -0.0248801 -0.0105985
+ 2.114e+11Hz -0.0248888 -0.0105862
+ 2.115e+11Hz -0.0248976 -0.0105739
+ 2.116e+11Hz -0.0249065 -0.0105616
+ 2.117e+11Hz -0.0249155 -0.0105494
+ 2.118e+11Hz -0.0249247 -0.0105372
+ 2.119e+11Hz -0.0249339 -0.0105249
+ 2.12e+11Hz -0.0249433 -0.0105127
+ 2.121e+11Hz -0.0249527 -0.0105005
+ 2.122e+11Hz -0.0249623 -0.0104883
+ 2.123e+11Hz -0.024972 -0.0104761
+ 2.124e+11Hz -0.0249819 -0.0104639
+ 2.125e+11Hz -0.0249918 -0.0104517
+ 2.126e+11Hz -0.0250019 -0.0104395
+ 2.127e+11Hz -0.0250121 -0.0104273
+ 2.128e+11Hz -0.0250225 -0.010415
+ 2.129e+11Hz -0.0250329 -0.0104028
+ 2.13e+11Hz -0.0250435 -0.0103905
+ 2.131e+11Hz -0.0250542 -0.0103783
+ 2.132e+11Hz -0.0250651 -0.010366
+ 2.133e+11Hz -0.025076 -0.0103536
+ 2.134e+11Hz -0.0250871 -0.0103413
+ 2.135e+11Hz -0.0250984 -0.0103289
+ 2.136e+11Hz -0.0251098 -0.0103165
+ 2.137e+11Hz -0.0251213 -0.010304
+ 2.138e+11Hz -0.0251329 -0.0102915
+ 2.139e+11Hz -0.0251447 -0.010279
+ 2.14e+11Hz -0.0251566 -0.0102664
+ 2.141e+11Hz -0.0251687 -0.0102538
+ 2.142e+11Hz -0.0251808 -0.0102411
+ 2.143e+11Hz -0.0251932 -0.0102283
+ 2.144e+11Hz -0.0252056 -0.0102155
+ 2.145e+11Hz -0.0252182 -0.0102026
+ 2.146e+11Hz -0.025231 -0.0101897
+ 2.147e+11Hz -0.0252438 -0.0101767
+ 2.148e+11Hz -0.0252569 -0.0101636
+ 2.149e+11Hz -0.02527 -0.0101504
+ 2.15e+11Hz -0.0252833 -0.0101372
+ 2.151e+11Hz -0.0252967 -0.0101239
+ 2.152e+11Hz -0.0253103 -0.0101105
+ 2.153e+11Hz -0.025324 -0.010097
+ 2.154e+11Hz -0.0253378 -0.0100834
+ 2.155e+11Hz -0.0253518 -0.0100697
+ 2.156e+11Hz -0.0253659 -0.0100559
+ 2.157e+11Hz -0.0253802 -0.010042
+ 2.158e+11Hz -0.0253946 -0.010028
+ 2.159e+11Hz -0.0254091 -0.0100139
+ 2.16e+11Hz -0.0254238 -0.00999965
+ 2.161e+11Hz -0.0254385 -0.0099853
+ 2.162e+11Hz -0.0254535 -0.00997083
+ 2.163e+11Hz -0.0254685 -0.00995624
+ 2.164e+11Hz -0.0254837 -0.00994151
+ 2.165e+11Hz -0.025499 -0.00992666
+ 2.166e+11Hz -0.0255145 -0.00991166
+ 2.167e+11Hz -0.02553 -0.00989653
+ 2.168e+11Hz -0.0255457 -0.00988125
+ 2.169e+11Hz -0.0255615 -0.00986583
+ 2.17e+11Hz -0.0255775 -0.00985026
+ 2.171e+11Hz -0.0255935 -0.00983453
+ 2.172e+11Hz -0.0256097 -0.00981864
+ 2.173e+11Hz -0.025626 -0.0098026
+ 2.174e+11Hz -0.0256424 -0.00978639
+ 2.175e+11Hz -0.025659 -0.00977001
+ 2.176e+11Hz -0.0256756 -0.00975347
+ 2.177e+11Hz -0.0256924 -0.00973675
+ 2.178e+11Hz -0.0257093 -0.00971985
+ 2.179e+11Hz -0.0257262 -0.00970276
+ 2.18e+11Hz -0.0257433 -0.0096855
+ 2.181e+11Hz -0.0257605 -0.00966805
+ 2.182e+11Hz -0.0257778 -0.0096504
+ 2.183e+11Hz -0.0257952 -0.00963256
+ 2.184e+11Hz -0.0258126 -0.00961452
+ 2.185e+11Hz -0.0258302 -0.00959629
+ 2.186e+11Hz -0.0258479 -0.00957785
+ 2.187e+11Hz -0.0258656 -0.0095592
+ 2.188e+11Hz -0.0258834 -0.00954034
+ 2.189e+11Hz -0.0259014 -0.00952126
+ 2.19e+11Hz -0.0259194 -0.00950197
+ 2.191e+11Hz -0.0259374 -0.00948247
+ 2.192e+11Hz -0.0259556 -0.00946273
+ 2.193e+11Hz -0.0259738 -0.00944278
+ 2.194e+11Hz -0.0259921 -0.00942259
+ 2.195e+11Hz -0.0260104 -0.00940218
+ 2.196e+11Hz -0.0260288 -0.00938153
+ 2.197e+11Hz -0.0260473 -0.00936064
+ 2.198e+11Hz -0.0260658 -0.00933951
+ 2.199e+11Hz -0.0260844 -0.00931815
+ 2.2e+11Hz -0.026103 -0.00929654
+ 2.201e+11Hz -0.0261217 -0.00927468
+ 2.202e+11Hz -0.0261404 -0.00925257
+ 2.203e+11Hz -0.0261591 -0.00923021
+ 2.204e+11Hz -0.0261779 -0.00920759
+ 2.205e+11Hz -0.0261967 -0.00918472
+ 2.206e+11Hz -0.0262156 -0.00916159
+ 2.207e+11Hz -0.0262344 -0.0091382
+ 2.208e+11Hz -0.0262533 -0.00911455
+ 2.209e+11Hz -0.0262722 -0.00909063
+ 2.21e+11Hz -0.0262911 -0.00906644
+ 2.211e+11Hz -0.0263099 -0.00904199
+ 2.212e+11Hz -0.0263288 -0.00901726
+ 2.213e+11Hz -0.0263477 -0.00899226
+ 2.214e+11Hz -0.0263666 -0.00896699
+ 2.215e+11Hz -0.0263855 -0.00894144
+ 2.216e+11Hz -0.0264044 -0.00891561
+ 2.217e+11Hz -0.0264232 -0.00888951
+ 2.218e+11Hz -0.026442 -0.00886312
+ 2.219e+11Hz -0.0264608 -0.00883645
+ 2.22e+11Hz -0.0264796 -0.0088095
+ 2.221e+11Hz -0.0264983 -0.00878227
+ 2.222e+11Hz -0.0265169 -0.00875475
+ 2.223e+11Hz -0.0265356 -0.00872694
+ 2.224e+11Hz -0.0265541 -0.00869884
+ 2.225e+11Hz -0.0265727 -0.00867046
+ 2.226e+11Hz -0.0265911 -0.00864179
+ 2.227e+11Hz -0.0266095 -0.00861283
+ 2.228e+11Hz -0.0266278 -0.00858358
+ 2.229e+11Hz -0.026646 -0.00855404
+ 2.23e+11Hz -0.0266642 -0.0085242
+ 2.231e+11Hz -0.0266823 -0.00849408
+ 2.232e+11Hz -0.0267003 -0.00846366
+ 2.233e+11Hz -0.0267181 -0.00843296
+ 2.234e+11Hz -0.0267359 -0.00840196
+ 2.235e+11Hz -0.0267536 -0.00837066
+ 2.236e+11Hz -0.0267712 -0.00833908
+ 2.237e+11Hz -0.0267886 -0.0083072
+ 2.238e+11Hz -0.026806 -0.00827504
+ 2.239e+11Hz -0.0268232 -0.00824258
+ 2.24e+11Hz -0.0268402 -0.00820983
+ 2.241e+11Hz -0.0268572 -0.00817679
+ 2.242e+11Hz -0.026874 -0.00814346
+ 2.243e+11Hz -0.0268906 -0.00810984
+ 2.244e+11Hz -0.0269071 -0.00807593
+ 2.245e+11Hz -0.0269235 -0.00804174
+ 2.246e+11Hz -0.0269397 -0.00800726
+ 2.247e+11Hz -0.0269557 -0.0079725
+ 2.248e+11Hz -0.0269716 -0.00793745
+ 2.249e+11Hz -0.0269872 -0.00790212
+ 2.25e+11Hz -0.0270027 -0.00786651
+ 2.251e+11Hz -0.027018 -0.00783062
+ 2.252e+11Hz -0.0270332 -0.00779445
+ 2.253e+11Hz -0.0270481 -0.007758
+ 2.254e+11Hz -0.0270628 -0.00772128
+ 2.255e+11Hz -0.0270773 -0.00768429
+ 2.256e+11Hz -0.0270917 -0.00764702
+ 2.257e+11Hz -0.0271058 -0.00760949
+ 2.258e+11Hz -0.0271196 -0.00757169
+ 2.259e+11Hz -0.0271333 -0.00753363
+ 2.26e+11Hz -0.0271467 -0.0074953
+ 2.261e+11Hz -0.0271599 -0.00745671
+ 2.262e+11Hz -0.0271729 -0.00741787
+ 2.263e+11Hz -0.0271856 -0.00737877
+ 2.264e+11Hz -0.0271981 -0.00733942
+ 2.265e+11Hz -0.0272103 -0.00729982
+ 2.266e+11Hz -0.0272222 -0.00725997
+ 2.267e+11Hz -0.0272339 -0.00721988
+ 2.268e+11Hz -0.0272453 -0.00717955
+ 2.269e+11Hz -0.0272565 -0.00713898
+ 2.27e+11Hz -0.0272674 -0.00709817
+ 2.271e+11Hz -0.027278 -0.00705714
+ 2.272e+11Hz -0.0272883 -0.00701587
+ 2.273e+11Hz -0.0272984 -0.00697438
+ 2.274e+11Hz -0.0273081 -0.00693267
+ 2.275e+11Hz -0.0273176 -0.00689075
+ 2.276e+11Hz -0.0273267 -0.00684861
+ 2.277e+11Hz -0.0273356 -0.00680626
+ 2.278e+11Hz -0.0273441 -0.0067637
+ 2.279e+11Hz -0.0273523 -0.00672094
+ 2.28e+11Hz -0.0273602 -0.00667798
+ 2.281e+11Hz -0.0273678 -0.00663483
+ 2.282e+11Hz -0.0273751 -0.00659148
+ 2.283e+11Hz -0.0273821 -0.00654795
+ 2.284e+11Hz -0.0273887 -0.00650424
+ 2.285e+11Hz -0.027395 -0.00646035
+ 2.286e+11Hz -0.0274009 -0.00641629
+ 2.287e+11Hz -0.0274065 -0.00637206
+ 2.288e+11Hz -0.0274118 -0.00632767
+ 2.289e+11Hz -0.0274167 -0.00628311
+ 2.29e+11Hz -0.0274213 -0.0062384
+ 2.291e+11Hz -0.0274255 -0.00619354
+ 2.292e+11Hz -0.0274294 -0.00614853
+ 2.293e+11Hz -0.0274329 -0.00610338
+ 2.294e+11Hz -0.0274361 -0.0060581
+ 2.295e+11Hz -0.0274388 -0.00601268
+ 2.296e+11Hz -0.0274413 -0.00596714
+ 2.297e+11Hz -0.0274433 -0.00592148
+ 2.298e+11Hz -0.027445 -0.0058757
+ 2.299e+11Hz -0.0274463 -0.00582981
+ 2.3e+11Hz -0.0274472 -0.00578382
+ 2.301e+11Hz -0.0274478 -0.00573772
+ 2.302e+11Hz -0.027448 -0.00569153
+ 2.303e+11Hz -0.0274478 -0.00564524
+ 2.304e+11Hz -0.0274472 -0.00559888
+ 2.305e+11Hz -0.0274462 -0.00555243
+ 2.306e+11Hz -0.0274449 -0.00550591
+ 2.307e+11Hz -0.0274431 -0.00545932
+ 2.308e+11Hz -0.027441 -0.00541266
+ 2.309e+11Hz -0.0274384 -0.00536595
+ 2.31e+11Hz -0.0274355 -0.00531919
+ 2.311e+11Hz -0.0274322 -0.00527237
+ 2.312e+11Hz -0.0274285 -0.00522552
+ 2.313e+11Hz -0.0274244 -0.00517863
+ 2.314e+11Hz -0.0274199 -0.00513171
+ 2.315e+11Hz -0.027415 -0.00508477
+ 2.316e+11Hz -0.0274097 -0.00503781
+ 2.317e+11Hz -0.027404 -0.00499083
+ 2.318e+11Hz -0.0273979 -0.00494384
+ 2.319e+11Hz -0.0273914 -0.00489686
+ 2.32e+11Hz -0.0273845 -0.00484988
+ 2.321e+11Hz -0.0273773 -0.0048029
+ 2.322e+11Hz -0.0273696 -0.00475594
+ 2.323e+11Hz -0.0273615 -0.004709
+ 2.324e+11Hz -0.027353 -0.00466209
+ 2.325e+11Hz -0.0273441 -0.00461521
+ 2.326e+11Hz -0.0273348 -0.00456836
+ 2.327e+11Hz -0.0273251 -0.00452156
+ 2.328e+11Hz -0.027315 -0.00447481
+ 2.329e+11Hz -0.0273045 -0.00442811
+ 2.33e+11Hz -0.0272936 -0.00438147
+ 2.331e+11Hz -0.0272824 -0.0043349
+ 2.332e+11Hz -0.0272707 -0.0042884
+ 2.333e+11Hz -0.0272586 -0.00424197
+ 2.334e+11Hz -0.0272461 -0.00419563
+ 2.335e+11Hz -0.0272333 -0.00414937
+ 2.336e+11Hz -0.02722 -0.00410321
+ 2.337e+11Hz -0.0272064 -0.00405715
+ 2.338e+11Hz -0.0271923 -0.00401119
+ 2.339e+11Hz -0.0271779 -0.00396534
+ 2.34e+11Hz -0.0271631 -0.0039196
+ 2.341e+11Hz -0.0271479 -0.00387399
+ 2.342e+11Hz -0.0271324 -0.0038285
+ 2.343e+11Hz -0.0271164 -0.00378314
+ 2.344e+11Hz -0.0271001 -0.00373791
+ 2.345e+11Hz -0.0270834 -0.00369283
+ 2.346e+11Hz -0.0270663 -0.00364789
+ 2.347e+11Hz -0.0270489 -0.00360311
+ 2.348e+11Hz -0.027031 -0.00355848
+ 2.349e+11Hz -0.0270129 -0.00351401
+ 2.35e+11Hz -0.0269943 -0.00346971
+ 2.351e+11Hz -0.0269754 -0.00342559
+ 2.352e+11Hz -0.0269561 -0.00338163
+ 2.353e+11Hz -0.0269365 -0.00333786
+ 2.354e+11Hz -0.0269165 -0.00329428
+ 2.355e+11Hz -0.0268962 -0.00325088
+ 2.356e+11Hz -0.0268755 -0.00320768
+ 2.357e+11Hz -0.0268545 -0.00316468
+ 2.358e+11Hz -0.0268331 -0.00312188
+ 2.359e+11Hz -0.0268114 -0.0030793
+ 2.36e+11Hz -0.0267894 -0.00303692
+ 2.361e+11Hz -0.026767 -0.00299476
+ 2.362e+11Hz -0.0267443 -0.00295283
+ 2.363e+11Hz -0.0267213 -0.00291112
+ 2.364e+11Hz -0.026698 -0.00286964
+ 2.365e+11Hz -0.0266743 -0.00282839
+ 2.366e+11Hz -0.0266503 -0.00278739
+ 2.367e+11Hz -0.0266261 -0.00274662
+ 2.368e+11Hz -0.0266015 -0.0027061
+ 2.369e+11Hz -0.0265766 -0.00266583
+ 2.37e+11Hz -0.0265514 -0.00262581
+ 2.371e+11Hz -0.0265259 -0.00258605
+ 2.372e+11Hz -0.0265002 -0.00254655
+ 2.373e+11Hz -0.0264741 -0.00250732
+ 2.374e+11Hz -0.0264478 -0.00246835
+ 2.375e+11Hz -0.0264212 -0.00242965
+ 2.376e+11Hz -0.0263943 -0.00239123
+ 2.377e+11Hz -0.0263671 -0.00235308
+ 2.378e+11Hz -0.0263397 -0.00231521
+ 2.379e+11Hz -0.026312 -0.00227762
+ 2.38e+11Hz -0.0262841 -0.00224033
+ 2.381e+11Hz -0.0262559 -0.00220331
+ 2.382e+11Hz -0.0262275 -0.00216659
+ 2.383e+11Hz -0.0261988 -0.00213017
+ 2.384e+11Hz -0.0261699 -0.00209404
+ 2.385e+11Hz -0.0261408 -0.00205821
+ 2.386e+11Hz -0.0261114 -0.00202268
+ 2.387e+11Hz -0.0260818 -0.00198746
+ 2.388e+11Hz -0.026052 -0.00195254
+ 2.389e+11Hz -0.0260219 -0.00191792
+ 2.39e+11Hz -0.0259917 -0.00188362
+ 2.391e+11Hz -0.0259613 -0.00184963
+ 2.392e+11Hz -0.0259306 -0.00181595
+ 2.393e+11Hz -0.0258998 -0.00178259
+ 2.394e+11Hz -0.0258687 -0.00174955
+ 2.395e+11Hz -0.0258375 -0.00171682
+ 2.396e+11Hz -0.0258061 -0.00168442
+ 2.397e+11Hz -0.0257746 -0.00165234
+ 2.398e+11Hz -0.0257428 -0.00162058
+ 2.399e+11Hz -0.0257109 -0.00158914
+ 2.4e+11Hz -0.0256788 -0.00155803
+ 2.401e+11Hz -0.0256466 -0.00152724
+ 2.402e+11Hz -0.0256142 -0.00149679
+ 2.403e+11Hz -0.0255817 -0.00146666
+ 2.404e+11Hz -0.025549 -0.00143686
+ 2.405e+11Hz -0.0255162 -0.00140739
+ 2.406e+11Hz -0.0254833 -0.00137825
+ 2.407e+11Hz -0.0254502 -0.00134944
+ 2.408e+11Hz -0.025417 -0.00132096
+ 2.409e+11Hz -0.0253837 -0.00129281
+ 2.41e+11Hz -0.0253503 -0.001265
+ 2.411e+11Hz -0.0253168 -0.00123752
+ 2.412e+11Hz -0.0252831 -0.00121037
+ 2.413e+11Hz -0.0252494 -0.00118355
+ 2.414e+11Hz -0.0252156 -0.00115707
+ 2.415e+11Hz -0.0251817 -0.00113092
+ 2.416e+11Hz -0.0251477 -0.0011051
+ 2.417e+11Hz -0.0251136 -0.00107961
+ 2.418e+11Hz -0.0250794 -0.00105445
+ 2.419e+11Hz -0.0250452 -0.00102962
+ 2.42e+11Hz -0.0250109 -0.00100513
+ 2.421e+11Hz -0.0249766 -0.000980965
+ 2.422e+11Hz -0.0249422 -0.000957129
+ 2.423e+11Hz -0.0249077 -0.000933622
+ 2.424e+11Hz -0.0248732 -0.000910443
+ 2.425e+11Hz -0.0248386 -0.00088759
+ 2.426e+11Hz -0.024804 -0.000865064
+ 2.427e+11Hz -0.0247694 -0.000842863
+ 2.428e+11Hz -0.0247347 -0.000820986
+ 2.429e+11Hz -0.0247001 -0.000799432
+ 2.43e+11Hz -0.0246653 -0.000778199
+ 2.431e+11Hz -0.0246306 -0.000757287
+ 2.432e+11Hz -0.0245959 -0.000736694
+ 2.433e+11Hz -0.0245611 -0.000716418
+ 2.434e+11Hz -0.0245264 -0.000696459
+ 2.435e+11Hz -0.0244916 -0.000676815
+ 2.436e+11Hz -0.0244568 -0.000657484
+ 2.437e+11Hz -0.0244221 -0.000638464
+ 2.438e+11Hz -0.0243873 -0.000619755
+ 2.439e+11Hz -0.0243526 -0.000601353
+ 2.44e+11Hz -0.0243179 -0.000583258
+ 2.441e+11Hz -0.0242832 -0.000565468
+ 2.442e+11Hz -0.0242485 -0.000547981
+ 2.443e+11Hz -0.0242139 -0.000530794
+ 2.444e+11Hz -0.0241793 -0.000513906
+ 2.445e+11Hz -0.0241447 -0.000497316
+ 2.446e+11Hz -0.0241101 -0.00048102
+ 2.447e+11Hz -0.0240756 -0.000465017
+ 2.448e+11Hz -0.0240412 -0.000449304
+ 2.449e+11Hz -0.0240068 -0.00043388
+ 2.45e+11Hz -0.0239724 -0.000418742
+ 2.451e+11Hz -0.0239381 -0.000403888
+ 2.452e+11Hz -0.0239039 -0.000389316
+ 2.453e+11Hz -0.0238697 -0.000375023
+ 2.454e+11Hz -0.0238356 -0.000361008
+ 2.455e+11Hz -0.0238015 -0.000347267
+ 2.456e+11Hz -0.0237676 -0.000333798
+ 2.457e+11Hz -0.0237337 -0.0003206
+ 2.458e+11Hz -0.0236998 -0.000307669
+ 2.459e+11Hz -0.0236661 -0.000295002
+ 2.46e+11Hz -0.0236324 -0.000282599
+ 2.461e+11Hz -0.0235988 -0.000270455
+ 2.462e+11Hz -0.0235653 -0.000258569
+ 2.463e+11Hz -0.0235319 -0.000246937
+ 2.464e+11Hz -0.0234985 -0.000235558
+ 2.465e+11Hz -0.0234653 -0.000224429
+ 2.466e+11Hz -0.0234321 -0.000213547
+ 2.467e+11Hz -0.0233991 -0.000202909
+ 2.468e+11Hz -0.0233662 -0.000192513
+ 2.469e+11Hz -0.0233333 -0.000182357
+ 2.47e+11Hz -0.0233006 -0.000172437
+ 2.471e+11Hz -0.0232679 -0.000162751
+ 2.472e+11Hz -0.0232354 -0.000153296
+ 2.473e+11Hz -0.023203 -0.00014407
+ 2.474e+11Hz -0.0231706 -0.00013507
+ 2.475e+11Hz -0.0231384 -0.000126293
+ 2.476e+11Hz -0.0231063 -0.000117737
+ 2.477e+11Hz -0.0230744 -0.000109399
+ 2.478e+11Hz -0.0230425 -0.000101277
+ 2.479e+11Hz -0.0230108 -9.33669e-05
+ 2.48e+11Hz -0.0229792 -8.5667e-05
+ 2.481e+11Hz -0.0229477 -7.81745e-05
+ 2.482e+11Hz -0.0229163 -7.08868e-05
+ 2.483e+11Hz -0.022885 -6.38012e-05
+ 2.484e+11Hz -0.0228539 -5.6915e-05
+ 2.485e+11Hz -0.0228229 -5.02257e-05
+ 2.486e+11Hz -0.0227921 -4.37307e-05
+ 2.487e+11Hz -0.0227613 -3.74273e-05
+ 2.488e+11Hz -0.0227307 -3.13131e-05
+ 2.489e+11Hz -0.0227002 -2.53853e-05
+ 2.49e+11Hz -0.0226699 -1.96415e-05
+ 2.491e+11Hz -0.0226397 -1.4079e-05
+ 2.492e+11Hz -0.0226096 -8.69551e-06
+ 2.493e+11Hz -0.0225796 -3.48836e-06
+ 2.494e+11Hz -0.0225498 1.5449e-06
+ 2.495e+11Hz -0.0225202 6.40676e-06
+ 2.496e+11Hz -0.0224906 1.10997e-05
+ 2.497e+11Hz -0.0224612 1.5626e-05
+ 2.498e+11Hz -0.022432 1.99883e-05
+ 2.499e+11Hz -0.0224029 2.41889e-05
+ 2.5e+11Hz -0.0223739 2.82301e-05
+ 2.501e+11Hz -0.022345 3.21144e-05
+ 2.502e+11Hz -0.0223163 3.5844e-05
+ 2.503e+11Hz -0.0222878 3.94213e-05
+ 2.504e+11Hz -0.0222594 4.28485e-05
+ 2.505e+11Hz -0.0222311 4.61279e-05
+ 2.506e+11Hz -0.022203 4.92618e-05
+ 2.507e+11Hz -0.022175 5.22523e-05
+ 2.508e+11Hz -0.0221471 5.51017e-05
+ 2.509e+11Hz -0.0221194 5.78121e-05
+ 2.51e+11Hz -0.0220919 6.03856e-05
+ 2.511e+11Hz -0.0220645 6.28245e-05
+ 2.512e+11Hz -0.0220372 6.51306e-05
+ 2.513e+11Hz -0.0220101 6.73063e-05
+ 2.514e+11Hz -0.0219831 6.93533e-05
+ 2.515e+11Hz -0.0219563 7.12739e-05
+ 2.516e+11Hz -0.0219296 7.307e-05
+ 2.517e+11Hz -0.0219031 7.47435e-05
+ 2.518e+11Hz -0.0218767 7.62963e-05
+ 2.519e+11Hz -0.0218505 7.77305e-05
+ 2.52e+11Hz -0.0218244 7.90478e-05
+ 2.521e+11Hz -0.0217984 8.02503e-05
+ 2.522e+11Hz -0.0217726 8.13396e-05
+ 2.523e+11Hz -0.021747 8.23176e-05
+ 2.524e+11Hz -0.0217215 8.31861e-05
+ 2.525e+11Hz -0.0216961 8.39469e-05
+ 2.526e+11Hz -0.0216709 8.46017e-05
+ 2.527e+11Hz -0.0216458 8.51522e-05
+ 2.528e+11Hz -0.0216209 8.56002e-05
+ 2.529e+11Hz -0.0215961 8.59473e-05
+ 2.53e+11Hz -0.0215715 8.61952e-05
+ 2.531e+11Hz -0.021547 8.63456e-05
+ 2.532e+11Hz -0.0215227 8.63999e-05
+ 2.533e+11Hz -0.0214985 8.63598e-05
+ 2.534e+11Hz -0.0214745 8.6227e-05
+ 2.535e+11Hz -0.0214506 8.60029e-05
+ 2.536e+11Hz -0.0214269 8.56891e-05
+ 2.537e+11Hz -0.0214033 8.52871e-05
+ 2.538e+11Hz -0.0213798 8.47985e-05
+ 2.539e+11Hz -0.0213565 8.42246e-05
+ 2.54e+11Hz -0.0213334 8.3567e-05
+ 2.541e+11Hz -0.0213104 8.28271e-05
+ 2.542e+11Hz -0.0212875 8.20064e-05
+ 2.543e+11Hz -0.0212648 8.11063e-05
+ 2.544e+11Hz -0.0212423 8.01282e-05
+ 2.545e+11Hz -0.0212199 7.90735e-05
+ 2.546e+11Hz -0.0211976 7.79437e-05
+ 2.547e+11Hz -0.0211755 7.674e-05
+ 2.548e+11Hz -0.0211536 7.54639e-05
+ 2.549e+11Hz -0.0211318 7.41168e-05
+ 2.55e+11Hz -0.0211101 7.26999e-05
+ 2.551e+11Hz -0.0210886 7.12146e-05
+ 2.552e+11Hz -0.0210673 6.96624e-05
+ 2.553e+11Hz -0.0210461 6.80445e-05
+ 2.554e+11Hz -0.021025 6.63622e-05
+ 2.555e+11Hz -0.0210041 6.4617e-05
+ 2.556e+11Hz -0.0209833 6.28101e-05
+ 2.557e+11Hz -0.0209627 6.09428e-05
+ 2.558e+11Hz -0.0209423 5.90166e-05
+ 2.559e+11Hz -0.020922 5.70326e-05
+ 2.56e+11Hz -0.0209018 5.49924e-05
+ 2.561e+11Hz -0.0208818 5.28972e-05
+ 2.562e+11Hz -0.020862 5.07483e-05
+ 2.563e+11Hz -0.0208423 4.85471e-05
+ 2.564e+11Hz -0.0208228 4.62949e-05
+ 2.565e+11Hz -0.0208034 4.39932e-05
+ 2.566e+11Hz -0.0207841 4.16432e-05
+ 2.567e+11Hz -0.0207651 3.92464e-05
+ 2.568e+11Hz -0.0207461 3.68041e-05
+ 2.569e+11Hz -0.0207274 3.43178e-05
+ 2.57e+11Hz -0.0207088 3.17889e-05
+ 2.571e+11Hz -0.0206903 2.92187e-05
+ 2.572e+11Hz -0.020672 2.66087e-05
+ 2.573e+11Hz -0.0206538 2.39604e-05
+ 2.574e+11Hz -0.0206359 2.12753e-05
+ 2.575e+11Hz -0.020618 1.85547e-05
+ 2.576e+11Hz -0.0206004 1.58003e-05
+ 2.577e+11Hz -0.0205828 1.30135e-05
+ 2.578e+11Hz -0.0205655 1.0196e-05
+ 2.579e+11Hz -0.0205483 7.34912e-06
+ 2.58e+11Hz -0.0205312 4.47462e-06
+ 2.581e+11Hz -0.0205144 1.57405e-06
+ 2.582e+11Hz -0.0204976 -1.35096e-06
+ 2.583e+11Hz -0.0204811 -4.29876e-06
+ 2.584e+11Hz -0.0204647 -7.26767e-06
+ 2.585e+11Hz -0.0204485 -1.0256e-05
+ 2.586e+11Hz -0.0204324 -1.3262e-05
+ 2.587e+11Hz -0.0204165 -1.6284e-05
+ 2.588e+11Hz -0.0204007 -1.93201e-05
+ 2.589e+11Hz -0.0203852 -2.23686e-05
+ 2.59e+11Hz -0.0203697 -2.54275e-05
+ 2.591e+11Hz -0.0203545 -2.84952e-05
+ 2.592e+11Hz -0.0203394 -3.15696e-05
+ 2.593e+11Hz -0.0203245 -3.46488e-05
+ 2.594e+11Hz -0.0203097 -3.77309e-05
+ 2.595e+11Hz -0.0202951 -4.08139e-05
+ 2.596e+11Hz -0.0202807 -4.38958e-05
+ 2.597e+11Hz -0.0202665 -4.69745e-05
+ 2.598e+11Hz -0.0202524 -5.00479e-05
+ 2.599e+11Hz -0.0202385 -5.3114e-05
+ 2.6e+11Hz -0.0202247 -5.61705e-05
+ 2.601e+11Hz -0.0202112 -5.92153e-05
+ 2.602e+11Hz -0.0201977 -6.22462e-05
+ 2.603e+11Hz -0.0201845 -6.5261e-05
+ 2.604e+11Hz -0.0201714 -6.82573e-05
+ 2.605e+11Hz -0.0201585 -7.12328e-05
+ 2.606e+11Hz -0.0201458 -7.41852e-05
+ 2.607e+11Hz -0.0201333 -7.71121e-05
+ 2.608e+11Hz -0.0201209 -8.00111e-05
+ 2.609e+11Hz -0.0201087 -8.28796e-05
+ 2.61e+11Hz -0.0200966 -8.57153e-05
+ 2.611e+11Hz -0.0200848 -8.85157e-05
+ 2.612e+11Hz -0.0200731 -9.1278e-05
+ 2.613e+11Hz -0.0200616 -9.39998e-05
+ 2.614e+11Hz -0.0200502 -9.66785e-05
+ 2.615e+11Hz -0.020039 -9.93113e-05
+ 2.616e+11Hz -0.020028 -0.000101896
+ 2.617e+11Hz -0.0200172 -0.000104429
+ 2.618e+11Hz -0.0200065 -0.000106908
+ 2.619e+11Hz -0.019996 -0.00010933
+ 2.62e+11Hz -0.0199857 -0.000111693
+ 2.621e+11Hz -0.0199756 -0.000113993
+ 2.622e+11Hz -0.0199656 -0.000116228
+ 2.623e+11Hz -0.0199558 -0.000118394
+ 2.624e+11Hz -0.0199462 -0.00012049
+ 2.625e+11Hz -0.0199367 -0.000122511
+ 2.626e+11Hz -0.0199274 -0.000124455
+ 2.627e+11Hz -0.0199183 -0.000126319
+ 2.628e+11Hz -0.0199094 -0.0001281
+ 2.629e+11Hz -0.0199006 -0.000129794
+ 2.63e+11Hz -0.019892 -0.000131399
+ 2.631e+11Hz -0.0198835 -0.000132912
+ 2.632e+11Hz -0.0198753 -0.000134329
+ 2.633e+11Hz -0.0198672 -0.000135647
+ 2.634e+11Hz -0.0198592 -0.000136863
+ 2.635e+11Hz -0.0198514 -0.000137973
+ 2.636e+11Hz -0.0198438 -0.000138976
+ 2.637e+11Hz -0.0198364 -0.000139866
+ 2.638e+11Hz -0.0198291 -0.000140642
+ 2.639e+11Hz -0.0198219 -0.0001413
+ 2.64e+11Hz -0.0198149 -0.000141836
+ 2.641e+11Hz -0.0198081 -0.000142247
+ 2.642e+11Hz -0.0198015 -0.00014253
+ 2.643e+11Hz -0.019795 -0.000142682
+ 2.644e+11Hz -0.0197886 -0.000142699
+ 2.645e+11Hz -0.0197824 -0.000142578
+ 2.646e+11Hz -0.0197764 -0.000142315
+ 2.647e+11Hz -0.0197705 -0.000141908
+ 2.648e+11Hz -0.0197647 -0.000141353
+ 2.649e+11Hz -0.0197591 -0.000140646
+ 2.65e+11Hz -0.0197536 -0.000139785
+ 2.651e+11Hz -0.0197483 -0.000138766
+ 2.652e+11Hz -0.0197431 -0.000137585
+ 2.653e+11Hz -0.0197381 -0.00013624
+ 2.654e+11Hz -0.0197332 -0.000134726
+ 2.655e+11Hz -0.0197284 -0.000133042
+ 2.656e+11Hz -0.0197237 -0.000131182
+ 2.657e+11Hz -0.0197192 -0.000129145
+ 2.658e+11Hz -0.0197148 -0.000126927
+ 2.659e+11Hz -0.0197105 -0.000124524
+ 2.66e+11Hz -0.0197064 -0.000121934
+ 2.661e+11Hz -0.0197023 -0.000119153
+ 2.662e+11Hz -0.0196984 -0.000116178
+ 2.663e+11Hz -0.0196946 -0.000113006
+ 2.664e+11Hz -0.0196909 -0.000109633
+ 2.665e+11Hz -0.0196873 -0.000106058
+ 2.666e+11Hz -0.0196838 -0.000102276
+ 2.667e+11Hz -0.0196804 -9.82843e-05
+ 2.668e+11Hz -0.0196771 -9.40805e-05
+ 2.669e+11Hz -0.0196739 -8.96614e-05
+ 2.67e+11Hz -0.0196708 -8.5024e-05
+ 2.671e+11Hz -0.0196678 -8.01655e-05
+ 2.672e+11Hz -0.0196648 -7.5083e-05
+ 2.673e+11Hz -0.019662 -6.97738e-05
+ 2.674e+11Hz -0.0196592 -6.42351e-05
+ 2.675e+11Hz -0.0196564 -5.84643e-05
+ 2.676e+11Hz -0.0196538 -5.24586e-05
+ 2.677e+11Hz -0.0196512 -4.62156e-05
+ 2.678e+11Hz -0.0196486 -3.97327e-05
+ 2.679e+11Hz -0.0196462 -3.30074e-05
+ 2.68e+11Hz -0.0196437 -2.60373e-05
+ 2.681e+11Hz -0.0196413 -1.88202e-05
+ 2.682e+11Hz -0.019639 -1.13536e-05
+ 2.683e+11Hz -0.0196367 -3.63541e-06
+ 2.684e+11Hz -0.0196344 4.33653e-06
+ 2.685e+11Hz -0.0196322 1.25643e-05
+ 2.686e+11Hz -0.01963 2.10499e-05
+ 2.687e+11Hz -0.0196278 2.97953e-05
+ 2.688e+11Hz -0.0196256 3.88023e-05
+ 2.689e+11Hz -0.0196234 4.80727e-05
+ 2.69e+11Hz -0.0196212 5.76082e-05
+ 2.691e+11Hz -0.0196191 6.74105e-05
+ 2.692e+11Hz -0.0196169 7.74809e-05
+ 2.693e+11Hz -0.0196147 8.78211e-05
+ 2.694e+11Hz -0.0196125 9.84323e-05
+ 2.695e+11Hz -0.0196103 0.000109316
+ 2.696e+11Hz -0.019608 0.000120473
+ 2.697e+11Hz -0.0196058 0.000131905
+ 2.698e+11Hz -0.0196035 0.000143612
+ 2.699e+11Hz -0.0196011 0.000155596
+ 2.7e+11Hz -0.0195987 0.000167857
+ 2.701e+11Hz -0.0195962 0.000180396
+ 2.702e+11Hz -0.0195937 0.000193214
+ 2.703e+11Hz -0.0195912 0.00020631
+ 2.704e+11Hz -0.0195885 0.000219687
+ 2.705e+11Hz -0.0195858 0.000233343
+ 2.706e+11Hz -0.019583 0.000247279
+ 2.707e+11Hz -0.0195801 0.000261495
+ 2.708e+11Hz -0.0195771 0.000275991
+ 2.709e+11Hz -0.0195741 0.000290768
+ 2.71e+11Hz -0.0195709 0.000305823
+ 2.711e+11Hz -0.0195676 0.000321159
+ 2.712e+11Hz -0.0195642 0.000336773
+ 2.713e+11Hz -0.0195607 0.000352665
+ 2.714e+11Hz -0.019557 0.000368835
+ 2.715e+11Hz -0.0195532 0.000385281
+ 2.716e+11Hz -0.0195493 0.000402004
+ 2.717e+11Hz -0.0195453 0.000419001
+ 2.718e+11Hz -0.019541 0.000436272
+ 2.719e+11Hz -0.0195367 0.000453815
+ 2.72e+11Hz -0.0195321 0.000471629
+ 2.721e+11Hz -0.0195274 0.000489712
+ 2.722e+11Hz -0.0195226 0.000508063
+ 2.723e+11Hz -0.0195175 0.00052668
+ 2.724e+11Hz -0.0195123 0.000545561
+ 2.725e+11Hz -0.0195069 0.000564704
+ 2.726e+11Hz -0.0195012 0.000584106
+ 2.727e+11Hz -0.0194954 0.000603767
+ 2.728e+11Hz -0.0194894 0.000623682
+ 2.729e+11Hz -0.0194831 0.000643851
+ 2.73e+11Hz -0.0194766 0.000664269
+ 2.731e+11Hz -0.0194699 0.000684935
+ 2.732e+11Hz -0.019463 0.000705845
+ 2.733e+11Hz -0.0194558 0.000726996
+ 2.734e+11Hz -0.0194484 0.000748386
+ 2.735e+11Hz -0.0194408 0.000770011
+ 2.736e+11Hz -0.0194329 0.000791868
+ 2.737e+11Hz -0.0194247 0.000813953
+ 2.738e+11Hz -0.0194162 0.000836262
+ 2.739e+11Hz -0.0194075 0.000858792
+ 2.74e+11Hz -0.0193985 0.000881539
+ 2.741e+11Hz -0.0193893 0.000904499
+ 2.742e+11Hz -0.0193797 0.000927668
+ 2.743e+11Hz -0.0193699 0.000951042
+ 2.744e+11Hz -0.0193597 0.000974616
+ 2.745e+11Hz -0.0193493 0.000998386
+ 2.746e+11Hz -0.0193385 0.00102235
+ 2.747e+11Hz -0.0193275 0.0010465
+ 2.748e+11Hz -0.0193161 0.00107083
+ 2.749e+11Hz -0.0193044 0.00109533
+ 2.75e+11Hz -0.0192923 0.00112001
+ 2.751e+11Hz -0.01928 0.00114486
+ 2.752e+11Hz -0.0192673 0.00116986
+ 2.753e+11Hz -0.0192542 0.00119503
+ 2.754e+11Hz -0.0192409 0.00122034
+ 2.755e+11Hz -0.0192271 0.0012458
+ 2.756e+11Hz -0.019213 0.0012714
+ 2.757e+11Hz -0.0191986 0.00129713
+ 2.758e+11Hz -0.0191838 0.00132299
+ 2.759e+11Hz -0.0191686 0.00134898
+ 2.76e+11Hz -0.0191531 0.00137508
+ 2.761e+11Hz -0.0191372 0.00140129
+ 2.762e+11Hz -0.0191209 0.0014276
+ 2.763e+11Hz -0.0191042 0.00145401
+ 2.764e+11Hz -0.0190872 0.00148051
+ 2.765e+11Hz -0.0190698 0.0015071
+ 2.766e+11Hz -0.0190519 0.00153376
+ 2.767e+11Hz -0.0190337 0.0015605
+ 2.768e+11Hz -0.0190151 0.0015873
+ 2.769e+11Hz -0.0189961 0.00161415
+ 2.77e+11Hz -0.0189767 0.00164106
+ 2.771e+11Hz -0.0189569 0.00166802
+ 2.772e+11Hz -0.0189367 0.001695
+ 2.773e+11Hz -0.0189161 0.00172202
+ 2.774e+11Hz -0.018895 0.00174907
+ 2.775e+11Hz -0.0188736 0.00177613
+ 2.776e+11Hz -0.0188518 0.00180319
+ 2.777e+11Hz -0.0188295 0.00183026
+ 2.778e+11Hz -0.0188068 0.00185732
+ 2.779e+11Hz -0.0187837 0.00188437
+ 2.78e+11Hz -0.0187602 0.0019114
+ 2.781e+11Hz -0.0187363 0.0019384
+ 2.782e+11Hz -0.0187119 0.00196536
+ 2.783e+11Hz -0.0186871 0.00199228
+ 2.784e+11Hz -0.0186619 0.00201915
+ 2.785e+11Hz -0.0186363 0.00204596
+ 2.786e+11Hz -0.0186103 0.0020727
+ 2.787e+11Hz -0.0185838 0.00209937
+ 2.788e+11Hz -0.0185569 0.00212596
+ 2.789e+11Hz -0.0185296 0.00215246
+ 2.79e+11Hz -0.0185019 0.00217886
+ 2.791e+11Hz -0.0184737 0.00220516
+ 2.792e+11Hz -0.0184451 0.00223134
+ 2.793e+11Hz -0.0184161 0.00225741
+ 2.794e+11Hz -0.0183867 0.00228334
+ 2.795e+11Hz -0.0183569 0.00230914
+ 2.796e+11Hz -0.0183266 0.0023348
+ 2.797e+11Hz -0.018296 0.00236031
+ 2.798e+11Hz -0.0182649 0.00238565
+ 2.799e+11Hz -0.0182334 0.00241084
+ 2.8e+11Hz -0.0182015 0.00243584
+ 2.801e+11Hz -0.0181691 0.00246067
+ 2.802e+11Hz -0.0181364 0.0024853
+ 2.803e+11Hz -0.0181033 0.00250974
+ 2.804e+11Hz -0.0180698 0.00253398
+ 2.805e+11Hz -0.0180358 0.002558
+ 2.806e+11Hz -0.0180015 0.00258181
+ 2.807e+11Hz -0.0179668 0.00260538
+ 2.808e+11Hz -0.0179317 0.00262873
+ 2.809e+11Hz -0.0178962 0.00265183
+ 2.81e+11Hz -0.0178603 0.00267468
+ 2.811e+11Hz -0.017824 0.00269728
+ 2.812e+11Hz -0.0177874 0.00271962
+ 2.813e+11Hz -0.0177504 0.00274168
+ 2.814e+11Hz -0.017713 0.00276347
+ 2.815e+11Hz -0.0176752 0.00278497
+ 2.816e+11Hz -0.0176371 0.00280619
+ 2.817e+11Hz -0.0175986 0.0028271
+ 2.818e+11Hz -0.0175598 0.00284772
+ 2.819e+11Hz -0.0175207 0.00286802
+ 2.82e+11Hz -0.0174811 0.002888
+ 2.821e+11Hz -0.0174413 0.00290766
+ 2.822e+11Hz -0.0174011 0.00292699
+ 2.823e+11Hz -0.0173606 0.00294599
+ 2.824e+11Hz -0.0173198 0.00296464
+ 2.825e+11Hz -0.0172786 0.00298294
+ 2.826e+11Hz -0.0172372 0.00300089
+ 2.827e+11Hz -0.0171954 0.00301848
+ 2.828e+11Hz -0.0171533 0.0030357
+ 2.829e+11Hz -0.017111 0.00305255
+ 2.83e+11Hz -0.0170683 0.00306903
+ 2.831e+11Hz -0.0170254 0.00308512
+ 2.832e+11Hz -0.0169822 0.00310083
+ 2.833e+11Hz -0.0169388 0.00311614
+ 2.834e+11Hz -0.016895 0.00313105
+ 2.835e+11Hz -0.016851 0.00314556
+ 2.836e+11Hz -0.0168068 0.00315967
+ 2.837e+11Hz -0.0167623 0.00317336
+ 2.838e+11Hz -0.0167176 0.00318664
+ 2.839e+11Hz -0.0166727 0.0031995
+ 2.84e+11Hz -0.0166275 0.00321193
+ 2.841e+11Hz -0.0165821 0.00322393
+ 2.842e+11Hz -0.0165366 0.0032355
+ 2.843e+11Hz -0.0164908 0.00324664
+ 2.844e+11Hz -0.0164448 0.00325733
+ 2.845e+11Hz -0.0163986 0.00326758
+ 2.846e+11Hz -0.0163523 0.00327739
+ 2.847e+11Hz -0.0163058 0.00328674
+ 2.848e+11Hz -0.0162591 0.00329564
+ 2.849e+11Hz -0.0162123 0.00330409
+ 2.85e+11Hz -0.0161653 0.00331208
+ 2.851e+11Hz -0.0161182 0.00331961
+ 2.852e+11Hz -0.016071 0.00332667
+ 2.853e+11Hz -0.0160236 0.00333327
+ 2.854e+11Hz -0.0159762 0.0033394
+ 2.855e+11Hz -0.0159286 0.00334506
+ 2.856e+11Hz -0.0158809 0.00335025
+ 2.857e+11Hz -0.0158331 0.00335497
+ 2.858e+11Hz -0.0157853 0.00335922
+ 2.859e+11Hz -0.0157373 0.00336299
+ 2.86e+11Hz -0.0156893 0.00336628
+ 2.861e+11Hz -0.0156413 0.0033691
+ 2.862e+11Hz -0.0155932 0.00337144
+ 2.863e+11Hz -0.015545 0.0033733
+ 2.864e+11Hz -0.0154969 0.00337469
+ 2.865e+11Hz -0.0154487 0.00337559
+ 2.866e+11Hz -0.0154004 0.00337602
+ 2.867e+11Hz -0.0153522 0.00337596
+ 2.868e+11Hz -0.015304 0.00337543
+ 2.869e+11Hz -0.0152558 0.00337442
+ 2.87e+11Hz -0.0152075 0.00337293
+ 2.871e+11Hz -0.0151594 0.00337097
+ 2.872e+11Hz -0.0151112 0.00336853
+ 2.873e+11Hz -0.0150631 0.00336562
+ 2.874e+11Hz -0.015015 0.00336223
+ 2.875e+11Hz -0.014967 0.00335837
+ 2.876e+11Hz -0.014919 0.00335404
+ 2.877e+11Hz -0.0148712 0.00334925
+ 2.878e+11Hz -0.0148234 0.00334398
+ 2.879e+11Hz -0.0147756 0.00333825
+ 2.88e+11Hz -0.014728 0.00333206
+ 2.881e+11Hz -0.0146805 0.00332541
+ 2.882e+11Hz -0.0146331 0.0033183
+ 2.883e+11Hz -0.0145858 0.00331074
+ 2.884e+11Hz -0.0145386 0.00330273
+ 2.885e+11Hz -0.0144916 0.00329427
+ 2.886e+11Hz -0.0144447 0.00328536
+ 2.887e+11Hz -0.014398 0.003276
+ 2.888e+11Hz -0.0143514 0.00326621
+ 2.889e+11Hz -0.0143049 0.00325599
+ 2.89e+11Hz -0.0142587 0.00324533
+ 2.891e+11Hz -0.0142126 0.00323425
+ 2.892e+11Hz -0.0141666 0.00322274
+ 2.893e+11Hz -0.0141209 0.00321081
+ 2.894e+11Hz -0.0140754 0.00319846
+ 2.895e+11Hz -0.0140301 0.0031857
+ 2.896e+11Hz -0.0139849 0.00317254
+ 2.897e+11Hz -0.01394 0.00315898
+ 2.898e+11Hz -0.0138954 0.00314501
+ 2.899e+11Hz -0.0138509 0.00313066
+ 2.9e+11Hz -0.0138067 0.00311591
+ 2.901e+11Hz -0.0137627 0.00310079
+ 2.902e+11Hz -0.0137189 0.00308528
+ 2.903e+11Hz -0.0136754 0.0030694
+ 2.904e+11Hz -0.0136322 0.00305316
+ 2.905e+11Hz -0.0135892 0.00303656
+ 2.906e+11Hz -0.0135465 0.00301959
+ 2.907e+11Hz -0.0135041 0.00300228
+ 2.908e+11Hz -0.0134619 0.00298463
+ 2.909e+11Hz -0.01342 0.00296663
+ 2.91e+11Hz -0.0133784 0.0029483
+ 2.911e+11Hz -0.0133371 0.00292965
+ 2.912e+11Hz -0.013296 0.00291067
+ 2.913e+11Hz -0.0132553 0.00289138
+ 2.914e+11Hz -0.0132149 0.00287178
+ 2.915e+11Hz -0.0131748 0.00285188
+ 2.916e+11Hz -0.013135 0.00283168
+ 2.917e+11Hz -0.0130955 0.0028112
+ 2.918e+11Hz -0.0130563 0.00279043
+ 2.919e+11Hz -0.0130175 0.00276938
+ 2.92e+11Hz -0.0129789 0.00274806
+ 2.921e+11Hz -0.0129407 0.00272648
+ 2.922e+11Hz -0.0129029 0.00270464
+ 2.923e+11Hz -0.0128653 0.00268255
+ 2.924e+11Hz -0.0128281 0.00266022
+ 2.925e+11Hz -0.0127913 0.00263765
+ 2.926e+11Hz -0.0127547 0.00261485
+ 2.927e+11Hz -0.0127186 0.00259183
+ 2.928e+11Hz -0.0126827 0.00256859
+ 2.929e+11Hz -0.0126472 0.00254514
+ 2.93e+11Hz -0.0126121 0.00252149
+ 2.931e+11Hz -0.0125773 0.00249764
+ 2.932e+11Hz -0.0125429 0.0024736
+ 2.933e+11Hz -0.0125088 0.00244938
+ 2.934e+11Hz -0.012475 0.00242498
+ 2.935e+11Hz -0.0124417 0.00240041
+ 2.936e+11Hz -0.0124087 0.00237569
+ 2.937e+11Hz -0.012376 0.0023508
+ 2.938e+11Hz -0.0123437 0.00232577
+ 2.939e+11Hz -0.0123117 0.00230059
+ 2.94e+11Hz -0.0122801 0.00227528
+ 2.941e+11Hz -0.0122489 0.00224984
+ 2.942e+11Hz -0.012218 0.00222428
+ 2.943e+11Hz -0.0121875 0.00219861
+ 2.944e+11Hz -0.0121574 0.00217282
+ 2.945e+11Hz -0.0121276 0.00214693
+ 2.946e+11Hz -0.0120981 0.00212095
+ 2.947e+11Hz -0.012069 0.00209488
+ 2.948e+11Hz -0.0120403 0.00206872
+ 2.949e+11Hz -0.0120119 0.00204249
+ 2.95e+11Hz -0.0119839 0.00201619
+ 2.951e+11Hz -0.0119562 0.00198983
+ 2.952e+11Hz -0.0119289 0.0019634
+ 2.953e+11Hz -0.0119019 0.00193693
+ 2.954e+11Hz -0.0118753 0.00191041
+ 2.955e+11Hz -0.011849 0.00188385
+ 2.956e+11Hz -0.0118231 0.00185725
+ 2.957e+11Hz -0.0117975 0.00183063
+ 2.958e+11Hz -0.0117722 0.00180398
+ 2.959e+11Hz -0.0117473 0.00177732
+ 2.96e+11Hz -0.0117228 0.00175065
+ 2.961e+11Hz -0.0116985 0.00172397
+ 2.962e+11Hz -0.0116746 0.0016973
+ 2.963e+11Hz -0.011651 0.00167063
+ 2.964e+11Hz -0.0116278 0.00164396
+ 2.965e+11Hz -0.0116048 0.00161732
+ 2.966e+11Hz -0.0115822 0.00159069
+ 2.967e+11Hz -0.0115599 0.00156409
+ 2.968e+11Hz -0.0115379 0.00153752
+ 2.969e+11Hz -0.0115163 0.00151099
+ 2.97e+11Hz -0.0114949 0.0014845
+ 2.971e+11Hz -0.0114738 0.00145805
+ 2.972e+11Hz -0.0114531 0.00143165
+ 2.973e+11Hz -0.0114326 0.0014053
+ 2.974e+11Hz -0.0114124 0.00137901
+ 2.975e+11Hz -0.0113926 0.00135278
+ 2.976e+11Hz -0.011373 0.00132662
+ 2.977e+11Hz -0.0113537 0.00130052
+ 2.978e+11Hz -0.0113347 0.0012745
+ 2.979e+11Hz -0.0113159 0.00124856
+ 2.98e+11Hz -0.0112974 0.00122269
+ 2.981e+11Hz -0.0112792 0.00119691
+ 2.982e+11Hz -0.0112613 0.00117122
+ 2.983e+11Hz -0.0112436 0.00114562
+ 2.984e+11Hz -0.0112262 0.00112011
+ 2.985e+11Hz -0.011209 0.0010947
+ 2.986e+11Hz -0.0111921 0.00106938
+ 2.987e+11Hz -0.0111754 0.00104417
+ 2.988e+11Hz -0.011159 0.00101906
+ 2.989e+11Hz -0.0111428 0.000994064
+ 2.99e+11Hz -0.0111268 0.000969174
+ 2.991e+11Hz -0.0111111 0.000944394
+ 2.992e+11Hz -0.0110956 0.000919729
+ 2.993e+11Hz -0.0110803 0.000895179
+ 2.994e+11Hz -0.0110652 0.000870747
+ 2.995e+11Hz -0.0110503 0.000846435
+ 2.996e+11Hz -0.0110357 0.000822244
+ 2.997e+11Hz -0.0110212 0.000798175
+ 2.998e+11Hz -0.0110069 0.000774231
+ 2.999e+11Hz -0.0109929 0.000750413
+ 3e+11Hz -0.010979 0.000726721
+ ]

.ENDS
.SUBCKT Sub_SPfile_X2 1 2 3
R1N 1 10 -50
R1P 10 11 100
R2N 2 20 -50
R2P 20 21 100

A11 %vd(10 3) %vd(11, 12) xfer1
.model xfer1 xfer R_I=true table=[
+ 0Hz 0.00482376 0
+ 1e+08Hz 0.00482395 1.93737e-06
+ 2e+08Hz 0.00482452 3.86743e-06
+ 3e+08Hz 0.00482548 5.78289e-06
+ 4e+08Hz 0.00482681 7.67645e-06
+ 5e+08Hz 0.00482853 9.54082e-06
+ 6e+08Hz 0.00483063 1.13687e-05
+ 7e+08Hz 0.0048331 1.3153e-05
+ 8e+08Hz 0.00483596 1.48863e-05
+ 9e+08Hz 0.00483919 1.65614e-05
+ 1e+09Hz 0.0048428 1.81712e-05
+ 1.1e+09Hz 0.00484679 1.97086e-05
+ 1.2e+09Hz 0.00485114 2.11664e-05
+ 1.3e+09Hz 0.00485587 2.25375e-05
+ 1.4e+09Hz 0.00486097 2.3815e-05
+ 1.5e+09Hz 0.00486643 2.49917e-05
+ 1.6e+09Hz 0.00487226 2.60609e-05
+ 1.7e+09Hz 0.00487846 2.70156e-05
+ 1.8e+09Hz 0.00488501 2.78489e-05
+ 1.9e+09Hz 0.00489192 2.85541e-05
+ 2e+09Hz 0.00489919 2.91245e-05
+ 2.1e+09Hz 0.00490681 2.95534e-05
+ 2.2e+09Hz 0.00491478 2.98342e-05
+ 2.3e+09Hz 0.00492309 2.99605e-05
+ 2.4e+09Hz 0.00493175 2.99257e-05
+ 2.5e+09Hz 0.00494075 2.97235e-05
+ 2.6e+09Hz 0.00495008 2.93477e-05
+ 2.7e+09Hz 0.00495975 2.87919e-05
+ 2.8e+09Hz 0.00496975 2.80502e-05
+ 2.9e+09Hz 0.00498007 2.71164e-05
+ 3e+09Hz 0.00499071 2.59846e-05
+ 3.1e+09Hz 0.00500167 2.4649e-05
+ 3.2e+09Hz 0.00501294 2.31038e-05
+ 3.3e+09Hz 0.00502452 2.13433e-05
+ 3.4e+09Hz 0.0050364 1.93619e-05
+ 3.5e+09Hz 0.00504859 1.71543e-05
+ 3.6e+09Hz 0.00506107 1.4715e-05
+ 3.7e+09Hz 0.00507383 1.20388e-05
+ 3.8e+09Hz 0.00508689 9.12049e-06
+ 3.9e+09Hz 0.00510022 5.9551e-06
+ 4e+09Hz 0.00511383 2.53768e-06
+ 4.1e+09Hz 0.00512771 -1.13658e-06
+ 4.2e+09Hz 0.00514185 -5.07238e-06
+ 4.3e+09Hz 0.00515626 -9.2743e-06
+ 4.4e+09Hz 0.00517091 -1.37468e-05
+ 4.5e+09Hz 0.00518582 -1.84942e-05
+ 4.6e+09Hz 0.00520097 -2.35208e-05
+ 4.7e+09Hz 0.00521636 -2.88306e-05
+ 4.8e+09Hz 0.00523198 -3.44276e-05
+ 4.9e+09Hz 0.00524782 -4.03157e-05
+ 5e+09Hz 0.00526389 -4.64986e-05
+ 5.1e+09Hz 0.00528017 -5.29798e-05
+ 5.2e+09Hz 0.00529666 -5.97629e-05
+ 5.3e+09Hz 0.00531335 -6.68512e-05
+ 5.4e+09Hz 0.00533024 -7.42479e-05
+ 5.5e+09Hz 0.00534732 -8.1956e-05
+ 5.6e+09Hz 0.00536459 -8.99785e-05
+ 5.7e+09Hz 0.00538203 -9.83183e-05
+ 5.8e+09Hz 0.00539964 -0.000106978
+ 5.9e+09Hz 0.00541742 -0.00011596
+ 6e+09Hz 0.00543536 -0.000125267
+ 6.1e+09Hz 0.00545346 -0.000134901
+ 6.2e+09Hz 0.0054717 -0.000144864
+ 6.3e+09Hz 0.00549008 -0.000155159
+ 6.4e+09Hz 0.00550859 -0.000165787
+ 6.5e+09Hz 0.00552723 -0.00017675
+ 6.6e+09Hz 0.005546 -0.000188049
+ 6.7e+09Hz 0.00556488 -0.000199686
+ 6.8e+09Hz 0.00558387 -0.000211663
+ 6.9e+09Hz 0.00560296 -0.00022398
+ 7e+09Hz 0.00562214 -0.000236638
+ 7.1e+09Hz 0.00564142 -0.000249639
+ 7.2e+09Hz 0.00566077 -0.000262984
+ 7.3e+09Hz 0.00568021 -0.000276673
+ 7.4e+09Hz 0.00569971 -0.000290706
+ 7.5e+09Hz 0.00571928 -0.000305084
+ 7.6e+09Hz 0.00573891 -0.000319807
+ 7.7e+09Hz 0.00575858 -0.000334876
+ 7.8e+09Hz 0.0057783 -0.00035029
+ 7.9e+09Hz 0.00579806 -0.00036605
+ 8e+09Hz 0.00581785 -0.000382155
+ 8.1e+09Hz 0.00583767 -0.000398604
+ 8.2e+09Hz 0.00585751 -0.000415398
+ 8.3e+09Hz 0.00587736 -0.000432536
+ 8.4e+09Hz 0.00589721 -0.000450016
+ 8.5e+09Hz 0.00591707 -0.000467839
+ 8.6e+09Hz 0.00593692 -0.000486003
+ 8.7e+09Hz 0.00595676 -0.000504507
+ 8.8e+09Hz 0.00597658 -0.00052335
+ 8.9e+09Hz 0.00599638 -0.000542531
+ 9e+09Hz 0.00601615 -0.000562048
+ 9.1e+09Hz 0.00603589 -0.0005819
+ 9.2e+09Hz 0.00605558 -0.000602085
+ 9.3e+09Hz 0.00607523 -0.000622601
+ 9.4e+09Hz 0.00609483 -0.000643447
+ 9.5e+09Hz 0.00611437 -0.00066462
+ 9.6e+09Hz 0.00613384 -0.000686119
+ 9.7e+09Hz 0.00615324 -0.000707941
+ 9.8e+09Hz 0.00617257 -0.000730084
+ 9.9e+09Hz 0.00619183 -0.000752546
+ 1e+10Hz 0.00621099 -0.000775324
+ 1.01e+10Hz 0.00623007 -0.000798416
+ 1.02e+10Hz 0.00624905 -0.000821819
+ 1.03e+10Hz 0.00626793 -0.000845531
+ 1.04e+10Hz 0.0062867 -0.000869548
+ 1.05e+10Hz 0.00630536 -0.000893868
+ 1.06e+10Hz 0.00632391 -0.000918487
+ 1.07e+10Hz 0.00634234 -0.000943403
+ 1.08e+10Hz 0.00636064 -0.000968612
+ 1.09e+10Hz 0.00637881 -0.000994112
+ 1.1e+10Hz 0.00639685 -0.0010199
+ 1.11e+10Hz 0.00641475 -0.00104597
+ 1.12e+10Hz 0.00643251 -0.00107232
+ 1.13e+10Hz 0.00645012 -0.00109895
+ 1.14e+10Hz 0.00646758 -0.00112585
+ 1.15e+10Hz 0.00648489 -0.00115302
+ 1.16e+10Hz 0.00650203 -0.00118045
+ 1.17e+10Hz 0.00651902 -0.00120815
+ 1.18e+10Hz 0.00653583 -0.00123611
+ 1.19e+10Hz 0.00655248 -0.00126432
+ 1.2e+10Hz 0.00656895 -0.00129278
+ 1.21e+10Hz 0.00658524 -0.00132148
+ 1.22e+10Hz 0.00660135 -0.00135043
+ 1.23e+10Hz 0.00661728 -0.00137962
+ 1.24e+10Hz 0.00663302 -0.00140904
+ 1.25e+10Hz 0.00664857 -0.00143869
+ 1.26e+10Hz 0.00666392 -0.00146857
+ 1.27e+10Hz 0.00667908 -0.00149867
+ 1.28e+10Hz 0.00669404 -0.00152899
+ 1.29e+10Hz 0.00670879 -0.00155951
+ 1.3e+10Hz 0.00672335 -0.00159025
+ 1.31e+10Hz 0.00673769 -0.00162119
+ 1.32e+10Hz 0.00675182 -0.00165234
+ 1.33e+10Hz 0.00676574 -0.00168367
+ 1.34e+10Hz 0.00677945 -0.0017152
+ 1.35e+10Hz 0.00679294 -0.00174692
+ 1.36e+10Hz 0.00680621 -0.00177882
+ 1.37e+10Hz 0.00681926 -0.00181089
+ 1.38e+10Hz 0.00683208 -0.00184314
+ 1.39e+10Hz 0.00684468 -0.00187555
+ 1.4e+10Hz 0.00685706 -0.00190813
+ 1.41e+10Hz 0.00686921 -0.00194087
+ 1.42e+10Hz 0.00688113 -0.00197377
+ 1.43e+10Hz 0.00689282 -0.00200681
+ 1.44e+10Hz 0.00690427 -0.00204001
+ 1.45e+10Hz 0.0069155 -0.00207334
+ 1.46e+10Hz 0.00692649 -0.00210681
+ 1.47e+10Hz 0.00693724 -0.00214041
+ 1.48e+10Hz 0.00694776 -0.00217414
+ 1.49e+10Hz 0.00695804 -0.00220799
+ 1.5e+10Hz 0.00696809 -0.00224196
+ 1.51e+10Hz 0.0069779 -0.00227604
+ 1.52e+10Hz 0.00698746 -0.00231024
+ 1.53e+10Hz 0.00699679 -0.00234454
+ 1.54e+10Hz 0.00700588 -0.00237894
+ 1.55e+10Hz 0.00701474 -0.00241344
+ 1.56e+10Hz 0.00702335 -0.00244802
+ 1.57e+10Hz 0.00703172 -0.0024827
+ 1.58e+10Hz 0.00703985 -0.00251746
+ 1.59e+10Hz 0.00704774 -0.0025523
+ 1.6e+10Hz 0.0070554 -0.00258721
+ 1.61e+10Hz 0.00706281 -0.00262219
+ 1.62e+10Hz 0.00706999 -0.00265724
+ 1.63e+10Hz 0.00707693 -0.00269235
+ 1.64e+10Hz 0.00708363 -0.00272752
+ 1.65e+10Hz 0.00709009 -0.00276274
+ 1.66e+10Hz 0.00709632 -0.00279801
+ 1.67e+10Hz 0.00710231 -0.00283332
+ 1.68e+10Hz 0.00710806 -0.00286868
+ 1.69e+10Hz 0.00711359 -0.00290407
+ 1.7e+10Hz 0.00711888 -0.0029395
+ 1.71e+10Hz 0.00712393 -0.00297496
+ 1.72e+10Hz 0.00712876 -0.00301044
+ 1.73e+10Hz 0.00713336 -0.00304594
+ 1.74e+10Hz 0.00713773 -0.00308147
+ 1.75e+10Hz 0.00714187 -0.003117
+ 1.76e+10Hz 0.00714579 -0.00315255
+ 1.77e+10Hz 0.00714948 -0.0031881
+ 1.78e+10Hz 0.00715295 -0.00322366
+ 1.79e+10Hz 0.00715621 -0.00325922
+ 1.8e+10Hz 0.00715924 -0.00329477
+ 1.81e+10Hz 0.00716205 -0.00333032
+ 1.82e+10Hz 0.00716465 -0.00336586
+ 1.83e+10Hz 0.00716703 -0.00340138
+ 1.84e+10Hz 0.00716921 -0.00343689
+ 1.85e+10Hz 0.00717117 -0.00347238
+ 1.86e+10Hz 0.00717293 -0.00350784
+ 1.87e+10Hz 0.00717447 -0.00354328
+ 1.88e+10Hz 0.00717582 -0.00357869
+ 1.89e+10Hz 0.00717696 -0.00361407
+ 1.9e+10Hz 0.00717791 -0.00364941
+ 1.91e+10Hz 0.00717866 -0.00368472
+ 1.92e+10Hz 0.00717921 -0.00371999
+ 1.93e+10Hz 0.00717957 -0.00375522
+ 1.94e+10Hz 0.00717974 -0.0037904
+ 1.95e+10Hz 0.00717972 -0.00382553
+ 1.96e+10Hz 0.00717951 -0.00386061
+ 1.97e+10Hz 0.00717912 -0.00389564
+ 1.98e+10Hz 0.00717856 -0.00393062
+ 1.99e+10Hz 0.00717781 -0.00396554
+ 2e+10Hz 0.00717689 -0.0040004
+ 2.01e+10Hz 0.00717579 -0.0040352
+ 2.02e+10Hz 0.00717453 -0.00406994
+ 2.03e+10Hz 0.00717309 -0.00410461
+ 2.04e+10Hz 0.00717149 -0.00413921
+ 2.05e+10Hz 0.00716973 -0.00417375
+ 2.06e+10Hz 0.00716781 -0.00420822
+ 2.07e+10Hz 0.00716573 -0.00424261
+ 2.08e+10Hz 0.0071635 -0.00427693
+ 2.09e+10Hz 0.00716111 -0.00431118
+ 2.1e+10Hz 0.00715858 -0.00434535
+ 2.11e+10Hz 0.0071559 -0.00437944
+ 2.12e+10Hz 0.00715308 -0.00441345
+ 2.13e+10Hz 0.00715011 -0.00444738
+ 2.14e+10Hz 0.00714701 -0.00448123
+ 2.15e+10Hz 0.00714377 -0.004515
+ 2.16e+10Hz 0.0071404 -0.00454868
+ 2.17e+10Hz 0.0071369 -0.00458228
+ 2.18e+10Hz 0.00713327 -0.0046158
+ 2.19e+10Hz 0.00712952 -0.00464922
+ 2.2e+10Hz 0.00712565 -0.00468256
+ 2.21e+10Hz 0.00712165 -0.00471582
+ 2.22e+10Hz 0.00711755 -0.00474898
+ 2.23e+10Hz 0.00711332 -0.00478206
+ 2.24e+10Hz 0.00710899 -0.00481504
+ 2.25e+10Hz 0.00710455 -0.00484794
+ 2.26e+10Hz 0.00710001 -0.00488074
+ 2.27e+10Hz 0.00709536 -0.00491346
+ 2.28e+10Hz 0.00709061 -0.00494608
+ 2.29e+10Hz 0.00708577 -0.00497862
+ 2.3e+10Hz 0.00708083 -0.00501106
+ 2.31e+10Hz 0.00707579 -0.00504341
+ 2.32e+10Hz 0.00707067 -0.00507567
+ 2.33e+10Hz 0.00706546 -0.00510784
+ 2.34e+10Hz 0.00706017 -0.00513992
+ 2.35e+10Hz 0.0070548 -0.00517191
+ 2.36e+10Hz 0.00704934 -0.00520381
+ 2.37e+10Hz 0.00704381 -0.00523561
+ 2.38e+10Hz 0.00703821 -0.00526733
+ 2.39e+10Hz 0.00703253 -0.00529896
+ 2.4e+10Hz 0.00702678 -0.0053305
+ 2.41e+10Hz 0.00702097 -0.00536195
+ 2.42e+10Hz 0.00701509 -0.00539332
+ 2.43e+10Hz 0.00700915 -0.00542459
+ 2.44e+10Hz 0.00700315 -0.00545578
+ 2.45e+10Hz 0.00699709 -0.00548688
+ 2.46e+10Hz 0.00699097 -0.0055179
+ 2.47e+10Hz 0.0069848 -0.00554884
+ 2.48e+10Hz 0.00697857 -0.00557969
+ 2.49e+10Hz 0.0069723 -0.00561046
+ 2.5e+10Hz 0.00696598 -0.00564114
+ 2.51e+10Hz 0.00695961 -0.00567175
+ 2.52e+10Hz 0.0069532 -0.00570228
+ 2.53e+10Hz 0.00694675 -0.00573272
+ 2.54e+10Hz 0.00694026 -0.00576309
+ 2.55e+10Hz 0.00693372 -0.00579339
+ 2.56e+10Hz 0.00692716 -0.00582361
+ 2.57e+10Hz 0.00692055 -0.00585375
+ 2.58e+10Hz 0.00691392 -0.00588382
+ 2.59e+10Hz 0.00690725 -0.00591382
+ 2.6e+10Hz 0.00690055 -0.00594375
+ 2.61e+10Hz 0.00689382 -0.00597361
+ 2.62e+10Hz 0.00688707 -0.0060034
+ 2.63e+10Hz 0.00688029 -0.00603313
+ 2.64e+10Hz 0.00687348 -0.00606279
+ 2.65e+10Hz 0.00686665 -0.00609239
+ 2.66e+10Hz 0.0068598 -0.00612192
+ 2.67e+10Hz 0.00685293 -0.00615139
+ 2.68e+10Hz 0.00684605 -0.00618081
+ 2.69e+10Hz 0.00683914 -0.00621016
+ 2.7e+10Hz 0.00683221 -0.00623947
+ 2.71e+10Hz 0.00682527 -0.00626871
+ 2.72e+10Hz 0.00681832 -0.0062979
+ 2.73e+10Hz 0.00681135 -0.00632704
+ 2.74e+10Hz 0.00680436 -0.00635613
+ 2.75e+10Hz 0.00679737 -0.00638517
+ 2.76e+10Hz 0.00679036 -0.00641417
+ 2.77e+10Hz 0.00678335 -0.00644311
+ 2.78e+10Hz 0.00677632 -0.00647202
+ 2.79e+10Hz 0.00676928 -0.00650088
+ 2.8e+10Hz 0.00676224 -0.0065297
+ 2.81e+10Hz 0.00675518 -0.00655848
+ 2.82e+10Hz 0.00674812 -0.00658722
+ 2.83e+10Hz 0.00674105 -0.00661593
+ 2.84e+10Hz 0.00673398 -0.0066446
+ 2.85e+10Hz 0.00672689 -0.00667324
+ 2.86e+10Hz 0.0067198 -0.00670184
+ 2.87e+10Hz 0.00671271 -0.00673042
+ 2.88e+10Hz 0.00670561 -0.00675897
+ 2.89e+10Hz 0.00669851 -0.00678749
+ 2.9e+10Hz 0.00669139 -0.00681599
+ 2.91e+10Hz 0.00668428 -0.00684446
+ 2.92e+10Hz 0.00667716 -0.00687291
+ 2.93e+10Hz 0.00667003 -0.00690134
+ 2.94e+10Hz 0.0066629 -0.00692975
+ 2.95e+10Hz 0.00665576 -0.00695814
+ 2.96e+10Hz 0.00664862 -0.00698652
+ 2.97e+10Hz 0.00664148 -0.00701488
+ 2.98e+10Hz 0.00663432 -0.00704322
+ 2.99e+10Hz 0.00662716 -0.00707156
+ 3e+10Hz 0.00662 -0.00709988
+ 3.01e+10Hz 0.00661283 -0.0071282
+ 3.02e+10Hz 0.00660565 -0.00715651
+ 3.03e+10Hz 0.00659846 -0.00718481
+ 3.04e+10Hz 0.00659127 -0.0072131
+ 3.05e+10Hz 0.00658407 -0.00724139
+ 3.06e+10Hz 0.00657686 -0.00726968
+ 3.07e+10Hz 0.00656964 -0.00729797
+ 3.08e+10Hz 0.00656241 -0.00732626
+ 3.09e+10Hz 0.00655517 -0.00735454
+ 3.1e+10Hz 0.00654792 -0.00738283
+ 3.11e+10Hz 0.00654066 -0.00741113
+ 3.12e+10Hz 0.00653339 -0.00743943
+ 3.13e+10Hz 0.0065261 -0.00746773
+ 3.14e+10Hz 0.0065188 -0.00749604
+ 3.15e+10Hz 0.00651149 -0.00752436
+ 3.16e+10Hz 0.00650416 -0.00755268
+ 3.17e+10Hz 0.00649682 -0.00758102
+ 3.18e+10Hz 0.00648946 -0.00760937
+ 3.19e+10Hz 0.00648208 -0.00763772
+ 3.2e+10Hz 0.00647468 -0.00766609
+ 3.21e+10Hz 0.00646726 -0.00769448
+ 3.22e+10Hz 0.00645983 -0.00772288
+ 3.23e+10Hz 0.00645237 -0.00775129
+ 3.24e+10Hz 0.00644489 -0.00777972
+ 3.25e+10Hz 0.00643738 -0.00780816
+ 3.26e+10Hz 0.00642986 -0.00783662
+ 3.27e+10Hz 0.0064223 -0.0078651
+ 3.28e+10Hz 0.00641473 -0.0078936
+ 3.29e+10Hz 0.00640712 -0.00792212
+ 3.3e+10Hz 0.00639949 -0.00795065
+ 3.31e+10Hz 0.00639182 -0.00797921
+ 3.32e+10Hz 0.00638413 -0.00800779
+ 3.33e+10Hz 0.00637641 -0.00803639
+ 3.34e+10Hz 0.00636865 -0.008065
+ 3.35e+10Hz 0.00636086 -0.00809365
+ 3.36e+10Hz 0.00635303 -0.00812231
+ 3.37e+10Hz 0.00634517 -0.008151
+ 3.38e+10Hz 0.00633728 -0.0081797
+ 3.39e+10Hz 0.00632934 -0.00820844
+ 3.4e+10Hz 0.00632137 -0.00823719
+ 3.41e+10Hz 0.00631335 -0.00826597
+ 3.42e+10Hz 0.0063053 -0.00829477
+ 3.43e+10Hz 0.0062972 -0.0083236
+ 3.44e+10Hz 0.00628906 -0.00835245
+ 3.45e+10Hz 0.00628087 -0.00838133
+ 3.46e+10Hz 0.00627264 -0.00841022
+ 3.47e+10Hz 0.00626436 -0.00843915
+ 3.48e+10Hz 0.00625603 -0.00846809
+ 3.49e+10Hz 0.00624766 -0.00849706
+ 3.5e+10Hz 0.00623923 -0.00852606
+ 3.51e+10Hz 0.00623075 -0.00855508
+ 3.52e+10Hz 0.00622222 -0.00858412
+ 3.53e+10Hz 0.00621364 -0.00861318
+ 3.54e+10Hz 0.006205 -0.00864227
+ 3.55e+10Hz 0.00619631 -0.00867138
+ 3.56e+10Hz 0.00618756 -0.00870052
+ 3.57e+10Hz 0.00617875 -0.00872968
+ 3.58e+10Hz 0.00616989 -0.00875885
+ 3.59e+10Hz 0.00616096 -0.00878805
+ 3.6e+10Hz 0.00615198 -0.00881728
+ 3.61e+10Hz 0.00614293 -0.00884652
+ 3.62e+10Hz 0.00613382 -0.00887578
+ 3.63e+10Hz 0.00612464 -0.00890507
+ 3.64e+10Hz 0.00611541 -0.00893437
+ 3.65e+10Hz 0.0061061 -0.00896369
+ 3.66e+10Hz 0.00609673 -0.00899303
+ 3.67e+10Hz 0.00608729 -0.00902239
+ 3.68e+10Hz 0.00607778 -0.00905177
+ 3.69e+10Hz 0.00606821 -0.00908116
+ 3.7e+10Hz 0.00605856 -0.00911057
+ 3.71e+10Hz 0.00604885 -0.00913999
+ 3.72e+10Hz 0.00603906 -0.00916943
+ 3.73e+10Hz 0.0060292 -0.00919888
+ 3.74e+10Hz 0.00601926 -0.00922835
+ 3.75e+10Hz 0.00600926 -0.00925783
+ 3.76e+10Hz 0.00599917 -0.00928732
+ 3.77e+10Hz 0.00598901 -0.00931682
+ 3.78e+10Hz 0.00597878 -0.00934633
+ 3.79e+10Hz 0.00596847 -0.00937585
+ 3.8e+10Hz 0.00595808 -0.00940538
+ 3.81e+10Hz 0.00594761 -0.00943492
+ 3.82e+10Hz 0.00593707 -0.00946447
+ 3.83e+10Hz 0.00592644 -0.00949402
+ 3.84e+10Hz 0.00591574 -0.00952358
+ 3.85e+10Hz 0.00590495 -0.00955314
+ 3.86e+10Hz 0.00589408 -0.0095827
+ 3.87e+10Hz 0.00588314 -0.00961227
+ 3.88e+10Hz 0.00587211 -0.00964184
+ 3.89e+10Hz 0.00586099 -0.00967141
+ 3.9e+10Hz 0.0058498 -0.00970098
+ 3.91e+10Hz 0.00583852 -0.00973055
+ 3.92e+10Hz 0.00582716 -0.00976011
+ 3.93e+10Hz 0.00581571 -0.00978968
+ 3.94e+10Hz 0.00580418 -0.00981924
+ 3.95e+10Hz 0.00579257 -0.00984879
+ 3.96e+10Hz 0.00578087 -0.00987834
+ 3.97e+10Hz 0.00576908 -0.00990788
+ 3.98e+10Hz 0.00575722 -0.00993741
+ 3.99e+10Hz 0.00574526 -0.00996694
+ 4e+10Hz 0.00573322 -0.00999645
+ 4.01e+10Hz 0.00572109 -0.010026
+ 4.02e+10Hz 0.00570888 -0.0100554
+ 4.03e+10Hz 0.00569658 -0.0100849
+ 4.04e+10Hz 0.00568419 -0.0101144
+ 4.05e+10Hz 0.00567172 -0.0101438
+ 4.06e+10Hz 0.00565916 -0.0101733
+ 4.07e+10Hz 0.00564652 -0.0102027
+ 4.08e+10Hz 0.00563379 -0.0102321
+ 4.09e+10Hz 0.00562097 -0.0102615
+ 4.1e+10Hz 0.00560807 -0.0102908
+ 4.11e+10Hz 0.00559508 -0.0103202
+ 4.12e+10Hz 0.00558201 -0.0103495
+ 4.13e+10Hz 0.00556884 -0.0103788
+ 4.14e+10Hz 0.0055556 -0.010408
+ 4.15e+10Hz 0.00554227 -0.0104373
+ 4.16e+10Hz 0.00552885 -0.0104665
+ 4.17e+10Hz 0.00551534 -0.0104957
+ 4.18e+10Hz 0.00550176 -0.0105248
+ 4.19e+10Hz 0.00548809 -0.010554
+ 4.2e+10Hz 0.00547433 -0.0105831
+ 4.21e+10Hz 0.00546049 -0.0106121
+ 4.22e+10Hz 0.00544656 -0.0106412
+ 4.23e+10Hz 0.00543256 -0.0106702
+ 4.24e+10Hz 0.00541846 -0.0106992
+ 4.25e+10Hz 0.00540429 -0.0107281
+ 4.26e+10Hz 0.00539004 -0.010757
+ 4.27e+10Hz 0.0053757 -0.0107859
+ 4.28e+10Hz 0.00536128 -0.0108147
+ 4.29e+10Hz 0.00534678 -0.0108435
+ 4.3e+10Hz 0.0053322 -0.0108723
+ 4.31e+10Hz 0.00531754 -0.010901
+ 4.32e+10Hz 0.0053028 -0.0109297
+ 4.33e+10Hz 0.00528798 -0.0109583
+ 4.34e+10Hz 0.00527308 -0.0109869
+ 4.35e+10Hz 0.00525811 -0.0110154
+ 4.36e+10Hz 0.00524306 -0.0110439
+ 4.37e+10Hz 0.00522793 -0.0110724
+ 4.38e+10Hz 0.00521272 -0.0111008
+ 4.39e+10Hz 0.00519744 -0.0111292
+ 4.4e+10Hz 0.00518209 -0.0111575
+ 4.41e+10Hz 0.00516666 -0.0111858
+ 4.42e+10Hz 0.00515116 -0.011214
+ 4.43e+10Hz 0.00513558 -0.0112422
+ 4.44e+10Hz 0.00511993 -0.0112703
+ 4.45e+10Hz 0.00510421 -0.0112984
+ 4.46e+10Hz 0.00508842 -0.0113265
+ 4.47e+10Hz 0.00507256 -0.0113545
+ 4.48e+10Hz 0.00505663 -0.0113824
+ 4.49e+10Hz 0.00504063 -0.0114103
+ 4.5e+10Hz 0.00502457 -0.0114381
+ 4.51e+10Hz 0.00500843 -0.0114659
+ 4.52e+10Hz 0.00499223 -0.0114936
+ 4.53e+10Hz 0.00497597 -0.0115213
+ 4.54e+10Hz 0.00495964 -0.0115489
+ 4.55e+10Hz 0.00494324 -0.0115765
+ 4.56e+10Hz 0.00492678 -0.011604
+ 4.57e+10Hz 0.00491026 -0.0116314
+ 4.58e+10Hz 0.00489368 -0.0116588
+ 4.59e+10Hz 0.00487703 -0.0116862
+ 4.6e+10Hz 0.00486033 -0.0117135
+ 4.61e+10Hz 0.00484356 -0.0117407
+ 4.62e+10Hz 0.00482674 -0.0117679
+ 4.63e+10Hz 0.00480986 -0.011795
+ 4.64e+10Hz 0.00479292 -0.011822
+ 4.65e+10Hz 0.00477592 -0.011849
+ 4.66e+10Hz 0.00475887 -0.011876
+ 4.67e+10Hz 0.00474177 -0.0119029
+ 4.68e+10Hz 0.00472461 -0.0119297
+ 4.69e+10Hz 0.0047074 -0.0119565
+ 4.7e+10Hz 0.00469013 -0.0119832
+ 4.71e+10Hz 0.00467281 -0.0120098
+ 4.72e+10Hz 0.00465544 -0.0120364
+ 4.73e+10Hz 0.00463803 -0.012063
+ 4.74e+10Hz 0.00462056 -0.0120895
+ 4.75e+10Hz 0.00460304 -0.0121159
+ 4.76e+10Hz 0.00458548 -0.0121422
+ 4.77e+10Hz 0.00456787 -0.0121685
+ 4.78e+10Hz 0.00455021 -0.0121948
+ 4.79e+10Hz 0.00453251 -0.012221
+ 4.8e+10Hz 0.00451476 -0.0122471
+ 4.81e+10Hz 0.00449697 -0.0122732
+ 4.82e+10Hz 0.00447914 -0.0122992
+ 4.83e+10Hz 0.00446126 -0.0123251
+ 4.84e+10Hz 0.00444334 -0.012351
+ 4.85e+10Hz 0.00442538 -0.0123769
+ 4.86e+10Hz 0.00440738 -0.0124027
+ 4.87e+10Hz 0.00438934 -0.0124284
+ 4.88e+10Hz 0.00437126 -0.0124541
+ 4.89e+10Hz 0.00435314 -0.0124797
+ 4.9e+10Hz 0.00433498 -0.0125052
+ 4.91e+10Hz 0.00431679 -0.0125307
+ 4.92e+10Hz 0.00429856 -0.0125561
+ 4.93e+10Hz 0.0042803 -0.0125815
+ 4.94e+10Hz 0.004262 -0.0126068
+ 4.95e+10Hz 0.00424366 -0.0126321
+ 4.96e+10Hz 0.00422529 -0.0126573
+ 4.97e+10Hz 0.00420689 -0.0126825
+ 4.98e+10Hz 0.00418846 -0.0127076
+ 4.99e+10Hz 0.00416999 -0.0127326
+ 5e+10Hz 0.00415149 -0.0127576
+ 5.01e+10Hz 0.00413296 -0.0127826
+ 5.02e+10Hz 0.0041144 -0.0128074
+ 5.03e+10Hz 0.00409581 -0.0128323
+ 5.04e+10Hz 0.00407719 -0.0128571
+ 5.05e+10Hz 0.00405854 -0.0128818
+ 5.06e+10Hz 0.00403987 -0.0129065
+ 5.07e+10Hz 0.00402116 -0.0129311
+ 5.08e+10Hz 0.00400243 -0.0129556
+ 5.09e+10Hz 0.00398367 -0.0129802
+ 5.1e+10Hz 0.00396488 -0.0130046
+ 5.11e+10Hz 0.00394607 -0.013029
+ 5.12e+10Hz 0.00392723 -0.0130534
+ 5.13e+10Hz 0.00390836 -0.0130777
+ 5.14e+10Hz 0.00388947 -0.013102
+ 5.15e+10Hz 0.00387056 -0.0131262
+ 5.16e+10Hz 0.00385162 -0.0131504
+ 5.17e+10Hz 0.00383265 -0.0131745
+ 5.18e+10Hz 0.00381367 -0.0131986
+ 5.19e+10Hz 0.00379466 -0.0132226
+ 5.2e+10Hz 0.00377562 -0.0132466
+ 5.21e+10Hz 0.00375656 -0.0132705
+ 5.22e+10Hz 0.00373748 -0.0132944
+ 5.23e+10Hz 0.00371838 -0.0133183
+ 5.24e+10Hz 0.00369925 -0.0133421
+ 5.25e+10Hz 0.00368011 -0.0133658
+ 5.26e+10Hz 0.00366094 -0.0133896
+ 5.27e+10Hz 0.00364175 -0.0134132
+ 5.28e+10Hz 0.00362253 -0.0134369
+ 5.29e+10Hz 0.0036033 -0.0134604
+ 5.3e+10Hz 0.00358404 -0.013484
+ 5.31e+10Hz 0.00356477 -0.0135075
+ 5.32e+10Hz 0.00354547 -0.013531
+ 5.33e+10Hz 0.00352615 -0.0135544
+ 5.34e+10Hz 0.00350681 -0.0135778
+ 5.35e+10Hz 0.00348745 -0.0136011
+ 5.36e+10Hz 0.00346807 -0.0136244
+ 5.37e+10Hz 0.00344867 -0.0136477
+ 5.38e+10Hz 0.00342925 -0.0136709
+ 5.39e+10Hz 0.0034098 -0.0136941
+ 5.4e+10Hz 0.00339034 -0.0137172
+ 5.41e+10Hz 0.00337085 -0.0137403
+ 5.42e+10Hz 0.00335135 -0.0137634
+ 5.43e+10Hz 0.00333182 -0.0137865
+ 5.44e+10Hz 0.00331228 -0.0138095
+ 5.45e+10Hz 0.00329271 -0.0138324
+ 5.46e+10Hz 0.00327312 -0.0138554
+ 5.47e+10Hz 0.00325351 -0.0138783
+ 5.48e+10Hz 0.00323388 -0.0139011
+ 5.49e+10Hz 0.00321423 -0.013924
+ 5.5e+10Hz 0.00319455 -0.0139468
+ 5.51e+10Hz 0.00317486 -0.0139695
+ 5.52e+10Hz 0.00315514 -0.0139923
+ 5.53e+10Hz 0.0031354 -0.014015
+ 5.54e+10Hz 0.00311564 -0.0140376
+ 5.55e+10Hz 0.00309586 -0.0140603
+ 5.56e+10Hz 0.00307606 -0.0140829
+ 5.57e+10Hz 0.00305623 -0.0141055
+ 5.58e+10Hz 0.00303638 -0.014128
+ 5.59e+10Hz 0.00301651 -0.0141505
+ 5.6e+10Hz 0.00299662 -0.014173
+ 5.61e+10Hz 0.0029767 -0.0141955
+ 5.62e+10Hz 0.00295676 -0.0142179
+ 5.63e+10Hz 0.00293679 -0.0142403
+ 5.64e+10Hz 0.0029168 -0.0142626
+ 5.65e+10Hz 0.00289679 -0.014285
+ 5.66e+10Hz 0.00287675 -0.0143073
+ 5.67e+10Hz 0.00285669 -0.0143296
+ 5.68e+10Hz 0.0028366 -0.0143518
+ 5.69e+10Hz 0.00281649 -0.014374
+ 5.7e+10Hz 0.00279635 -0.0143962
+ 5.71e+10Hz 0.00277619 -0.0144184
+ 5.72e+10Hz 0.002756 -0.0144406
+ 5.73e+10Hz 0.00273579 -0.0144627
+ 5.74e+10Hz 0.00271554 -0.0144848
+ 5.75e+10Hz 0.00269527 -0.0145068
+ 5.76e+10Hz 0.00267498 -0.0145288
+ 5.77e+10Hz 0.00265465 -0.0145509
+ 5.78e+10Hz 0.0026343 -0.0145728
+ 5.79e+10Hz 0.00261392 -0.0145948
+ 5.8e+10Hz 0.00259351 -0.0146167
+ 5.81e+10Hz 0.00257308 -0.0146386
+ 5.82e+10Hz 0.00255261 -0.0146605
+ 5.83e+10Hz 0.00253212 -0.0146823
+ 5.84e+10Hz 0.00251159 -0.0147042
+ 5.85e+10Hz 0.00249104 -0.014726
+ 5.86e+10Hz 0.00247045 -0.0147477
+ 5.87e+10Hz 0.00244984 -0.0147695
+ 5.88e+10Hz 0.00242919 -0.0147912
+ 5.89e+10Hz 0.00240851 -0.0148129
+ 5.9e+10Hz 0.00238781 -0.0148345
+ 5.91e+10Hz 0.00236707 -0.0148562
+ 5.92e+10Hz 0.00234629 -0.0148778
+ 5.93e+10Hz 0.00232549 -0.0148994
+ 5.94e+10Hz 0.00230465 -0.0149209
+ 5.95e+10Hz 0.00228378 -0.0149425
+ 5.96e+10Hz 0.00226287 -0.014964
+ 5.97e+10Hz 0.00224194 -0.0149854
+ 5.98e+10Hz 0.00222096 -0.0150069
+ 5.99e+10Hz 0.00219996 -0.0150283
+ 6e+10Hz 0.00217892 -0.0150497
+ 6.01e+10Hz 0.00215784 -0.0150711
+ 6.02e+10Hz 0.00213673 -0.0150924
+ 6.03e+10Hz 0.00211559 -0.0151137
+ 6.04e+10Hz 0.00209441 -0.015135
+ 6.05e+10Hz 0.00207319 -0.0151563
+ 6.06e+10Hz 0.00205194 -0.0151775
+ 6.07e+10Hz 0.00203065 -0.0151987
+ 6.08e+10Hz 0.00200932 -0.0152199
+ 6.09e+10Hz 0.00198796 -0.015241
+ 6.1e+10Hz 0.00196656 -0.0152621
+ 6.11e+10Hz 0.00194512 -0.0152832
+ 6.12e+10Hz 0.00192364 -0.0153043
+ 6.13e+10Hz 0.00190213 -0.0153253
+ 6.14e+10Hz 0.00188058 -0.0153463
+ 6.15e+10Hz 0.00185899 -0.0153672
+ 6.16e+10Hz 0.00183736 -0.0153882
+ 6.17e+10Hz 0.0018157 -0.0154091
+ 6.18e+10Hz 0.00179399 -0.0154299
+ 6.19e+10Hz 0.00177225 -0.0154508
+ 6.2e+10Hz 0.00175047 -0.0154716
+ 6.21e+10Hz 0.00172865 -0.0154924
+ 6.22e+10Hz 0.00170678 -0.0155131
+ 6.23e+10Hz 0.00168488 -0.0155338
+ 6.24e+10Hz 0.00166294 -0.0155545
+ 6.25e+10Hz 0.00164096 -0.0155751
+ 6.26e+10Hz 0.00161894 -0.0155957
+ 6.27e+10Hz 0.00159688 -0.0156163
+ 6.28e+10Hz 0.00157478 -0.0156368
+ 6.29e+10Hz 0.00155264 -0.0156574
+ 6.3e+10Hz 0.00153046 -0.0156778
+ 6.31e+10Hz 0.00150824 -0.0156983
+ 6.32e+10Hz 0.00148597 -0.0157187
+ 6.33e+10Hz 0.00146367 -0.015739
+ 6.34e+10Hz 0.00144133 -0.0157593
+ 6.35e+10Hz 0.00141894 -0.0157796
+ 6.36e+10Hz 0.00139652 -0.0157999
+ 6.37e+10Hz 0.00137405 -0.0158201
+ 6.38e+10Hz 0.00135155 -0.0158403
+ 6.39e+10Hz 0.001329 -0.0158604
+ 6.4e+10Hz 0.00130641 -0.0158805
+ 6.41e+10Hz 0.00128378 -0.0159006
+ 6.42e+10Hz 0.00126111 -0.0159206
+ 6.43e+10Hz 0.00123841 -0.0159406
+ 6.44e+10Hz 0.00121566 -0.0159605
+ 6.45e+10Hz 0.00119286 -0.0159804
+ 6.46e+10Hz 0.00117003 -0.0160003
+ 6.47e+10Hz 0.00114716 -0.0160201
+ 6.48e+10Hz 0.00112425 -0.0160399
+ 6.49e+10Hz 0.0011013 -0.0160596
+ 6.5e+10Hz 0.0010783 -0.0160793
+ 6.51e+10Hz 0.00105527 -0.0160989
+ 6.52e+10Hz 0.0010322 -0.0161185
+ 6.53e+10Hz 0.00100909 -0.0161381
+ 6.54e+10Hz 0.000985935 -0.0161576
+ 6.55e+10Hz 0.000962743 -0.0161771
+ 6.56e+10Hz 0.000939512 -0.0161965
+ 6.57e+10Hz 0.000916242 -0.0162159
+ 6.58e+10Hz 0.000892933 -0.0162352
+ 6.59e+10Hz 0.000869584 -0.0162545
+ 6.6e+10Hz 0.000846197 -0.0162737
+ 6.61e+10Hz 0.000822772 -0.0162929
+ 6.62e+10Hz 0.000799308 -0.0163121
+ 6.63e+10Hz 0.000775805 -0.0163312
+ 6.64e+10Hz 0.000752265 -0.0163502
+ 6.65e+10Hz 0.000728688 -0.0163693
+ 6.66e+10Hz 0.000705072 -0.0163882
+ 6.67e+10Hz 0.00068142 -0.0164071
+ 6.68e+10Hz 0.00065773 -0.016426
+ 6.69e+10Hz 0.000634004 -0.0164448
+ 6.7e+10Hz 0.000610241 -0.0164636
+ 6.71e+10Hz 0.000586442 -0.0164823
+ 6.72e+10Hz 0.000562607 -0.0165009
+ 6.73e+10Hz 0.000538736 -0.0165195
+ 6.74e+10Hz 0.00051483 -0.0165381
+ 6.75e+10Hz 0.000490889 -0.0165566
+ 6.76e+10Hz 0.000466913 -0.0165751
+ 6.77e+10Hz 0.000442902 -0.0165935
+ 6.78e+10Hz 0.000418857 -0.0166118
+ 6.79e+10Hz 0.000394778 -0.0166301
+ 6.8e+10Hz 0.000370666 -0.0166484
+ 6.81e+10Hz 0.00034652 -0.0166666
+ 6.82e+10Hz 0.000322341 -0.0166847
+ 6.83e+10Hz 0.00029813 -0.0167028
+ 6.84e+10Hz 0.000273886 -0.0167209
+ 6.85e+10Hz 0.000249611 -0.0167388
+ 6.86e+10Hz 0.000225304 -0.0167568
+ 6.87e+10Hz 0.000200965 -0.0167747
+ 6.88e+10Hz 0.000176596 -0.0167925
+ 6.89e+10Hz 0.000152196 -0.0168102
+ 6.9e+10Hz 0.000127766 -0.016828
+ 6.91e+10Hz 0.000103306 -0.0168456
+ 6.92e+10Hz 7.88161e-05 -0.0168632
+ 6.93e+10Hz 5.42975e-05 -0.0168808
+ 6.94e+10Hz 2.97502e-05 -0.0168983
+ 6.95e+10Hz 5.17445e-06 -0.0169157
+ 6.96e+10Hz -1.94293e-05 -0.0169331
+ 6.97e+10Hz -4.40606e-05 -0.0169504
+ 6.98e+10Hz -6.87192e-05 -0.0169677
+ 6.99e+10Hz -9.34047e-05 -0.0169849
+ 7e+10Hz -0.000118117 -0.0170021
+ 7.01e+10Hz -0.000142855 -0.0170192
+ 7.02e+10Hz -0.000167619 -0.0170362
+ 7.03e+10Hz -0.000192408 -0.0170532
+ 7.04e+10Hz -0.000217222 -0.0170701
+ 7.05e+10Hz -0.00024206 -0.017087
+ 7.06e+10Hz -0.000266923 -0.0171039
+ 7.07e+10Hz -0.00029181 -0.0171206
+ 7.08e+10Hz -0.00031672 -0.0171373
+ 7.09e+10Hz -0.000341654 -0.017154
+ 7.1e+10Hz -0.000366609 -0.0171706
+ 7.11e+10Hz -0.000391588 -0.0171871
+ 7.12e+10Hz -0.000416588 -0.0172036
+ 7.13e+10Hz -0.000441609 -0.01722
+ 7.14e+10Hz -0.000466652 -0.0172364
+ 7.15e+10Hz -0.000491716 -0.0172527
+ 7.16e+10Hz -0.0005168 -0.017269
+ 7.17e+10Hz -0.000541904 -0.0172852
+ 7.18e+10Hz -0.000567028 -0.0173013
+ 7.19e+10Hz -0.000592171 -0.0173174
+ 7.2e+10Hz -0.000617333 -0.0173335
+ 7.21e+10Hz -0.000642514 -0.0173494
+ 7.22e+10Hz -0.000667713 -0.0173654
+ 7.23e+10Hz -0.000692929 -0.0173812
+ 7.24e+10Hz -0.000718164 -0.017397
+ 7.25e+10Hz -0.000743415 -0.0174128
+ 7.26e+10Hz -0.000768684 -0.0174285
+ 7.27e+10Hz -0.000793969 -0.0174441
+ 7.28e+10Hz -0.00081927 -0.0174597
+ 7.29e+10Hz -0.000844587 -0.0174752
+ 7.3e+10Hz -0.000869919 -0.0174907
+ 7.31e+10Hz -0.000895267 -0.0175061
+ 7.32e+10Hz -0.000920629 -0.0175215
+ 7.33e+10Hz -0.000946006 -0.0175368
+ 7.34e+10Hz -0.000971398 -0.017552
+ 7.35e+10Hz -0.000996803 -0.0175672
+ 7.36e+10Hz -0.00102222 -0.0175824
+ 7.37e+10Hz -0.00104765 -0.0175975
+ 7.38e+10Hz -0.0010731 -0.0176125
+ 7.39e+10Hz -0.00109856 -0.0176275
+ 7.4e+10Hz -0.00112403 -0.0176424
+ 7.41e+10Hz -0.00114951 -0.0176573
+ 7.42e+10Hz -0.00117501 -0.0176721
+ 7.43e+10Hz -0.00120051 -0.0176869
+ 7.44e+10Hz -0.00122603 -0.0177016
+ 7.45e+10Hz -0.00125156 -0.0177162
+ 7.46e+10Hz -0.0012771 -0.0177308
+ 7.47e+10Hz -0.00130265 -0.0177454
+ 7.48e+10Hz -0.00132821 -0.0177599
+ 7.49e+10Hz -0.00135379 -0.0177743
+ 7.5e+10Hz -0.00137937 -0.0177887
+ 7.51e+10Hz -0.00140496 -0.0178031
+ 7.52e+10Hz -0.00143056 -0.0178174
+ 7.53e+10Hz -0.00145617 -0.0178316
+ 7.54e+10Hz -0.00148179 -0.0178458
+ 7.55e+10Hz -0.00150742 -0.0178599
+ 7.56e+10Hz -0.00153306 -0.017874
+ 7.57e+10Hz -0.00155871 -0.0178881
+ 7.58e+10Hz -0.00158436 -0.0179021
+ 7.59e+10Hz -0.00161003 -0.017916
+ 7.6e+10Hz -0.0016357 -0.0179299
+ 7.61e+10Hz -0.00166138 -0.0179437
+ 7.62e+10Hz -0.00168707 -0.0179575
+ 7.63e+10Hz -0.00171277 -0.0179712
+ 7.64e+10Hz -0.00173847 -0.0179849
+ 7.65e+10Hz -0.00176418 -0.0179986
+ 7.66e+10Hz -0.0017899 -0.0180121
+ 7.67e+10Hz -0.00181563 -0.0180257
+ 7.68e+10Hz -0.00184136 -0.0180392
+ 7.69e+10Hz -0.0018671 -0.0180526
+ 7.7e+10Hz -0.00189285 -0.018066
+ 7.71e+10Hz -0.00191861 -0.0180794
+ 7.72e+10Hz -0.00194437 -0.0180927
+ 7.73e+10Hz -0.00197014 -0.0181059
+ 7.74e+10Hz -0.00199592 -0.0181191
+ 7.75e+10Hz -0.0020217 -0.0181323
+ 7.76e+10Hz -0.00204749 -0.0181454
+ 7.77e+10Hz -0.00207328 -0.0181585
+ 7.78e+10Hz -0.00209909 -0.0181715
+ 7.79e+10Hz -0.0021249 -0.0181845
+ 7.8e+10Hz -0.00215071 -0.0181974
+ 7.81e+10Hz -0.00217654 -0.0182103
+ 7.82e+10Hz -0.00220237 -0.0182231
+ 7.83e+10Hz -0.0022282 -0.0182359
+ 7.84e+10Hz -0.00225405 -0.0182487
+ 7.85e+10Hz -0.0022799 -0.0182614
+ 7.86e+10Hz -0.00230575 -0.018274
+ 7.87e+10Hz -0.00233162 -0.0182867
+ 7.88e+10Hz -0.00235749 -0.0182992
+ 7.89e+10Hz -0.00238336 -0.0183118
+ 7.9e+10Hz -0.00240925 -0.0183242
+ 7.91e+10Hz -0.00243514 -0.0183367
+ 7.92e+10Hz -0.00246103 -0.0183491
+ 7.93e+10Hz -0.00248694 -0.0183614
+ 7.94e+10Hz -0.00251285 -0.0183737
+ 7.95e+10Hz -0.00253876 -0.018386
+ 7.96e+10Hz -0.00256469 -0.0183982
+ 7.97e+10Hz -0.00259062 -0.0184104
+ 7.98e+10Hz -0.00261656 -0.0184226
+ 7.99e+10Hz -0.00264251 -0.0184347
+ 8e+10Hz -0.00266846 -0.0184467
+ 8.01e+10Hz -0.00269442 -0.0184587
+ 8.02e+10Hz -0.00272039 -0.0184707
+ 8.03e+10Hz -0.00274637 -0.0184826
+ 8.04e+10Hz -0.00277235 -0.0184945
+ 8.05e+10Hz -0.00279834 -0.0185064
+ 8.06e+10Hz -0.00282434 -0.0185182
+ 8.07e+10Hz -0.00285035 -0.0185299
+ 8.08e+10Hz -0.00287637 -0.0185417
+ 8.09e+10Hz -0.00290239 -0.0185534
+ 8.1e+10Hz -0.00292842 -0.018565
+ 8.11e+10Hz -0.00295446 -0.0185766
+ 8.12e+10Hz -0.00298051 -0.0185882
+ 8.13e+10Hz -0.00300657 -0.0185997
+ 8.14e+10Hz -0.00303264 -0.0186111
+ 8.15e+10Hz -0.00305872 -0.0186226
+ 8.16e+10Hz -0.0030848 -0.018634
+ 8.17e+10Hz -0.00311089 -0.0186453
+ 8.18e+10Hz -0.003137 -0.0186567
+ 8.19e+10Hz -0.00316311 -0.0186679
+ 8.2e+10Hz -0.00318923 -0.0186792
+ 8.21e+10Hz -0.00321537 -0.0186904
+ 8.22e+10Hz -0.00324151 -0.0187015
+ 8.23e+10Hz -0.00326766 -0.0187126
+ 8.24e+10Hz -0.00329382 -0.0187237
+ 8.25e+10Hz -0.00332 -0.0187347
+ 8.26e+10Hz -0.00334618 -0.0187457
+ 8.27e+10Hz -0.00337237 -0.0187567
+ 8.28e+10Hz -0.00339858 -0.0187676
+ 8.29e+10Hz -0.00342479 -0.0187784
+ 8.3e+10Hz -0.00345102 -0.0187893
+ 8.31e+10Hz -0.00347725 -0.0188001
+ 8.32e+10Hz -0.0035035 -0.0188108
+ 8.33e+10Hz -0.00352976 -0.0188215
+ 8.34e+10Hz -0.00355603 -0.0188322
+ 8.35e+10Hz -0.00358231 -0.0188428
+ 8.36e+10Hz -0.00360861 -0.0188534
+ 8.37e+10Hz -0.00363491 -0.0188639
+ 8.38e+10Hz -0.00366123 -0.0188744
+ 8.39e+10Hz -0.00368756 -0.0188849
+ 8.4e+10Hz -0.0037139 -0.0188953
+ 8.41e+10Hz -0.00374026 -0.0189057
+ 8.42e+10Hz -0.00376662 -0.018916
+ 8.43e+10Hz -0.003793 -0.0189263
+ 8.44e+10Hz -0.00381939 -0.0189366
+ 8.45e+10Hz -0.0038458 -0.0189468
+ 8.46e+10Hz -0.00387221 -0.018957
+ 8.47e+10Hz -0.00389864 -0.0189671
+ 8.48e+10Hz -0.00392508 -0.0189772
+ 8.49e+10Hz -0.00395154 -0.0189872
+ 8.5e+10Hz -0.00397801 -0.0189972
+ 8.51e+10Hz -0.00400449 -0.0190072
+ 8.52e+10Hz -0.00403099 -0.0190171
+ 8.53e+10Hz -0.00405749 -0.019027
+ 8.54e+10Hz -0.00408402 -0.0190368
+ 8.55e+10Hz -0.00411055 -0.0190466
+ 8.56e+10Hz -0.0041371 -0.0190563
+ 8.57e+10Hz -0.00416367 -0.019066
+ 8.58e+10Hz -0.00419024 -0.0190757
+ 8.59e+10Hz -0.00421683 -0.0190853
+ 8.6e+10Hz -0.00424344 -0.0190948
+ 8.61e+10Hz -0.00427006 -0.0191044
+ 8.62e+10Hz -0.00429669 -0.0191138
+ 8.63e+10Hz -0.00432333 -0.0191233
+ 8.64e+10Hz -0.00435 -0.0191327
+ 8.65e+10Hz -0.00437667 -0.019142
+ 8.66e+10Hz -0.00440336 -0.0191513
+ 8.67e+10Hz -0.00443006 -0.0191606
+ 8.68e+10Hz -0.00445678 -0.0191698
+ 8.69e+10Hz -0.00448351 -0.0191789
+ 8.7e+10Hz -0.00451025 -0.0191881
+ 8.71e+10Hz -0.00453701 -0.0191971
+ 8.72e+10Hz -0.00456379 -0.0192062
+ 8.73e+10Hz -0.00459057 -0.0192151
+ 8.74e+10Hz -0.00461738 -0.0192241
+ 8.75e+10Hz -0.00464419 -0.0192329
+ 8.76e+10Hz -0.00467102 -0.0192418
+ 8.77e+10Hz -0.00469786 -0.0192506
+ 8.78e+10Hz -0.00472472 -0.0192593
+ 8.79e+10Hz -0.00475159 -0.019268
+ 8.8e+10Hz -0.00477848 -0.0192766
+ 8.81e+10Hz -0.00480538 -0.0192852
+ 8.82e+10Hz -0.00483229 -0.0192938
+ 8.83e+10Hz -0.00485922 -0.0193023
+ 8.84e+10Hz -0.00488616 -0.0193107
+ 8.85e+10Hz -0.00491311 -0.0193191
+ 8.86e+10Hz -0.00494008 -0.0193275
+ 8.87e+10Hz -0.00496706 -0.0193358
+ 8.88e+10Hz -0.00499405 -0.019344
+ 8.89e+10Hz -0.00502106 -0.0193522
+ 8.9e+10Hz -0.00504808 -0.0193604
+ 8.91e+10Hz -0.00507512 -0.0193685
+ 8.92e+10Hz -0.00510216 -0.0193765
+ 8.93e+10Hz -0.00512922 -0.0193845
+ 8.94e+10Hz -0.00515629 -0.0193925
+ 8.95e+10Hz -0.00518338 -0.0194004
+ 8.96e+10Hz -0.00521047 -0.0194082
+ 8.97e+10Hz -0.00523758 -0.019416
+ 8.98e+10Hz -0.0052647 -0.0194237
+ 8.99e+10Hz -0.00529184 -0.0194314
+ 9e+10Hz -0.00531898 -0.019439
+ 9.01e+10Hz -0.00534614 -0.0194466
+ 9.02e+10Hz -0.0053733 -0.0194541
+ 9.03e+10Hz -0.00540048 -0.0194616
+ 9.04e+10Hz -0.00542767 -0.019469
+ 9.05e+10Hz -0.00545487 -0.0194764
+ 9.06e+10Hz -0.00548208 -0.0194837
+ 9.07e+10Hz -0.00550931 -0.0194909
+ 9.08e+10Hz -0.00553654 -0.0194981
+ 9.09e+10Hz -0.00556378 -0.0195053
+ 9.1e+10Hz -0.00559103 -0.0195124
+ 9.11e+10Hz -0.00561829 -0.0195194
+ 9.12e+10Hz -0.00564557 -0.0195264
+ 9.13e+10Hz -0.00567285 -0.0195333
+ 9.14e+10Hz -0.00570014 -0.0195402
+ 9.15e+10Hz -0.00572743 -0.019547
+ 9.16e+10Hz -0.00575474 -0.0195537
+ 9.17e+10Hz -0.00578206 -0.0195604
+ 9.18e+10Hz -0.00580938 -0.0195671
+ 9.19e+10Hz -0.00583671 -0.0195737
+ 9.2e+10Hz -0.00586405 -0.0195802
+ 9.21e+10Hz -0.0058914 -0.0195867
+ 9.22e+10Hz -0.00591875 -0.0195931
+ 9.23e+10Hz -0.00594611 -0.0195994
+ 9.24e+10Hz -0.00597347 -0.0196057
+ 9.25e+10Hz -0.00600085 -0.019612
+ 9.26e+10Hz -0.00602823 -0.0196182
+ 9.27e+10Hz -0.00605561 -0.0196243
+ 9.28e+10Hz -0.006083 -0.0196304
+ 9.29e+10Hz -0.00611039 -0.0196364
+ 9.3e+10Hz -0.00613779 -0.0196423
+ 9.31e+10Hz -0.0061652 -0.0196482
+ 9.32e+10Hz -0.00619261 -0.019654
+ 9.33e+10Hz -0.00622002 -0.0196598
+ 9.34e+10Hz -0.00624744 -0.0196655
+ 9.35e+10Hz -0.00627485 -0.0196712
+ 9.36e+10Hz -0.00630228 -0.0196768
+ 9.37e+10Hz -0.0063297 -0.0196823
+ 9.38e+10Hz -0.00635713 -0.0196878
+ 9.39e+10Hz -0.00638456 -0.0196932
+ 9.4e+10Hz -0.00641199 -0.0196986
+ 9.41e+10Hz -0.00643943 -0.0197039
+ 9.42e+10Hz -0.00646686 -0.0197091
+ 9.43e+10Hz -0.0064943 -0.0197143
+ 9.44e+10Hz -0.00652173 -0.0197194
+ 9.45e+10Hz -0.00654917 -0.0197245
+ 9.46e+10Hz -0.0065766 -0.0197295
+ 9.47e+10Hz -0.00660404 -0.0197344
+ 9.48e+10Hz -0.00663148 -0.0197393
+ 9.49e+10Hz -0.00665891 -0.0197441
+ 9.5e+10Hz -0.00668634 -0.0197489
+ 9.51e+10Hz -0.00671377 -0.0197536
+ 9.52e+10Hz -0.0067412 -0.0197582
+ 9.53e+10Hz -0.00676863 -0.0197628
+ 9.54e+10Hz -0.00679605 -0.0197673
+ 9.55e+10Hz -0.00682347 -0.0197718
+ 9.56e+10Hz -0.00685089 -0.0197762
+ 9.57e+10Hz -0.00687831 -0.0197805
+ 9.58e+10Hz -0.00690572 -0.0197848
+ 9.59e+10Hz -0.00693312 -0.019789
+ 9.6e+10Hz -0.00696052 -0.0197932
+ 9.61e+10Hz -0.00698792 -0.0197973
+ 9.62e+10Hz -0.00701531 -0.0198014
+ 9.63e+10Hz -0.0070427 -0.0198053
+ 9.64e+10Hz -0.00707008 -0.0198093
+ 9.65e+10Hz -0.00709745 -0.0198131
+ 9.66e+10Hz -0.00712482 -0.0198169
+ 9.67e+10Hz -0.00715218 -0.0198207
+ 9.68e+10Hz -0.00717953 -0.0198243
+ 9.69e+10Hz -0.00720688 -0.019828
+ 9.7e+10Hz -0.00723421 -0.0198315
+ 9.71e+10Hz -0.00726154 -0.019835
+ 9.72e+10Hz -0.00728887 -0.0198385
+ 9.73e+10Hz -0.00731618 -0.0198418
+ 9.74e+10Hz -0.00734348 -0.0198452
+ 9.75e+10Hz -0.00737078 -0.0198484
+ 9.76e+10Hz -0.00739806 -0.0198516
+ 9.77e+10Hz -0.00742533 -0.0198548
+ 9.78e+10Hz -0.0074526 -0.0198579
+ 9.79e+10Hz -0.00747985 -0.0198609
+ 9.8e+10Hz -0.0075071 -0.0198639
+ 9.81e+10Hz -0.00753433 -0.0198668
+ 9.82e+10Hz -0.00756155 -0.0198696
+ 9.83e+10Hz -0.00758876 -0.0198724
+ 9.84e+10Hz -0.00761595 -0.0198752
+ 9.85e+10Hz -0.00764314 -0.0198778
+ 9.86e+10Hz -0.00767031 -0.0198805
+ 9.87e+10Hz -0.00769747 -0.019883
+ 9.88e+10Hz -0.00772461 -0.0198855
+ 9.89e+10Hz -0.00775175 -0.019888
+ 9.9e+10Hz -0.00777887 -0.0198904
+ 9.91e+10Hz -0.00780597 -0.0198927
+ 9.92e+10Hz -0.00783306 -0.019895
+ 9.93e+10Hz -0.00786014 -0.0198972
+ 9.94e+10Hz -0.0078872 -0.0198993
+ 9.95e+10Hz -0.00791425 -0.0199014
+ 9.96e+10Hz -0.00794128 -0.0199035
+ 9.97e+10Hz -0.00796829 -0.0199055
+ 9.98e+10Hz -0.0079953 -0.0199074
+ 9.99e+10Hz -0.00802228 -0.0199093
+ 1e+11Hz -0.00804925 -0.0199111
+ 1.001e+11Hz -0.0080762 -0.0199129
+ 1.002e+11Hz -0.00810314 -0.0199146
+ 1.003e+11Hz -0.00813006 -0.0199162
+ 1.004e+11Hz -0.00815696 -0.0199178
+ 1.005e+11Hz -0.00818384 -0.0199194
+ 1.006e+11Hz -0.00821071 -0.0199209
+ 1.007e+11Hz -0.00823756 -0.0199223
+ 1.008e+11Hz -0.00826439 -0.0199237
+ 1.009e+11Hz -0.00829121 -0.019925
+ 1.01e+11Hz -0.008318 -0.0199263
+ 1.011e+11Hz -0.00834478 -0.0199275
+ 1.012e+11Hz -0.00837154 -0.0199287
+ 1.013e+11Hz -0.00839828 -0.0199298
+ 1.014e+11Hz -0.008425 -0.0199309
+ 1.015e+11Hz -0.0084517 -0.0199319
+ 1.016e+11Hz -0.00847838 -0.0199328
+ 1.017e+11Hz -0.00850504 -0.0199337
+ 1.018e+11Hz -0.00853169 -0.0199346
+ 1.019e+11Hz -0.00855831 -0.0199354
+ 1.02e+11Hz -0.00858491 -0.0199361
+ 1.021e+11Hz -0.0086115 -0.0199368
+ 1.022e+11Hz -0.00863806 -0.0199374
+ 1.023e+11Hz -0.0086646 -0.019938
+ 1.024e+11Hz -0.00869113 -0.0199386
+ 1.025e+11Hz -0.00871763 -0.019939
+ 1.026e+11Hz -0.00874411 -0.0199395
+ 1.027e+11Hz -0.00877057 -0.0199399
+ 1.028e+11Hz -0.00879701 -0.0199402
+ 1.029e+11Hz -0.00882343 -0.0199405
+ 1.03e+11Hz -0.00884982 -0.0199407
+ 1.031e+11Hz -0.0088762 -0.0199409
+ 1.032e+11Hz -0.00890255 -0.019941
+ 1.033e+11Hz -0.00892888 -0.0199411
+ 1.034e+11Hz -0.00895519 -0.0199412
+ 1.035e+11Hz -0.00898148 -0.0199412
+ 1.036e+11Hz -0.00900775 -0.0199411
+ 1.037e+11Hz -0.00903399 -0.019941
+ 1.038e+11Hz -0.00906022 -0.0199408
+ 1.039e+11Hz -0.00908642 -0.0199406
+ 1.04e+11Hz -0.0091126 -0.0199404
+ 1.041e+11Hz -0.00913875 -0.0199401
+ 1.042e+11Hz -0.00916489 -0.0199397
+ 1.043e+11Hz -0.009191 -0.0199393
+ 1.044e+11Hz -0.00921709 -0.0199389
+ 1.045e+11Hz -0.00924315 -0.0199384
+ 1.046e+11Hz -0.0092692 -0.0199378
+ 1.047e+11Hz -0.00929522 -0.0199373
+ 1.048e+11Hz -0.00932122 -0.0199366
+ 1.049e+11Hz -0.00934719 -0.0199359
+ 1.05e+11Hz -0.00937315 -0.0199352
+ 1.051e+11Hz -0.00939908 -0.0199345
+ 1.052e+11Hz -0.00942498 -0.0199336
+ 1.053e+11Hz -0.00945087 -0.0199328
+ 1.054e+11Hz -0.00947673 -0.0199319
+ 1.055e+11Hz -0.00950257 -0.0199309
+ 1.056e+11Hz -0.00952838 -0.0199299
+ 1.057e+11Hz -0.00955417 -0.0199289
+ 1.058e+11Hz -0.00957994 -0.0199278
+ 1.059e+11Hz -0.00960569 -0.0199267
+ 1.06e+11Hz -0.00963141 -0.0199255
+ 1.061e+11Hz -0.00965711 -0.0199243
+ 1.062e+11Hz -0.00968279 -0.019923
+ 1.063e+11Hz -0.00970844 -0.0199217
+ 1.064e+11Hz -0.00973407 -0.0199203
+ 1.065e+11Hz -0.00975968 -0.0199189
+ 1.066e+11Hz -0.00978526 -0.0199175
+ 1.067e+11Hz -0.00981082 -0.019916
+ 1.068e+11Hz -0.00983636 -0.0199145
+ 1.069e+11Hz -0.00986187 -0.0199129
+ 1.07e+11Hz -0.00988736 -0.0199113
+ 1.071e+11Hz -0.00991283 -0.0199096
+ 1.072e+11Hz -0.00993828 -0.019908
+ 1.073e+11Hz -0.0099637 -0.0199062
+ 1.074e+11Hz -0.00998909 -0.0199044
+ 1.075e+11Hz -0.0100145 -0.0199026
+ 1.076e+11Hz -0.0100398 -0.0199007
+ 1.077e+11Hz -0.0100651 -0.0198988
+ 1.078e+11Hz -0.0100905 -0.0198969
+ 1.079e+11Hz -0.0101157 -0.0198949
+ 1.08e+11Hz -0.010141 -0.0198928
+ 1.081e+11Hz -0.0101662 -0.0198908
+ 1.082e+11Hz -0.0101914 -0.0198886
+ 1.083e+11Hz -0.0102166 -0.0198865
+ 1.084e+11Hz -0.0102418 -0.0198843
+ 1.085e+11Hz -0.0102669 -0.019882
+ 1.086e+11Hz -0.0102921 -0.0198797
+ 1.087e+11Hz -0.0103172 -0.0198774
+ 1.088e+11Hz -0.0103422 -0.019875
+ 1.089e+11Hz -0.0103673 -0.0198726
+ 1.09e+11Hz -0.0103923 -0.0198702
+ 1.091e+11Hz -0.0104173 -0.0198677
+ 1.092e+11Hz -0.0104423 -0.0198652
+ 1.093e+11Hz -0.0104672 -0.0198626
+ 1.094e+11Hz -0.0104922 -0.01986
+ 1.095e+11Hz -0.0105171 -0.0198573
+ 1.096e+11Hz -0.010542 -0.0198546
+ 1.097e+11Hz -0.0105668 -0.0198519
+ 1.098e+11Hz -0.0105917 -0.0198491
+ 1.099e+11Hz -0.0106165 -0.0198463
+ 1.1e+11Hz -0.0106413 -0.0198434
+ 1.101e+11Hz -0.0106661 -0.0198405
+ 1.102e+11Hz -0.0106908 -0.0198376
+ 1.103e+11Hz -0.0107155 -0.0198346
+ 1.104e+11Hz -0.0107403 -0.0198316
+ 1.105e+11Hz -0.0107649 -0.0198285
+ 1.106e+11Hz -0.0107896 -0.0198254
+ 1.107e+11Hz -0.0108142 -0.0198223
+ 1.108e+11Hz -0.0108388 -0.0198191
+ 1.109e+11Hz -0.0108634 -0.0198159
+ 1.11e+11Hz -0.010888 -0.0198126
+ 1.111e+11Hz -0.0109125 -0.0198093
+ 1.112e+11Hz -0.010937 -0.019806
+ 1.113e+11Hz -0.0109615 -0.0198026
+ 1.114e+11Hz -0.010986 -0.0197992
+ 1.115e+11Hz -0.0110105 -0.0197957
+ 1.116e+11Hz -0.0110349 -0.0197922
+ 1.117e+11Hz -0.0110593 -0.0197887
+ 1.118e+11Hz -0.0110837 -0.0197851
+ 1.119e+11Hz -0.011108 -0.0197815
+ 1.12e+11Hz -0.0111324 -0.0197778
+ 1.121e+11Hz -0.0111567 -0.0197741
+ 1.122e+11Hz -0.011181 -0.0197704
+ 1.123e+11Hz -0.0112052 -0.0197666
+ 1.124e+11Hz -0.0112295 -0.0197628
+ 1.125e+11Hz -0.0112537 -0.0197589
+ 1.126e+11Hz -0.0112779 -0.019755
+ 1.127e+11Hz -0.011302 -0.0197511
+ 1.128e+11Hz -0.0113262 -0.0197471
+ 1.129e+11Hz -0.0113503 -0.0197431
+ 1.13e+11Hz -0.0113744 -0.019739
+ 1.131e+11Hz -0.0113985 -0.0197349
+ 1.132e+11Hz -0.0114225 -0.0197308
+ 1.133e+11Hz -0.0114466 -0.0197266
+ 1.134e+11Hz -0.0114706 -0.0197224
+ 1.135e+11Hz -0.0114945 -0.0197181
+ 1.136e+11Hz -0.0115185 -0.0197138
+ 1.137e+11Hz -0.0115424 -0.0197095
+ 1.138e+11Hz -0.0115663 -0.0197051
+ 1.139e+11Hz -0.0115902 -0.0197007
+ 1.14e+11Hz -0.0116141 -0.0196962
+ 1.141e+11Hz -0.0116379 -0.0196917
+ 1.142e+11Hz -0.0116617 -0.0196872
+ 1.143e+11Hz -0.0116855 -0.0196826
+ 1.144e+11Hz -0.0117093 -0.019678
+ 1.145e+11Hz -0.011733 -0.0196733
+ 1.146e+11Hz -0.0117567 -0.0196686
+ 1.147e+11Hz -0.0117804 -0.0196638
+ 1.148e+11Hz -0.0118041 -0.0196591
+ 1.149e+11Hz -0.0118277 -0.0196542
+ 1.15e+11Hz -0.0118513 -0.0196494
+ 1.151e+11Hz -0.0118749 -0.0196445
+ 1.152e+11Hz -0.0118985 -0.0196395
+ 1.153e+11Hz -0.011922 -0.0196345
+ 1.154e+11Hz -0.0119455 -0.0196295
+ 1.155e+11Hz -0.011969 -0.0196245
+ 1.156e+11Hz -0.0119925 -0.0196194
+ 1.157e+11Hz -0.0120159 -0.0196142
+ 1.158e+11Hz -0.0120393 -0.019609
+ 1.159e+11Hz -0.0120627 -0.0196038
+ 1.16e+11Hz -0.012086 -0.0195985
+ 1.161e+11Hz -0.0121094 -0.0195932
+ 1.162e+11Hz -0.0121327 -0.0195879
+ 1.163e+11Hz -0.0121559 -0.0195825
+ 1.164e+11Hz -0.0121792 -0.019577
+ 1.165e+11Hz -0.0122024 -0.0195716
+ 1.166e+11Hz -0.0122256 -0.0195661
+ 1.167e+11Hz -0.0122488 -0.0195605
+ 1.168e+11Hz -0.0122719 -0.0195549
+ 1.169e+11Hz -0.012295 -0.0195493
+ 1.17e+11Hz -0.0123181 -0.0195436
+ 1.171e+11Hz -0.0123412 -0.0195379
+ 1.172e+11Hz -0.0123642 -0.0195322
+ 1.173e+11Hz -0.0123872 -0.0195264
+ 1.174e+11Hz -0.0124102 -0.0195205
+ 1.175e+11Hz -0.0124331 -0.0195147
+ 1.176e+11Hz -0.012456 -0.0195087
+ 1.177e+11Hz -0.0124789 -0.0195028
+ 1.178e+11Hz -0.0125018 -0.0194968
+ 1.179e+11Hz -0.0125246 -0.0194908
+ 1.18e+11Hz -0.0125474 -0.0194847
+ 1.181e+11Hz -0.0125702 -0.0194786
+ 1.182e+11Hz -0.0125929 -0.0194724
+ 1.183e+11Hz -0.0126157 -0.0194662
+ 1.184e+11Hz -0.0126383 -0.01946
+ 1.185e+11Hz -0.012661 -0.0194537
+ 1.186e+11Hz -0.0126836 -0.0194474
+ 1.187e+11Hz -0.0127062 -0.019441
+ 1.188e+11Hz -0.0127288 -0.0194346
+ 1.189e+11Hz -0.0127513 -0.0194282
+ 1.19e+11Hz -0.0127738 -0.0194217
+ 1.191e+11Hz -0.0127963 -0.0194152
+ 1.192e+11Hz -0.0128187 -0.0194086
+ 1.193e+11Hz -0.0128411 -0.019402
+ 1.194e+11Hz -0.0128635 -0.0193954
+ 1.195e+11Hz -0.0128859 -0.0193887
+ 1.196e+11Hz -0.0129082 -0.019382
+ 1.197e+11Hz -0.0129304 -0.0193752
+ 1.198e+11Hz -0.0129527 -0.0193684
+ 1.199e+11Hz -0.0129749 -0.0193616
+ 1.2e+11Hz -0.0129971 -0.0193547
+ 1.201e+11Hz -0.0130192 -0.0193478
+ 1.202e+11Hz -0.0130414 -0.0193409
+ 1.203e+11Hz -0.0130635 -0.0193339
+ 1.204e+11Hz -0.0130855 -0.0193268
+ 1.205e+11Hz -0.0131075 -0.0193198
+ 1.206e+11Hz -0.0131295 -0.0193126
+ 1.207e+11Hz -0.0131515 -0.0193055
+ 1.208e+11Hz -0.0131734 -0.0192983
+ 1.209e+11Hz -0.0131953 -0.0192911
+ 1.21e+11Hz -0.0132171 -0.0192838
+ 1.211e+11Hz -0.0132389 -0.0192765
+ 1.212e+11Hz -0.0132607 -0.0192692
+ 1.213e+11Hz -0.0132824 -0.0192618
+ 1.214e+11Hz -0.0133041 -0.0192544
+ 1.215e+11Hz -0.0133258 -0.0192469
+ 1.216e+11Hz -0.0133475 -0.0192394
+ 1.217e+11Hz -0.0133691 -0.0192319
+ 1.218e+11Hz -0.0133906 -0.0192243
+ 1.219e+11Hz -0.0134122 -0.0192167
+ 1.22e+11Hz -0.0134336 -0.019209
+ 1.221e+11Hz -0.0134551 -0.0192013
+ 1.222e+11Hz -0.0134765 -0.0191936
+ 1.223e+11Hz -0.0134979 -0.0191859
+ 1.224e+11Hz -0.0135192 -0.0191781
+ 1.225e+11Hz -0.0135405 -0.0191702
+ 1.226e+11Hz -0.0135618 -0.0191624
+ 1.227e+11Hz -0.013583 -0.0191544
+ 1.228e+11Hz -0.0136042 -0.0191465
+ 1.229e+11Hz -0.0136254 -0.0191385
+ 1.23e+11Hz -0.0136465 -0.0191305
+ 1.231e+11Hz -0.0136676 -0.0191225
+ 1.232e+11Hz -0.0136886 -0.0191144
+ 1.233e+11Hz -0.0137096 -0.0191062
+ 1.234e+11Hz -0.0137306 -0.0190981
+ 1.235e+11Hz -0.0137515 -0.0190899
+ 1.236e+11Hz -0.0137724 -0.0190816
+ 1.237e+11Hz -0.0137932 -0.0190734
+ 1.238e+11Hz -0.013814 -0.0190651
+ 1.239e+11Hz -0.0138348 -0.0190567
+ 1.24e+11Hz -0.0138555 -0.0190484
+ 1.241e+11Hz -0.0138762 -0.01904
+ 1.242e+11Hz -0.0138969 -0.0190315
+ 1.243e+11Hz -0.0139175 -0.019023
+ 1.244e+11Hz -0.013938 -0.0190145
+ 1.245e+11Hz -0.0139585 -0.019006
+ 1.246e+11Hz -0.013979 -0.0189974
+ 1.247e+11Hz -0.0139995 -0.0189888
+ 1.248e+11Hz -0.0140199 -0.0189802
+ 1.249e+11Hz -0.0140402 -0.0189715
+ 1.25e+11Hz -0.0140605 -0.0189628
+ 1.251e+11Hz -0.0140808 -0.018954
+ 1.252e+11Hz -0.014101 -0.0189452
+ 1.253e+11Hz -0.0141212 -0.0189364
+ 1.254e+11Hz -0.0141414 -0.0189276
+ 1.255e+11Hz -0.0141615 -0.0189187
+ 1.256e+11Hz -0.0141815 -0.0189098
+ 1.257e+11Hz -0.0142015 -0.0189009
+ 1.258e+11Hz -0.0142215 -0.0188919
+ 1.259e+11Hz -0.0142414 -0.0188829
+ 1.26e+11Hz -0.0142613 -0.0188739
+ 1.261e+11Hz -0.0142812 -0.0188648
+ 1.262e+11Hz -0.014301 -0.0188557
+ 1.263e+11Hz -0.0143207 -0.0188466
+ 1.264e+11Hz -0.0143404 -0.0188375
+ 1.265e+11Hz -0.0143601 -0.0188283
+ 1.266e+11Hz -0.0143797 -0.0188191
+ 1.267e+11Hz -0.0143993 -0.0188098
+ 1.268e+11Hz -0.0144188 -0.0188006
+ 1.269e+11Hz -0.0144383 -0.0187913
+ 1.27e+11Hz -0.0144578 -0.018782
+ 1.271e+11Hz -0.0144772 -0.0187726
+ 1.272e+11Hz -0.0144965 -0.0187632
+ 1.273e+11Hz -0.0145159 -0.0187538
+ 1.274e+11Hz -0.0145351 -0.0187444
+ 1.275e+11Hz -0.0145543 -0.0187349
+ 1.276e+11Hz -0.0145735 -0.0187254
+ 1.277e+11Hz -0.0145926 -0.0187159
+ 1.278e+11Hz -0.0146117 -0.0187063
+ 1.279e+11Hz -0.0146308 -0.0186968
+ 1.28e+11Hz -0.0146498 -0.0186872
+ 1.281e+11Hz -0.0146687 -0.0186775
+ 1.282e+11Hz -0.0146876 -0.0186679
+ 1.283e+11Hz -0.0147065 -0.0186582
+ 1.284e+11Hz -0.0147253 -0.0186485
+ 1.285e+11Hz -0.0147441 -0.0186388
+ 1.286e+11Hz -0.0147628 -0.018629
+ 1.287e+11Hz -0.0147814 -0.0186192
+ 1.288e+11Hz -0.0148001 -0.0186094
+ 1.289e+11Hz -0.0148186 -0.0185996
+ 1.29e+11Hz -0.0148372 -0.0185897
+ 1.291e+11Hz -0.0148557 -0.0185799
+ 1.292e+11Hz -0.0148741 -0.01857
+ 1.293e+11Hz -0.0148925 -0.01856
+ 1.294e+11Hz -0.0149108 -0.0185501
+ 1.295e+11Hz -0.0149291 -0.0185401
+ 1.296e+11Hz -0.0149474 -0.0185301
+ 1.297e+11Hz -0.0149656 -0.0185201
+ 1.298e+11Hz -0.0149838 -0.0185101
+ 1.299e+11Hz -0.0150019 -0.0185
+ 1.3e+11Hz -0.0150199 -0.0184899
+ 1.301e+11Hz -0.0150379 -0.0184798
+ 1.302e+11Hz -0.0150559 -0.0184697
+ 1.303e+11Hz -0.0150738 -0.0184595
+ 1.304e+11Hz -0.0150917 -0.0184494
+ 1.305e+11Hz -0.0151095 -0.0184392
+ 1.306e+11Hz -0.0151273 -0.018429
+ 1.307e+11Hz -0.015145 -0.0184187
+ 1.308e+11Hz -0.0151627 -0.0184085
+ 1.309e+11Hz -0.0151804 -0.0183982
+ 1.31e+11Hz -0.0151979 -0.0183879
+ 1.311e+11Hz -0.0152155 -0.0183776
+ 1.312e+11Hz -0.015233 -0.0183673
+ 1.313e+11Hz -0.0152504 -0.018357
+ 1.314e+11Hz -0.0152678 -0.0183466
+ 1.315e+11Hz -0.0152852 -0.0183362
+ 1.316e+11Hz -0.0153025 -0.0183258
+ 1.317e+11Hz -0.0153197 -0.0183154
+ 1.318e+11Hz -0.0153369 -0.018305
+ 1.319e+11Hz -0.0153541 -0.0182945
+ 1.32e+11Hz -0.0153712 -0.018284
+ 1.321e+11Hz -0.0153883 -0.0182735
+ 1.322e+11Hz -0.0154053 -0.018263
+ 1.323e+11Hz -0.0154222 -0.0182525
+ 1.324e+11Hz -0.0154392 -0.018242
+ 1.325e+11Hz -0.015456 -0.0182314
+ 1.326e+11Hz -0.0154729 -0.0182209
+ 1.327e+11Hz -0.0154896 -0.0182103
+ 1.328e+11Hz -0.0155064 -0.0181997
+ 1.329e+11Hz -0.015523 -0.0181891
+ 1.33e+11Hz -0.0155397 -0.0181784
+ 1.331e+11Hz -0.0155562 -0.0181678
+ 1.332e+11Hz -0.0155728 -0.0181571
+ 1.333e+11Hz -0.0155893 -0.0181464
+ 1.334e+11Hz -0.0156057 -0.0181358
+ 1.335e+11Hz -0.0156221 -0.0181251
+ 1.336e+11Hz -0.0156384 -0.0181143
+ 1.337e+11Hz -0.0156547 -0.0181036
+ 1.338e+11Hz -0.015671 -0.0180929
+ 1.339e+11Hz -0.0156872 -0.0180821
+ 1.34e+11Hz -0.0157033 -0.0180714
+ 1.341e+11Hz -0.0157194 -0.0180606
+ 1.342e+11Hz -0.0157355 -0.0180498
+ 1.343e+11Hz -0.0157515 -0.018039
+ 1.344e+11Hz -0.0157674 -0.0180282
+ 1.345e+11Hz -0.0157833 -0.0180173
+ 1.346e+11Hz -0.0157992 -0.0180065
+ 1.347e+11Hz -0.015815 -0.0179956
+ 1.348e+11Hz -0.0158308 -0.0179848
+ 1.349e+11Hz -0.0158465 -0.0179739
+ 1.35e+11Hz -0.0158622 -0.017963
+ 1.351e+11Hz -0.0158778 -0.0179521
+ 1.352e+11Hz -0.0158933 -0.0179412
+ 1.353e+11Hz -0.0159089 -0.0179303
+ 1.354e+11Hz -0.0159243 -0.0179194
+ 1.355e+11Hz -0.0159398 -0.0179084
+ 1.356e+11Hz -0.0159552 -0.0178975
+ 1.357e+11Hz -0.0159705 -0.0178865
+ 1.358e+11Hz -0.0159858 -0.0178756
+ 1.359e+11Hz -0.016001 -0.0178646
+ 1.36e+11Hz -0.0160162 -0.0178536
+ 1.361e+11Hz -0.0160313 -0.0178426
+ 1.362e+11Hz -0.0160464 -0.0178316
+ 1.363e+11Hz -0.0160615 -0.0178206
+ 1.364e+11Hz -0.0160765 -0.0178096
+ 1.365e+11Hz -0.0160914 -0.0177986
+ 1.366e+11Hz -0.0161063 -0.0177876
+ 1.367e+11Hz -0.0161212 -0.0177765
+ 1.368e+11Hz -0.016136 -0.0177655
+ 1.369e+11Hz -0.0161507 -0.0177544
+ 1.37e+11Hz -0.0161654 -0.0177434
+ 1.371e+11Hz -0.0161801 -0.0177323
+ 1.372e+11Hz -0.0161947 -0.0177212
+ 1.373e+11Hz -0.0162093 -0.0177101
+ 1.374e+11Hz -0.0162238 -0.0176991
+ 1.375e+11Hz -0.0162383 -0.017688
+ 1.376e+11Hz -0.0162527 -0.0176769
+ 1.377e+11Hz -0.0162671 -0.0176658
+ 1.378e+11Hz -0.0162814 -0.0176547
+ 1.379e+11Hz -0.0162957 -0.0176436
+ 1.38e+11Hz -0.0163099 -0.0176324
+ 1.381e+11Hz -0.0163241 -0.0176213
+ 1.382e+11Hz -0.0163382 -0.0176102
+ 1.383e+11Hz -0.0163523 -0.0175991
+ 1.384e+11Hz -0.0163663 -0.0175879
+ 1.385e+11Hz -0.0163803 -0.0175768
+ 1.386e+11Hz -0.0163943 -0.0175656
+ 1.387e+11Hz -0.0164082 -0.0175545
+ 1.388e+11Hz -0.016422 -0.0175433
+ 1.389e+11Hz -0.0164358 -0.0175322
+ 1.39e+11Hz -0.0164495 -0.017521
+ 1.391e+11Hz -0.0164633 -0.0175099
+ 1.392e+11Hz -0.0164769 -0.0174987
+ 1.393e+11Hz -0.0164905 -0.0174875
+ 1.394e+11Hz -0.0165041 -0.0174764
+ 1.395e+11Hz -0.0165176 -0.0174652
+ 1.396e+11Hz -0.016531 -0.017454
+ 1.397e+11Hz -0.0165445 -0.0174429
+ 1.398e+11Hz -0.0165578 -0.0174317
+ 1.399e+11Hz -0.0165711 -0.0174205
+ 1.4e+11Hz -0.0165844 -0.0174093
+ 1.401e+11Hz -0.0165976 -0.0173981
+ 1.402e+11Hz -0.0166108 -0.017387
+ 1.403e+11Hz -0.0166239 -0.0173758
+ 1.404e+11Hz -0.016637 -0.0173646
+ 1.405e+11Hz -0.0166501 -0.0173534
+ 1.406e+11Hz -0.016663 -0.0173422
+ 1.407e+11Hz -0.016676 -0.017331
+ 1.408e+11Hz -0.0166889 -0.0173199
+ 1.409e+11Hz -0.0167017 -0.0173087
+ 1.41e+11Hz -0.0167145 -0.0172975
+ 1.411e+11Hz -0.0167272 -0.0172863
+ 1.412e+11Hz -0.0167399 -0.0172751
+ 1.413e+11Hz -0.0167526 -0.017264
+ 1.414e+11Hz -0.0167652 -0.0172528
+ 1.415e+11Hz -0.0167777 -0.0172416
+ 1.416e+11Hz -0.0167902 -0.0172304
+ 1.417e+11Hz -0.0168027 -0.0172193
+ 1.418e+11Hz -0.0168151 -0.0172081
+ 1.419e+11Hz -0.0168274 -0.0171969
+ 1.42e+11Hz -0.0168398 -0.0171858
+ 1.421e+11Hz -0.016852 -0.0171746
+ 1.422e+11Hz -0.0168642 -0.0171634
+ 1.423e+11Hz -0.0168764 -0.0171523
+ 1.424e+11Hz -0.0168885 -0.0171411
+ 1.425e+11Hz -0.0169006 -0.01713
+ 1.426e+11Hz -0.0169126 -0.0171189
+ 1.427e+11Hz -0.0169246 -0.0171077
+ 1.428e+11Hz -0.0169365 -0.0170966
+ 1.429e+11Hz -0.0169484 -0.0170855
+ 1.43e+11Hz -0.0169602 -0.0170743
+ 1.431e+11Hz -0.016972 -0.0170632
+ 1.432e+11Hz -0.0169837 -0.0170521
+ 1.433e+11Hz -0.0169954 -0.017041
+ 1.434e+11Hz -0.017007 -0.0170299
+ 1.435e+11Hz -0.0170186 -0.0170188
+ 1.436e+11Hz -0.0170301 -0.0170077
+ 1.437e+11Hz -0.0170416 -0.0169966
+ 1.438e+11Hz -0.017053 -0.0169856
+ 1.439e+11Hz -0.0170644 -0.0169745
+ 1.44e+11Hz -0.0170757 -0.0169634
+ 1.441e+11Hz -0.017087 -0.0169524
+ 1.442e+11Hz -0.0170983 -0.0169413
+ 1.443e+11Hz -0.0171094 -0.0169303
+ 1.444e+11Hz -0.0171206 -0.0169193
+ 1.445e+11Hz -0.0171317 -0.0169083
+ 1.446e+11Hz -0.0171427 -0.0168973
+ 1.447e+11Hz -0.0171537 -0.0168863
+ 1.448e+11Hz -0.0171646 -0.0168753
+ 1.449e+11Hz -0.0171755 -0.0168643
+ 1.45e+11Hz -0.0171864 -0.0168533
+ 1.451e+11Hz -0.0171972 -0.0168424
+ 1.452e+11Hz -0.0172079 -0.0168314
+ 1.453e+11Hz -0.0172186 -0.0168205
+ 1.454e+11Hz -0.0172293 -0.0168096
+ 1.455e+11Hz -0.0172399 -0.0167987
+ 1.456e+11Hz -0.0172504 -0.0167878
+ 1.457e+11Hz -0.0172609 -0.0167769
+ 1.458e+11Hz -0.0172714 -0.016766
+ 1.459e+11Hz -0.0172818 -0.0167551
+ 1.46e+11Hz -0.0172921 -0.0167443
+ 1.461e+11Hz -0.0173024 -0.0167335
+ 1.462e+11Hz -0.0173127 -0.0167227
+ 1.463e+11Hz -0.0173229 -0.0167119
+ 1.464e+11Hz -0.017333 -0.0167011
+ 1.465e+11Hz -0.0173432 -0.0166903
+ 1.466e+11Hz -0.0173532 -0.0166795
+ 1.467e+11Hz -0.0173632 -0.0166688
+ 1.468e+11Hz -0.0173732 -0.0166581
+ 1.469e+11Hz -0.0173831 -0.0166474
+ 1.47e+11Hz -0.017393 -0.0166367
+ 1.471e+11Hz -0.0174028 -0.016626
+ 1.472e+11Hz -0.0174125 -0.0166154
+ 1.473e+11Hz -0.0174222 -0.0166047
+ 1.474e+11Hz -0.0174319 -0.0165941
+ 1.475e+11Hz -0.0174415 -0.0165835
+ 1.476e+11Hz -0.0174511 -0.0165729
+ 1.477e+11Hz -0.0174606 -0.0165624
+ 1.478e+11Hz -0.0174701 -0.0165518
+ 1.479e+11Hz -0.0174795 -0.0165413
+ 1.48e+11Hz -0.0174889 -0.0165308
+ 1.481e+11Hz -0.0174982 -0.0165203
+ 1.482e+11Hz -0.0175074 -0.0165099
+ 1.483e+11Hz -0.0175167 -0.0164994
+ 1.484e+11Hz -0.0175258 -0.016489
+ 1.485e+11Hz -0.017535 -0.0164787
+ 1.486e+11Hz -0.0175441 -0.0164683
+ 1.487e+11Hz -0.0175531 -0.0164579
+ 1.488e+11Hz -0.0175621 -0.0164476
+ 1.489e+11Hz -0.017571 -0.0164373
+ 1.49e+11Hz -0.0175799 -0.0164271
+ 1.491e+11Hz -0.0175887 -0.0164168
+ 1.492e+11Hz -0.0175975 -0.0164066
+ 1.493e+11Hz -0.0176063 -0.0163964
+ 1.494e+11Hz -0.0176149 -0.0163863
+ 1.495e+11Hz -0.0176236 -0.0163762
+ 1.496e+11Hz -0.0176322 -0.016366
+ 1.497e+11Hz -0.0176407 -0.016356
+ 1.498e+11Hz -0.0176492 -0.0163459
+ 1.499e+11Hz -0.0176577 -0.0163359
+ 1.5e+11Hz -0.0176661 -0.0163259
+ 1.501e+11Hz -0.0176745 -0.016316
+ 1.502e+11Hz -0.0176828 -0.016306
+ 1.503e+11Hz -0.0176911 -0.0162961
+ 1.504e+11Hz -0.0176993 -0.0162863
+ 1.505e+11Hz -0.0177075 -0.0162764
+ 1.506e+11Hz -0.0177156 -0.0162666
+ 1.507e+11Hz -0.0177237 -0.0162569
+ 1.508e+11Hz -0.0177317 -0.0162471
+ 1.509e+11Hz -0.0177397 -0.0162374
+ 1.51e+11Hz -0.0177477 -0.0162278
+ 1.511e+11Hz -0.0177556 -0.0162181
+ 1.512e+11Hz -0.0177634 -0.0162085
+ 1.513e+11Hz -0.0177713 -0.016199
+ 1.514e+11Hz -0.017779 -0.0161895
+ 1.515e+11Hz -0.0177868 -0.01618
+ 1.516e+11Hz -0.0177944 -0.0161705
+ 1.517e+11Hz -0.0178021 -0.0161611
+ 1.518e+11Hz -0.0178097 -0.0161518
+ 1.519e+11Hz -0.0178172 -0.0161424
+ 1.52e+11Hz -0.0178247 -0.0161331
+ 1.521e+11Hz -0.0178322 -0.0161239
+ 1.522e+11Hz -0.0178396 -0.0161147
+ 1.523e+11Hz -0.017847 -0.0161055
+ 1.524e+11Hz -0.0178544 -0.0160964
+ 1.525e+11Hz -0.0178617 -0.0160873
+ 1.526e+11Hz -0.0178689 -0.0160782
+ 1.527e+11Hz -0.0178762 -0.0160692
+ 1.528e+11Hz -0.0178833 -0.0160603
+ 1.529e+11Hz -0.0178905 -0.0160513
+ 1.53e+11Hz -0.0178976 -0.0160425
+ 1.531e+11Hz -0.0179046 -0.0160336
+ 1.532e+11Hz -0.0179117 -0.0160249
+ 1.533e+11Hz -0.0179187 -0.0160161
+ 1.534e+11Hz -0.0179256 -0.0160074
+ 1.535e+11Hz -0.0179325 -0.0159988
+ 1.536e+11Hz -0.0179394 -0.0159902
+ 1.537e+11Hz -0.0179462 -0.0159817
+ 1.538e+11Hz -0.017953 -0.0159732
+ 1.539e+11Hz -0.0179598 -0.0159647
+ 1.54e+11Hz -0.0179665 -0.0159563
+ 1.541e+11Hz -0.0179732 -0.015948
+ 1.542e+11Hz -0.0179799 -0.0159397
+ 1.543e+11Hz -0.0179865 -0.0159314
+ 1.544e+11Hz -0.0179931 -0.0159232
+ 1.545e+11Hz -0.0179996 -0.0159151
+ 1.546e+11Hz -0.0180062 -0.015907
+ 1.547e+11Hz -0.0180126 -0.0158989
+ 1.548e+11Hz -0.0180191 -0.0158909
+ 1.549e+11Hz -0.0180255 -0.015883
+ 1.55e+11Hz -0.0180319 -0.0158751
+ 1.551e+11Hz -0.0180383 -0.0158673
+ 1.552e+11Hz -0.0180446 -0.0158595
+ 1.553e+11Hz -0.0180509 -0.0158518
+ 1.554e+11Hz -0.0180572 -0.0158442
+ 1.555e+11Hz -0.0180635 -0.0158366
+ 1.556e+11Hz -0.0180697 -0.015829
+ 1.557e+11Hz -0.0180759 -0.0158215
+ 1.558e+11Hz -0.0180821 -0.0158141
+ 1.559e+11Hz -0.0180882 -0.0158067
+ 1.56e+11Hz -0.0180943 -0.0157994
+ 1.561e+11Hz -0.0181004 -0.0157922
+ 1.562e+11Hz -0.0181065 -0.015785
+ 1.563e+11Hz -0.0181126 -0.0157779
+ 1.564e+11Hz -0.0181186 -0.0157708
+ 1.565e+11Hz -0.0181246 -0.0157638
+ 1.566e+11Hz -0.0181306 -0.0157568
+ 1.567e+11Hz -0.0181365 -0.0157499
+ 1.568e+11Hz -0.0181425 -0.0157431
+ 1.569e+11Hz -0.0181484 -0.0157364
+ 1.57e+11Hz -0.0181543 -0.0157297
+ 1.571e+11Hz -0.0181602 -0.015723
+ 1.572e+11Hz -0.0181661 -0.0157164
+ 1.573e+11Hz -0.0181719 -0.0157099
+ 1.574e+11Hz -0.0181778 -0.0157035
+ 1.575e+11Hz -0.0181836 -0.0156971
+ 1.576e+11Hz -0.0181894 -0.0156908
+ 1.577e+11Hz -0.0181952 -0.0156845
+ 1.578e+11Hz -0.018201 -0.0156784
+ 1.579e+11Hz -0.0182068 -0.0156722
+ 1.58e+11Hz -0.0182125 -0.0156662
+ 1.581e+11Hz -0.0182183 -0.0156602
+ 1.582e+11Hz -0.018224 -0.0156543
+ 1.583e+11Hz -0.0182298 -0.0156484
+ 1.584e+11Hz -0.0182355 -0.0156427
+ 1.585e+11Hz -0.0182412 -0.0156369
+ 1.586e+11Hz -0.0182469 -0.0156313
+ 1.587e+11Hz -0.0182526 -0.0156257
+ 1.588e+11Hz -0.0182583 -0.0156202
+ 1.589e+11Hz -0.018264 -0.0156148
+ 1.59e+11Hz -0.0182697 -0.0156094
+ 1.591e+11Hz -0.0182754 -0.0156041
+ 1.592e+11Hz -0.0182811 -0.0155988
+ 1.593e+11Hz -0.0182868 -0.0155937
+ 1.594e+11Hz -0.0182925 -0.0155886
+ 1.595e+11Hz -0.0182982 -0.0155835
+ 1.596e+11Hz -0.0183039 -0.0155786
+ 1.597e+11Hz -0.0183096 -0.0155737
+ 1.598e+11Hz -0.0183153 -0.0155689
+ 1.599e+11Hz -0.018321 -0.0155641
+ 1.6e+11Hz -0.0183267 -0.0155595
+ 1.601e+11Hz -0.0183325 -0.0155549
+ 1.602e+11Hz -0.0183382 -0.0155503
+ 1.603e+11Hz -0.0183439 -0.0155459
+ 1.604e+11Hz -0.0183497 -0.0155415
+ 1.605e+11Hz -0.0183555 -0.0155371
+ 1.606e+11Hz -0.0183612 -0.0155329
+ 1.607e+11Hz -0.018367 -0.0155287
+ 1.608e+11Hz -0.0183728 -0.0155246
+ 1.609e+11Hz -0.0183786 -0.0155206
+ 1.61e+11Hz -0.0183845 -0.0155166
+ 1.611e+11Hz -0.0183903 -0.0155127
+ 1.612e+11Hz -0.0183962 -0.0155089
+ 1.613e+11Hz -0.0184021 -0.0155051
+ 1.614e+11Hz -0.018408 -0.0155014
+ 1.615e+11Hz -0.0184139 -0.0154978
+ 1.616e+11Hz -0.0184199 -0.0154943
+ 1.617e+11Hz -0.0184258 -0.0154908
+ 1.618e+11Hz -0.0184318 -0.0154874
+ 1.619e+11Hz -0.0184378 -0.0154841
+ 1.62e+11Hz -0.0184439 -0.0154808
+ 1.621e+11Hz -0.0184499 -0.0154776
+ 1.622e+11Hz -0.018456 -0.0154745
+ 1.623e+11Hz -0.0184622 -0.0154714
+ 1.624e+11Hz -0.0184683 -0.0154684
+ 1.625e+11Hz -0.0184745 -0.0154655
+ 1.626e+11Hz -0.0184807 -0.0154627
+ 1.627e+11Hz -0.018487 -0.0154599
+ 1.628e+11Hz -0.0184933 -0.0154572
+ 1.629e+11Hz -0.0184996 -0.0154546
+ 1.63e+11Hz -0.0185059 -0.015452
+ 1.631e+11Hz -0.0185123 -0.0154495
+ 1.632e+11Hz -0.0185187 -0.0154471
+ 1.633e+11Hz -0.0185252 -0.0154447
+ 1.634e+11Hz -0.0185317 -0.0154424
+ 1.635e+11Hz -0.0185383 -0.0154402
+ 1.636e+11Hz -0.0185448 -0.015438
+ 1.637e+11Hz -0.0185515 -0.0154359
+ 1.638e+11Hz -0.0185582 -0.0154339
+ 1.639e+11Hz -0.0185649 -0.0154319
+ 1.64e+11Hz -0.0185716 -0.01543
+ 1.641e+11Hz -0.0185785 -0.0154281
+ 1.642e+11Hz -0.0185853 -0.0154264
+ 1.643e+11Hz -0.0185922 -0.0154247
+ 1.644e+11Hz -0.0185992 -0.015423
+ 1.645e+11Hz -0.0186062 -0.0154214
+ 1.646e+11Hz -0.0186132 -0.0154199
+ 1.647e+11Hz -0.0186204 -0.0154184
+ 1.648e+11Hz -0.0186275 -0.015417
+ 1.649e+11Hz -0.0186347 -0.0154157
+ 1.65e+11Hz -0.018642 -0.0154144
+ 1.651e+11Hz -0.0186494 -0.0154132
+ 1.652e+11Hz -0.0186567 -0.015412
+ 1.653e+11Hz -0.0186642 -0.0154109
+ 1.654e+11Hz -0.0186717 -0.0154098
+ 1.655e+11Hz -0.0186793 -0.0154088
+ 1.656e+11Hz -0.0186869 -0.0154079
+ 1.657e+11Hz -0.0186946 -0.015407
+ 1.658e+11Hz -0.0187023 -0.0154062
+ 1.659e+11Hz -0.0187102 -0.0154054
+ 1.66e+11Hz -0.0187181 -0.0154047
+ 1.661e+11Hz -0.018726 -0.015404
+ 1.662e+11Hz -0.018734 -0.0154034
+ 1.663e+11Hz -0.0187421 -0.0154028
+ 1.664e+11Hz -0.0187503 -0.0154023
+ 1.665e+11Hz -0.0187585 -0.0154018
+ 1.666e+11Hz -0.0187668 -0.0154014
+ 1.667e+11Hz -0.0187751 -0.0154011
+ 1.668e+11Hz -0.0187836 -0.0154007
+ 1.669e+11Hz -0.0187921 -0.0154005
+ 1.67e+11Hz -0.0188007 -0.0154002
+ 1.671e+11Hz -0.0188093 -0.0154
+ 1.672e+11Hz -0.0188181 -0.0153999
+ 1.673e+11Hz -0.0188269 -0.0153998
+ 1.674e+11Hz -0.0188358 -0.0153997
+ 1.675e+11Hz -0.0188447 -0.0153997
+ 1.676e+11Hz -0.0188538 -0.0153997
+ 1.677e+11Hz -0.0188629 -0.0153998
+ 1.678e+11Hz -0.0188721 -0.0153999
+ 1.679e+11Hz -0.0188814 -0.0154
+ 1.68e+11Hz -0.0188908 -0.0154002
+ 1.681e+11Hz -0.0189002 -0.0154004
+ 1.682e+11Hz -0.0189097 -0.0154007
+ 1.683e+11Hz -0.0189194 -0.015401
+ 1.684e+11Hz -0.0189291 -0.0154013
+ 1.685e+11Hz -0.0189388 -0.0154016
+ 1.686e+11Hz -0.0189487 -0.015402
+ 1.687e+11Hz -0.0189587 -0.0154024
+ 1.688e+11Hz -0.0189687 -0.0154028
+ 1.689e+11Hz -0.0189789 -0.0154033
+ 1.69e+11Hz -0.0189891 -0.0154037
+ 1.691e+11Hz -0.0189994 -0.0154043
+ 1.692e+11Hz -0.0190098 -0.0154048
+ 1.693e+11Hz -0.0190203 -0.0154053
+ 1.694e+11Hz -0.0190309 -0.0154059
+ 1.695e+11Hz -0.0190415 -0.0154065
+ 1.696e+11Hz -0.0190523 -0.0154071
+ 1.697e+11Hz -0.0190632 -0.0154078
+ 1.698e+11Hz -0.0190741 -0.0154084
+ 1.699e+11Hz -0.0190852 -0.0154091
+ 1.7e+11Hz -0.0190963 -0.0154098
+ 1.701e+11Hz -0.0191075 -0.0154105
+ 1.702e+11Hz -0.0191189 -0.0154112
+ 1.703e+11Hz -0.0191303 -0.0154119
+ 1.704e+11Hz -0.0191418 -0.0154126
+ 1.705e+11Hz -0.0191534 -0.0154133
+ 1.706e+11Hz -0.0191651 -0.0154141
+ 1.707e+11Hz -0.0191769 -0.0154148
+ 1.708e+11Hz -0.0191889 -0.0154156
+ 1.709e+11Hz -0.0192009 -0.0154163
+ 1.71e+11Hz -0.019213 -0.0154171
+ 1.711e+11Hz -0.0192252 -0.0154179
+ 1.712e+11Hz -0.0192375 -0.0154186
+ 1.713e+11Hz -0.0192499 -0.0154194
+ 1.714e+11Hz -0.0192623 -0.0154201
+ 1.715e+11Hz -0.0192749 -0.0154209
+ 1.716e+11Hz -0.0192876 -0.0154216
+ 1.717e+11Hz -0.0193004 -0.0154224
+ 1.718e+11Hz -0.0193133 -0.0154231
+ 1.719e+11Hz -0.0193263 -0.0154238
+ 1.72e+11Hz -0.0193394 -0.0154246
+ 1.721e+11Hz -0.0193526 -0.0154253
+ 1.722e+11Hz -0.0193659 -0.015426
+ 1.723e+11Hz -0.0193793 -0.0154266
+ 1.724e+11Hz -0.0193928 -0.0154273
+ 1.725e+11Hz -0.0194064 -0.0154279
+ 1.726e+11Hz -0.0194201 -0.0154285
+ 1.727e+11Hz -0.0194339 -0.0154292
+ 1.728e+11Hz -0.0194478 -0.0154297
+ 1.729e+11Hz -0.0194618 -0.0154303
+ 1.73e+11Hz -0.0194759 -0.0154308
+ 1.731e+11Hz -0.0194901 -0.0154313
+ 1.732e+11Hz -0.0195044 -0.0154318
+ 1.733e+11Hz -0.0195188 -0.0154323
+ 1.734e+11Hz -0.0195334 -0.0154327
+ 1.735e+11Hz -0.019548 -0.0154331
+ 1.736e+11Hz -0.0195627 -0.0154335
+ 1.737e+11Hz -0.0195775 -0.0154338
+ 1.738e+11Hz -0.0195924 -0.0154341
+ 1.739e+11Hz -0.0196074 -0.0154343
+ 1.74e+11Hz -0.0196225 -0.0154346
+ 1.741e+11Hz -0.0196377 -0.0154348
+ 1.742e+11Hz -0.019653 -0.0154349
+ 1.743e+11Hz -0.0196684 -0.015435
+ 1.744e+11Hz -0.0196839 -0.0154351
+ 1.745e+11Hz -0.0196995 -0.0154351
+ 1.746e+11Hz -0.0197153 -0.015435
+ 1.747e+11Hz -0.0197311 -0.015435
+ 1.748e+11Hz -0.019747 -0.0154348
+ 1.749e+11Hz -0.019763 -0.0154347
+ 1.75e+11Hz -0.019779 -0.0154344
+ 1.751e+11Hz -0.0197952 -0.0154342
+ 1.752e+11Hz -0.0198115 -0.0154338
+ 1.753e+11Hz -0.0198279 -0.0154335
+ 1.754e+11Hz -0.0198444 -0.015433
+ 1.755e+11Hz -0.019861 -0.0154325
+ 1.756e+11Hz -0.0198776 -0.015432
+ 1.757e+11Hz -0.0198944 -0.0154313
+ 1.758e+11Hz -0.0199112 -0.0154307
+ 1.759e+11Hz -0.0199282 -0.0154299
+ 1.76e+11Hz -0.0199452 -0.0154291
+ 1.761e+11Hz -0.0199624 -0.0154283
+ 1.762e+11Hz -0.0199796 -0.0154273
+ 1.763e+11Hz -0.0199969 -0.0154263
+ 1.764e+11Hz -0.0200143 -0.0154252
+ 1.765e+11Hz -0.0200318 -0.0154241
+ 1.766e+11Hz -0.0200494 -0.0154229
+ 1.767e+11Hz -0.020067 -0.0154216
+ 1.768e+11Hz -0.0200848 -0.0154202
+ 1.769e+11Hz -0.0201026 -0.0154188
+ 1.77e+11Hz -0.0201206 -0.0154173
+ 1.771e+11Hz -0.0201386 -0.0154157
+ 1.772e+11Hz -0.0201567 -0.015414
+ 1.773e+11Hz -0.0201749 -0.0154123
+ 1.774e+11Hz -0.0201931 -0.0154105
+ 1.775e+11Hz -0.0202115 -0.0154086
+ 1.776e+11Hz -0.0202299 -0.0154066
+ 1.777e+11Hz -0.0202484 -0.0154045
+ 1.778e+11Hz -0.020267 -0.0154023
+ 1.779e+11Hz -0.0202857 -0.0154001
+ 1.78e+11Hz -0.0203044 -0.0153977
+ 1.781e+11Hz -0.0203232 -0.0153953
+ 1.782e+11Hz -0.0203421 -0.0153928
+ 1.783e+11Hz -0.0203611 -0.0153902
+ 1.784e+11Hz -0.0203801 -0.0153875
+ 1.785e+11Hz -0.0203993 -0.0153847
+ 1.786e+11Hz -0.0204184 -0.0153818
+ 1.787e+11Hz -0.0204377 -0.0153788
+ 1.788e+11Hz -0.020457 -0.0153757
+ 1.789e+11Hz -0.0204764 -0.0153726
+ 1.79e+11Hz -0.0204959 -0.0153693
+ 1.791e+11Hz -0.0205154 -0.0153659
+ 1.792e+11Hz -0.020535 -0.0153624
+ 1.793e+11Hz -0.0205547 -0.0153589
+ 1.794e+11Hz -0.0205744 -0.0153552
+ 1.795e+11Hz -0.0205942 -0.0153514
+ 1.796e+11Hz -0.0206141 -0.0153475
+ 1.797e+11Hz -0.020634 -0.0153435
+ 1.798e+11Hz -0.020654 -0.0153394
+ 1.799e+11Hz -0.020674 -0.0153352
+ 1.8e+11Hz -0.0206941 -0.0153309
+ 1.801e+11Hz -0.0207143 -0.0153265
+ 1.802e+11Hz -0.0207345 -0.015322
+ 1.803e+11Hz -0.0207547 -0.0153174
+ 1.804e+11Hz -0.020775 -0.0153126
+ 1.805e+11Hz -0.0207954 -0.0153078
+ 1.806e+11Hz -0.0208158 -0.0153028
+ 1.807e+11Hz -0.0208363 -0.0152977
+ 1.808e+11Hz -0.0208568 -0.0152925
+ 1.809e+11Hz -0.0208773 -0.0152872
+ 1.81e+11Hz -0.0208979 -0.0152818
+ 1.811e+11Hz -0.0209186 -0.0152762
+ 1.812e+11Hz -0.0209392 -0.0152706
+ 1.813e+11Hz -0.02096 -0.0152648
+ 1.814e+11Hz -0.0209807 -0.0152589
+ 1.815e+11Hz -0.0210015 -0.0152529
+ 1.816e+11Hz -0.0210224 -0.0152467
+ 1.817e+11Hz -0.0210433 -0.0152405
+ 1.818e+11Hz -0.0210642 -0.0152341
+ 1.819e+11Hz -0.0210851 -0.0152276
+ 1.82e+11Hz -0.0211061 -0.015221
+ 1.821e+11Hz -0.0211271 -0.0152143
+ 1.822e+11Hz -0.0211481 -0.0152074
+ 1.823e+11Hz -0.0211692 -0.0152004
+ 1.824e+11Hz -0.0211903 -0.0151933
+ 1.825e+11Hz -0.0212114 -0.0151861
+ 1.826e+11Hz -0.0212325 -0.0151787
+ 1.827e+11Hz -0.0212537 -0.0151712
+ 1.828e+11Hz -0.0212749 -0.0151636
+ 1.829e+11Hz -0.0212961 -0.0151559
+ 1.83e+11Hz -0.0213173 -0.015148
+ 1.831e+11Hz -0.0213385 -0.0151401
+ 1.832e+11Hz -0.0213598 -0.015132
+ 1.833e+11Hz -0.021381 -0.0151237
+ 1.834e+11Hz -0.0214023 -0.0151154
+ 1.835e+11Hz -0.0214236 -0.0151069
+ 1.836e+11Hz -0.0214449 -0.0150982
+ 1.837e+11Hz -0.0214662 -0.0150895
+ 1.838e+11Hz -0.0214875 -0.0150806
+ 1.839e+11Hz -0.0215088 -0.0150716
+ 1.84e+11Hz -0.0215301 -0.0150625
+ 1.841e+11Hz -0.0215515 -0.0150532
+ 1.842e+11Hz -0.0215728 -0.0150438
+ 1.843e+11Hz -0.0215941 -0.0150343
+ 1.844e+11Hz -0.0216154 -0.0150247
+ 1.845e+11Hz -0.0216367 -0.0150149
+ 1.846e+11Hz -0.021658 -0.015005
+ 1.847e+11Hz -0.0216793 -0.014995
+ 1.848e+11Hz -0.0217006 -0.0149848
+ 1.849e+11Hz -0.0217219 -0.0149745
+ 1.85e+11Hz -0.0217432 -0.0149641
+ 1.851e+11Hz -0.0217644 -0.0149536
+ 1.852e+11Hz -0.0217857 -0.0149429
+ 1.853e+11Hz -0.0218069 -0.0149321
+ 1.854e+11Hz -0.0218281 -0.0149212
+ 1.855e+11Hz -0.0218493 -0.0149101
+ 1.856e+11Hz -0.0218705 -0.0148989
+ 1.857e+11Hz -0.0218916 -0.0148876
+ 1.858e+11Hz -0.0219128 -0.0148761
+ 1.859e+11Hz -0.0219339 -0.0148646
+ 1.86e+11Hz -0.0219549 -0.0148529
+ 1.861e+11Hz -0.021976 -0.014841
+ 1.862e+11Hz -0.021997 -0.0148291
+ 1.863e+11Hz -0.022018 -0.014817
+ 1.864e+11Hz -0.022039 -0.0148048
+ 1.865e+11Hz -0.0220599 -0.0147925
+ 1.866e+11Hz -0.0220808 -0.01478
+ 1.867e+11Hz -0.0221016 -0.0147674
+ 1.868e+11Hz -0.0221224 -0.0147547
+ 1.869e+11Hz -0.0221432 -0.0147419
+ 1.87e+11Hz -0.0221639 -0.0147289
+ 1.871e+11Hz -0.0221846 -0.0147158
+ 1.872e+11Hz -0.0222053 -0.0147026
+ 1.873e+11Hz -0.0222259 -0.0146893
+ 1.874e+11Hz -0.0222464 -0.0146758
+ 1.875e+11Hz -0.0222669 -0.0146623
+ 1.876e+11Hz -0.0222874 -0.0146486
+ 1.877e+11Hz -0.0223078 -0.0146348
+ 1.878e+11Hz -0.0223282 -0.0146208
+ 1.879e+11Hz -0.0223485 -0.0146068
+ 1.88e+11Hz -0.0223687 -0.0145926
+ 1.881e+11Hz -0.0223889 -0.0145783
+ 1.882e+11Hz -0.022409 -0.0145639
+ 1.883e+11Hz -0.0224291 -0.0145494
+ 1.884e+11Hz -0.0224491 -0.0145347
+ 1.885e+11Hz -0.0224691 -0.01452
+ 1.886e+11Hz -0.022489 -0.0145051
+ 1.887e+11Hz -0.0225088 -0.0144901
+ 1.888e+11Hz -0.0225286 -0.014475
+ 1.889e+11Hz -0.0225482 -0.0144598
+ 1.89e+11Hz -0.0225679 -0.0144445
+ 1.891e+11Hz -0.0225874 -0.0144291
+ 1.892e+11Hz -0.0226069 -0.0144135
+ 1.893e+11Hz -0.0226263 -0.0143979
+ 1.894e+11Hz -0.0226457 -0.0143821
+ 1.895e+11Hz -0.0226649 -0.0143663
+ 1.896e+11Hz -0.0226841 -0.0143503
+ 1.897e+11Hz -0.0227032 -0.0143342
+ 1.898e+11Hz -0.0227223 -0.014318
+ 1.899e+11Hz -0.0227412 -0.0143017
+ 1.9e+11Hz -0.0227601 -0.0142854
+ 1.901e+11Hz -0.0227789 -0.0142689
+ 1.902e+11Hz -0.0227976 -0.0142523
+ 1.903e+11Hz -0.0228162 -0.0142356
+ 1.904e+11Hz -0.0228348 -0.0142188
+ 1.905e+11Hz -0.0228532 -0.0142019
+ 1.906e+11Hz -0.0228716 -0.014185
+ 1.907e+11Hz -0.0228899 -0.0141679
+ 1.908e+11Hz -0.0229081 -0.0141507
+ 1.909e+11Hz -0.0229262 -0.0141335
+ 1.91e+11Hz -0.0229442 -0.0141161
+ 1.911e+11Hz -0.0229621 -0.0140987
+ 1.912e+11Hz -0.0229799 -0.0140812
+ 1.913e+11Hz -0.0229976 -0.0140635
+ 1.914e+11Hz -0.0230153 -0.0140458
+ 1.915e+11Hz -0.0230328 -0.014028
+ 1.916e+11Hz -0.0230503 -0.0140102
+ 1.917e+11Hz -0.0230676 -0.0139922
+ 1.918e+11Hz -0.0230848 -0.0139742
+ 1.919e+11Hz -0.023102 -0.0139561
+ 1.92e+11Hz -0.023119 -0.0139379
+ 1.921e+11Hz -0.023136 -0.0139196
+ 1.922e+11Hz -0.0231528 -0.0139013
+ 1.923e+11Hz -0.0231695 -0.0138828
+ 1.924e+11Hz -0.0231862 -0.0138644
+ 1.925e+11Hz -0.0232027 -0.0138458
+ 1.926e+11Hz -0.0232191 -0.0138271
+ 1.927e+11Hz -0.0232354 -0.0138084
+ 1.928e+11Hz -0.0232516 -0.0137897
+ 1.929e+11Hz -0.0232677 -0.0137708
+ 1.93e+11Hz -0.0232837 -0.0137519
+ 1.931e+11Hz -0.0232996 -0.013733
+ 1.932e+11Hz -0.0233154 -0.0137139
+ 1.933e+11Hz -0.0233311 -0.0136948
+ 1.934e+11Hz -0.0233466 -0.0136757
+ 1.935e+11Hz -0.0233621 -0.0136565
+ 1.936e+11Hz -0.0233774 -0.0136372
+ 1.937e+11Hz -0.0233926 -0.0136179
+ 1.938e+11Hz -0.0234077 -0.0135985
+ 1.939e+11Hz -0.0234227 -0.0135791
+ 1.94e+11Hz -0.0234376 -0.0135596
+ 1.941e+11Hz -0.0234523 -0.0135401
+ 1.942e+11Hz -0.023467 -0.0135206
+ 1.943e+11Hz -0.0234815 -0.0135009
+ 1.944e+11Hz -0.0234959 -0.0134813
+ 1.945e+11Hz -0.0235102 -0.0134616
+ 1.946e+11Hz -0.0235244 -0.0134419
+ 1.947e+11Hz -0.0235385 -0.0134221
+ 1.948e+11Hz -0.0235525 -0.0134023
+ 1.949e+11Hz -0.0235663 -0.0133824
+ 1.95e+11Hz -0.02358 -0.0133625
+ 1.951e+11Hz -0.0235936 -0.0133426
+ 1.952e+11Hz -0.0236071 -0.0133227
+ 1.953e+11Hz -0.0236205 -0.0133027
+ 1.954e+11Hz -0.0236337 -0.0132827
+ 1.955e+11Hz -0.0236469 -0.0132627
+ 1.956e+11Hz -0.0236599 -0.0132426
+ 1.957e+11Hz -0.0236728 -0.0132226
+ 1.958e+11Hz -0.0236856 -0.0132025
+ 1.959e+11Hz -0.0236982 -0.0131824
+ 1.96e+11Hz -0.0237108 -0.0131622
+ 1.961e+11Hz -0.0237232 -0.0131421
+ 1.962e+11Hz -0.0237355 -0.0131219
+ 1.963e+11Hz -0.0237477 -0.0131018
+ 1.964e+11Hz -0.0237598 -0.0130816
+ 1.965e+11Hz -0.0237718 -0.0130614
+ 1.966e+11Hz -0.0237836 -0.0130412
+ 1.967e+11Hz -0.0237953 -0.013021
+ 1.968e+11Hz -0.0238069 -0.0130008
+ 1.969e+11Hz -0.0238184 -0.0129806
+ 1.97e+11Hz -0.0238298 -0.0129604
+ 1.971e+11Hz -0.0238411 -0.0129402
+ 1.972e+11Hz -0.0238522 -0.01292
+ 1.973e+11Hz -0.0238633 -0.0128998
+ 1.974e+11Hz -0.0238742 -0.0128796
+ 1.975e+11Hz -0.023885 -0.0128594
+ 1.976e+11Hz -0.0238957 -0.0128392
+ 1.977e+11Hz -0.0239063 -0.012819
+ 1.978e+11Hz -0.0239168 -0.0127989
+ 1.979e+11Hz -0.0239271 -0.0127787
+ 1.98e+11Hz -0.0239374 -0.0127586
+ 1.981e+11Hz -0.0239475 -0.0127385
+ 1.982e+11Hz -0.0239575 -0.0127184
+ 1.983e+11Hz -0.0239675 -0.0126984
+ 1.984e+11Hz -0.0239773 -0.0126783
+ 1.985e+11Hz -0.023987 -0.0126583
+ 1.986e+11Hz -0.0239966 -0.0126383
+ 1.987e+11Hz -0.0240061 -0.0126183
+ 1.988e+11Hz -0.0240155 -0.0125984
+ 1.989e+11Hz -0.0240247 -0.0125785
+ 1.99e+11Hz -0.0240339 -0.0125586
+ 1.991e+11Hz -0.024043 -0.0125388
+ 1.992e+11Hz -0.024052 -0.012519
+ 1.993e+11Hz -0.0240608 -0.0124992
+ 1.994e+11Hz -0.0240696 -0.0124795
+ 1.995e+11Hz -0.0240783 -0.0124598
+ 1.996e+11Hz -0.0240869 -0.0124401
+ 1.997e+11Hz -0.0240954 -0.0124205
+ 1.998e+11Hz -0.0241037 -0.0124009
+ 1.999e+11Hz -0.024112 -0.0123814
+ 2e+11Hz -0.0241202 -0.0123619
+ 2.001e+11Hz -0.0241283 -0.0123425
+ 2.002e+11Hz -0.0241364 -0.0123231
+ 2.003e+11Hz -0.0241443 -0.0123038
+ 2.004e+11Hz -0.0241521 -0.0122845
+ 2.005e+11Hz -0.0241599 -0.0122653
+ 2.006e+11Hz -0.0241675 -0.0122461
+ 2.007e+11Hz -0.0241751 -0.012227
+ 2.008e+11Hz -0.0241826 -0.0122079
+ 2.009e+11Hz -0.02419 -0.0121889
+ 2.01e+11Hz -0.0241974 -0.01217
+ 2.011e+11Hz -0.0242046 -0.0121511
+ 2.012e+11Hz -0.0242118 -0.0121323
+ 2.013e+11Hz -0.0242189 -0.0121136
+ 2.014e+11Hz -0.024226 -0.0120949
+ 2.015e+11Hz -0.0242329 -0.0120762
+ 2.016e+11Hz -0.0242398 -0.0120577
+ 2.017e+11Hz -0.0242466 -0.0120392
+ 2.018e+11Hz -0.0242534 -0.0120208
+ 2.019e+11Hz -0.0242601 -0.0120024
+ 2.02e+11Hz -0.0242667 -0.0119841
+ 2.021e+11Hz -0.0242732 -0.0119659
+ 2.022e+11Hz -0.0242797 -0.0119478
+ 2.023e+11Hz -0.0242861 -0.0119297
+ 2.024e+11Hz -0.0242925 -0.0119118
+ 2.025e+11Hz -0.0242988 -0.0118938
+ 2.026e+11Hz -0.0243051 -0.011876
+ 2.027e+11Hz -0.0243113 -0.0118582
+ 2.028e+11Hz -0.0243175 -0.0118406
+ 2.029e+11Hz -0.0243236 -0.011823
+ 2.03e+11Hz -0.0243296 -0.0118054
+ 2.031e+11Hz -0.0243357 -0.011788
+ 2.032e+11Hz -0.0243416 -0.0117706
+ 2.033e+11Hz -0.0243476 -0.0117533
+ 2.034e+11Hz -0.0243535 -0.0117361
+ 2.035e+11Hz -0.0243593 -0.011719
+ 2.036e+11Hz -0.0243651 -0.011702
+ 2.037e+11Hz -0.0243709 -0.011685
+ 2.038e+11Hz -0.0243767 -0.0116682
+ 2.039e+11Hz -0.0243824 -0.0116514
+ 2.04e+11Hz -0.0243881 -0.0116347
+ 2.041e+11Hz -0.0243938 -0.0116181
+ 2.042e+11Hz -0.0243994 -0.0116016
+ 2.043e+11Hz -0.024405 -0.0115851
+ 2.044e+11Hz -0.0244106 -0.0115688
+ 2.045e+11Hz -0.0244162 -0.0115525
+ 2.046e+11Hz -0.0244218 -0.0115363
+ 2.047e+11Hz -0.0244273 -0.0115202
+ 2.048e+11Hz -0.0244329 -0.0115042
+ 2.049e+11Hz -0.0244384 -0.0114883
+ 2.05e+11Hz -0.0244439 -0.0114724
+ 2.051e+11Hz -0.0244495 -0.0114567
+ 2.052e+11Hz -0.024455 -0.011441
+ 2.053e+11Hz -0.0244605 -0.0114254
+ 2.054e+11Hz -0.024466 -0.0114099
+ 2.055e+11Hz -0.0244715 -0.0113945
+ 2.056e+11Hz -0.0244771 -0.0113792
+ 2.057e+11Hz -0.0244826 -0.011364
+ 2.058e+11Hz -0.0244881 -0.0113489
+ 2.059e+11Hz -0.0244937 -0.0113338
+ 2.06e+11Hz -0.0244993 -0.0113188
+ 2.061e+11Hz -0.0245049 -0.0113039
+ 2.062e+11Hz -0.0245105 -0.0112891
+ 2.063e+11Hz -0.0245161 -0.0112744
+ 2.064e+11Hz -0.0245217 -0.0112598
+ 2.065e+11Hz -0.0245274 -0.0112452
+ 2.066e+11Hz -0.0245331 -0.0112307
+ 2.067e+11Hz -0.0245389 -0.0112163
+ 2.068e+11Hz -0.0245446 -0.011202
+ 2.069e+11Hz -0.0245504 -0.0111878
+ 2.07e+11Hz -0.0245563 -0.0111737
+ 2.071e+11Hz -0.0245621 -0.0111596
+ 2.072e+11Hz -0.024568 -0.0111456
+ 2.073e+11Hz -0.024574 -0.0111317
+ 2.074e+11Hz -0.02458 -0.0111178
+ 2.075e+11Hz -0.0245861 -0.0111041
+ 2.076e+11Hz -0.0245921 -0.0110904
+ 2.077e+11Hz -0.0245983 -0.0110768
+ 2.078e+11Hz -0.0246045 -0.0110632
+ 2.079e+11Hz -0.0246107 -0.0110497
+ 2.08e+11Hz -0.0246171 -0.0110363
+ 2.081e+11Hz -0.0246234 -0.011023
+ 2.082e+11Hz -0.0246299 -0.0110097
+ 2.083e+11Hz -0.0246364 -0.0109965
+ 2.084e+11Hz -0.0246429 -0.0109834
+ 2.085e+11Hz -0.0246496 -0.0109703
+ 2.086e+11Hz -0.0246563 -0.0109573
+ 2.087e+11Hz -0.024663 -0.0109444
+ 2.088e+11Hz -0.0246699 -0.0109315
+ 2.089e+11Hz -0.0246768 -0.0109186
+ 2.09e+11Hz -0.0246838 -0.0109058
+ 2.091e+11Hz -0.0246909 -0.0108931
+ 2.092e+11Hz -0.024698 -0.0108804
+ 2.093e+11Hz -0.0247053 -0.0108678
+ 2.094e+11Hz -0.0247126 -0.0108553
+ 2.095e+11Hz -0.02472 -0.0108427
+ 2.096e+11Hz -0.0247275 -0.0108302
+ 2.097e+11Hz -0.0247351 -0.0108178
+ 2.098e+11Hz -0.0247428 -0.0108054
+ 2.099e+11Hz -0.0247505 -0.0107931
+ 2.1e+11Hz -0.0247584 -0.0107807
+ 2.101e+11Hz -0.0247664 -0.0107685
+ 2.102e+11Hz -0.0247744 -0.0107562
+ 2.103e+11Hz -0.0247826 -0.010744
+ 2.104e+11Hz -0.0247909 -0.0107318
+ 2.105e+11Hz -0.0247992 -0.0107197
+ 2.106e+11Hz -0.0248077 -0.0107075
+ 2.107e+11Hz -0.0248163 -0.0106954
+ 2.108e+11Hz -0.024825 -0.0106833
+ 2.109e+11Hz -0.0248338 -0.0106712
+ 2.11e+11Hz -0.0248427 -0.0106592
+ 2.111e+11Hz -0.0248517 -0.0106472
+ 2.112e+11Hz -0.0248608 -0.0106351
+ 2.113e+11Hz -0.02487 -0.0106231
+ 2.114e+11Hz -0.0248794 -0.0106111
+ 2.115e+11Hz -0.0248889 -0.0105991
+ 2.116e+11Hz -0.0248985 -0.0105871
+ 2.117e+11Hz -0.0249082 -0.0105751
+ 2.118e+11Hz -0.024918 -0.010563
+ 2.119e+11Hz -0.024928 -0.010551
+ 2.12e+11Hz -0.024938 -0.010539
+ 2.121e+11Hz -0.0249482 -0.0105269
+ 2.122e+11Hz -0.0249586 -0.0105149
+ 2.123e+11Hz -0.024969 -0.0105028
+ 2.124e+11Hz -0.0249796 -0.0104907
+ 2.125e+11Hz -0.0249903 -0.0104786
+ 2.126e+11Hz -0.0250011 -0.0104665
+ 2.127e+11Hz -0.025012 -0.0104543
+ 2.128e+11Hz -0.0250231 -0.0104421
+ 2.129e+11Hz -0.0250343 -0.0104299
+ 2.13e+11Hz -0.0250456 -0.0104176
+ 2.131e+11Hz -0.0250571 -0.0104053
+ 2.132e+11Hz -0.0250687 -0.0103929
+ 2.133e+11Hz -0.0250804 -0.0103805
+ 2.134e+11Hz -0.0250923 -0.0103681
+ 2.135e+11Hz -0.0251043 -0.0103556
+ 2.136e+11Hz -0.0251164 -0.010343
+ 2.137e+11Hz -0.0251286 -0.0103304
+ 2.138e+11Hz -0.025141 -0.0103177
+ 2.139e+11Hz -0.0251535 -0.010305
+ 2.14e+11Hz -0.0251661 -0.0102922
+ 2.141e+11Hz -0.0251789 -0.0102793
+ 2.142e+11Hz -0.0251918 -0.0102663
+ 2.143e+11Hz -0.0252048 -0.0102533
+ 2.144e+11Hz -0.025218 -0.0102402
+ 2.145e+11Hz -0.0252313 -0.010227
+ 2.146e+11Hz -0.0252447 -0.0102137
+ 2.147e+11Hz -0.0252583 -0.0102004
+ 2.148e+11Hz -0.0252719 -0.0101869
+ 2.149e+11Hz -0.0252857 -0.0101733
+ 2.15e+11Hz -0.0252997 -0.0101597
+ 2.151e+11Hz -0.0253137 -0.0101459
+ 2.152e+11Hz -0.0253279 -0.0101321
+ 2.153e+11Hz -0.0253422 -0.0101181
+ 2.154e+11Hz -0.0253567 -0.010104
+ 2.155e+11Hz -0.0253713 -0.0100898
+ 2.156e+11Hz -0.0253859 -0.0100755
+ 2.157e+11Hz -0.0254008 -0.0100611
+ 2.158e+11Hz -0.0254157 -0.0100466
+ 2.159e+11Hz -0.0254307 -0.0100319
+ 2.16e+11Hz -0.0254459 -0.0100171
+ 2.161e+11Hz -0.0254612 -0.0100021
+ 2.162e+11Hz -0.0254766 -0.00998704
+ 2.163e+11Hz -0.0254921 -0.00997182
+ 2.164e+11Hz -0.0255078 -0.00995646
+ 2.165e+11Hz -0.0255235 -0.00994096
+ 2.166e+11Hz -0.0255394 -0.0099253
+ 2.167e+11Hz -0.0255553 -0.00990949
+ 2.168e+11Hz -0.0255714 -0.00989353
+ 2.169e+11Hz -0.0255876 -0.00987741
+ 2.17e+11Hz -0.0256039 -0.00986113
+ 2.171e+11Hz -0.0256203 -0.00984469
+ 2.172e+11Hz -0.0256368 -0.00982807
+ 2.173e+11Hz -0.0256533 -0.00981129
+ 2.174e+11Hz -0.02567 -0.00979434
+ 2.175e+11Hz -0.0256868 -0.00977721
+ 2.176e+11Hz -0.0257037 -0.0097599
+ 2.177e+11Hz -0.0257206 -0.00974241
+ 2.178e+11Hz -0.0257377 -0.00972474
+ 2.179e+11Hz -0.0257548 -0.00970688
+ 2.18e+11Hz -0.025772 -0.00968883
+ 2.181e+11Hz -0.0257893 -0.00967059
+ 2.182e+11Hz -0.0258067 -0.00965215
+ 2.183e+11Hz -0.0258242 -0.00963351
+ 2.184e+11Hz -0.0258417 -0.00961468
+ 2.185e+11Hz -0.0258593 -0.00959564
+ 2.186e+11Hz -0.025877 -0.00957639
+ 2.187e+11Hz -0.0258947 -0.00955694
+ 2.188e+11Hz -0.0259125 -0.00953728
+ 2.189e+11Hz -0.0259304 -0.0095174
+ 2.19e+11Hz -0.0259483 -0.00949731
+ 2.191e+11Hz -0.0259663 -0.00947699
+ 2.192e+11Hz -0.0259843 -0.00945646
+ 2.193e+11Hz -0.0260024 -0.00943571
+ 2.194e+11Hz -0.0260205 -0.00941473
+ 2.195e+11Hz -0.0260386 -0.00939352
+ 2.196e+11Hz -0.0260568 -0.00937209
+ 2.197e+11Hz -0.0260751 -0.00935042
+ 2.198e+11Hz -0.0260933 -0.00932852
+ 2.199e+11Hz -0.0261116 -0.00930638
+ 2.2e+11Hz -0.02613 -0.00928401
+ 2.201e+11Hz -0.0261483 -0.00926139
+ 2.202e+11Hz -0.0261667 -0.00923854
+ 2.203e+11Hz -0.0261851 -0.00921544
+ 2.204e+11Hz -0.0262035 -0.00919209
+ 2.205e+11Hz -0.0262219 -0.0091685
+ 2.206e+11Hz -0.0262403 -0.00914466
+ 2.207e+11Hz -0.0262587 -0.00912057
+ 2.208e+11Hz -0.0262771 -0.00909623
+ 2.209e+11Hz -0.0262955 -0.00907164
+ 2.21e+11Hz -0.0263139 -0.00904679
+ 2.211e+11Hz -0.0263323 -0.00902169
+ 2.212e+11Hz -0.0263506 -0.00899633
+ 2.213e+11Hz -0.026369 -0.00897071
+ 2.214e+11Hz -0.0263873 -0.00894483
+ 2.215e+11Hz -0.0264056 -0.00891869
+ 2.216e+11Hz -0.0264238 -0.00889229
+ 2.217e+11Hz -0.026442 -0.00886562
+ 2.218e+11Hz -0.0264602 -0.00883869
+ 2.219e+11Hz -0.0264783 -0.0088115
+ 2.22e+11Hz -0.0264964 -0.00878404
+ 2.221e+11Hz -0.0265144 -0.00875631
+ 2.222e+11Hz -0.0265324 -0.00872832
+ 2.223e+11Hz -0.0265503 -0.00870006
+ 2.224e+11Hz -0.0265682 -0.00867153
+ 2.225e+11Hz -0.0265859 -0.00864274
+ 2.226e+11Hz -0.0266036 -0.00861367
+ 2.227e+11Hz -0.0266213 -0.00858434
+ 2.228e+11Hz -0.0266388 -0.00855473
+ 2.229e+11Hz -0.0266563 -0.00852486
+ 2.23e+11Hz -0.0266736 -0.00849471
+ 2.231e+11Hz -0.0266909 -0.0084643
+ 2.232e+11Hz -0.0267081 -0.00843362
+ 2.233e+11Hz -0.0267251 -0.00840266
+ 2.234e+11Hz -0.0267421 -0.00837144
+ 2.235e+11Hz -0.0267589 -0.00833994
+ 2.236e+11Hz -0.0267757 -0.00830818
+ 2.237e+11Hz -0.0267923 -0.00827615
+ 2.238e+11Hz -0.0268087 -0.00824385
+ 2.239e+11Hz -0.0268251 -0.00821128
+ 2.24e+11Hz -0.0268413 -0.00817845
+ 2.241e+11Hz -0.0268574 -0.00814535
+ 2.242e+11Hz -0.0268733 -0.00811198
+ 2.243e+11Hz -0.0268891 -0.00807835
+ 2.244e+11Hz -0.0269047 -0.00804445
+ 2.245e+11Hz -0.0269202 -0.00801029
+ 2.246e+11Hz -0.0269355 -0.00797587
+ 2.247e+11Hz -0.0269507 -0.00794119
+ 2.248e+11Hz -0.0269657 -0.00790625
+ 2.249e+11Hz -0.0269805 -0.00787105
+ 2.25e+11Hz -0.0269951 -0.00783559
+ 2.251e+11Hz -0.0270096 -0.00779987
+ 2.252e+11Hz -0.0270238 -0.00776391
+ 2.253e+11Hz -0.0270379 -0.00772769
+ 2.254e+11Hz -0.0270518 -0.00769121
+ 2.255e+11Hz -0.0270655 -0.00765449
+ 2.256e+11Hz -0.027079 -0.00761752
+ 2.257e+11Hz -0.0270922 -0.00758031
+ 2.258e+11Hz -0.0271053 -0.00754285
+ 2.259e+11Hz -0.0271182 -0.00750515
+ 2.26e+11Hz -0.0271308 -0.00746721
+ 2.261e+11Hz -0.0271432 -0.00742904
+ 2.262e+11Hz -0.0271554 -0.00739062
+ 2.263e+11Hz -0.0271673 -0.00735198
+ 2.264e+11Hz -0.027179 -0.0073131
+ 2.265e+11Hz -0.0271905 -0.007274
+ 2.266e+11Hz -0.0272017 -0.00723467
+ 2.267e+11Hz -0.0272127 -0.00719512
+ 2.268e+11Hz -0.0272234 -0.00715534
+ 2.269e+11Hz -0.0272339 -0.00711535
+ 2.27e+11Hz -0.0272441 -0.00707515
+ 2.271e+11Hz -0.027254 -0.00703473
+ 2.272e+11Hz -0.0272637 -0.0069941
+ 2.273e+11Hz -0.0272731 -0.00695327
+ 2.274e+11Hz -0.0272823 -0.00691223
+ 2.275e+11Hz -0.0272911 -0.00687099
+ 2.276e+11Hz -0.0272997 -0.00682956
+ 2.277e+11Hz -0.027308 -0.00678793
+ 2.278e+11Hz -0.027316 -0.00674611
+ 2.279e+11Hz -0.0273237 -0.00670411
+ 2.28e+11Hz -0.0273311 -0.00666192
+ 2.281e+11Hz -0.0273383 -0.00661955
+ 2.282e+11Hz -0.0273451 -0.00657701
+ 2.283e+11Hz -0.0273516 -0.00653429
+ 2.284e+11Hz -0.0273578 -0.0064914
+ 2.285e+11Hz -0.0273637 -0.00644835
+ 2.286e+11Hz -0.0273693 -0.00640514
+ 2.287e+11Hz -0.0273746 -0.00636176
+ 2.288e+11Hz -0.0273795 -0.00631824
+ 2.289e+11Hz -0.0273841 -0.00627456
+ 2.29e+11Hz -0.0273884 -0.00623074
+ 2.291e+11Hz -0.0273924 -0.00618678
+ 2.292e+11Hz -0.0273961 -0.00614267
+ 2.293e+11Hz -0.0273994 -0.00609844
+ 2.294e+11Hz -0.0274024 -0.00605407
+ 2.295e+11Hz -0.027405 -0.00600958
+ 2.296e+11Hz -0.0274073 -0.00596497
+ 2.297e+11Hz -0.0274092 -0.00592024
+ 2.298e+11Hz -0.0274109 -0.0058754
+ 2.299e+11Hz -0.0274121 -0.00583045
+ 2.3e+11Hz -0.027413 -0.00578539
+ 2.301e+11Hz -0.0274136 -0.00574024
+ 2.302e+11Hz -0.0274138 -0.00569499
+ 2.303e+11Hz -0.0274137 -0.00564965
+ 2.304e+11Hz -0.0274131 -0.00560423
+ 2.305e+11Hz -0.0274123 -0.00555873
+ 2.306e+11Hz -0.0274111 -0.00551315
+ 2.307e+11Hz -0.0274095 -0.0054675
+ 2.308e+11Hz -0.0274075 -0.00542178
+ 2.309e+11Hz -0.0274052 -0.005376
+ 2.31e+11Hz -0.0274025 -0.00533016
+ 2.311e+11Hz -0.0273995 -0.00528427
+ 2.312e+11Hz -0.0273961 -0.00523833
+ 2.313e+11Hz -0.0273923 -0.00519235
+ 2.314e+11Hz -0.0273881 -0.00514633
+ 2.315e+11Hz -0.0273836 -0.00510028
+ 2.316e+11Hz -0.0273787 -0.0050542
+ 2.317e+11Hz -0.0273734 -0.0050081
+ 2.318e+11Hz -0.0273678 -0.00496198
+ 2.319e+11Hz -0.0273617 -0.00491584
+ 2.32e+11Hz -0.0273553 -0.0048697
+ 2.321e+11Hz -0.0273485 -0.00482355
+ 2.322e+11Hz -0.0273414 -0.00477741
+ 2.323e+11Hz -0.0273339 -0.00473127
+ 2.324e+11Hz -0.0273259 -0.00468514
+ 2.325e+11Hz -0.0273177 -0.00463904
+ 2.326e+11Hz -0.027309 -0.00459295
+ 2.327e+11Hz -0.0272999 -0.00454689
+ 2.328e+11Hz -0.0272905 -0.00450086
+ 2.329e+11Hz -0.0272807 -0.00445486
+ 2.33e+11Hz -0.0272705 -0.00440891
+ 2.331e+11Hz -0.02726 -0.00436301
+ 2.332e+11Hz -0.027249 -0.00431716
+ 2.333e+11Hz -0.0272377 -0.00427136
+ 2.334e+11Hz -0.0272261 -0.00422563
+ 2.335e+11Hz -0.027214 -0.00417996
+ 2.336e+11Hz -0.0272016 -0.00413437
+ 2.337e+11Hz -0.0271888 -0.00408885
+ 2.338e+11Hz -0.0271756 -0.00404342
+ 2.339e+11Hz -0.027162 -0.00399807
+ 2.34e+11Hz -0.0271481 -0.00395281
+ 2.341e+11Hz -0.0271338 -0.00390765
+ 2.342e+11Hz -0.0271191 -0.00386259
+ 2.343e+11Hz -0.0271041 -0.00381764
+ 2.344e+11Hz -0.0270887 -0.00377279
+ 2.345e+11Hz -0.027073 -0.00372807
+ 2.346e+11Hz -0.0270568 -0.00368346
+ 2.347e+11Hz -0.0270404 -0.00363898
+ 2.348e+11Hz -0.0270235 -0.00359464
+ 2.349e+11Hz -0.0270063 -0.00355042
+ 2.35e+11Hz -0.0269888 -0.00350635
+ 2.351e+11Hz -0.0269709 -0.00346242
+ 2.352e+11Hz -0.0269526 -0.00341864
+ 2.353e+11Hz -0.026934 -0.00337501
+ 2.354e+11Hz -0.026915 -0.00333154
+ 2.355e+11Hz -0.0268957 -0.00328823
+ 2.356e+11Hz -0.0268761 -0.00324509
+ 2.357e+11Hz -0.0268561 -0.00320213
+ 2.358e+11Hz -0.0268357 -0.00315934
+ 2.359e+11Hz -0.0268151 -0.00311673
+ 2.36e+11Hz -0.0267941 -0.0030743
+ 2.361e+11Hz -0.0267727 -0.00303206
+ 2.362e+11Hz -0.0267511 -0.00299002
+ 2.363e+11Hz -0.0267291 -0.00294817
+ 2.364e+11Hz -0.0267068 -0.00290653
+ 2.365e+11Hz -0.0266842 -0.00286509
+ 2.366e+11Hz -0.0266612 -0.00282386
+ 2.367e+11Hz -0.026638 -0.00278284
+ 2.368e+11Hz -0.0266144 -0.00274204
+ 2.369e+11Hz -0.0265905 -0.00270146
+ 2.37e+11Hz -0.0265663 -0.00266111
+ 2.371e+11Hz -0.0265418 -0.00262099
+ 2.372e+11Hz -0.026517 -0.0025811
+ 2.373e+11Hz -0.026492 -0.00254144
+ 2.374e+11Hz -0.0264666 -0.00250203
+ 2.375e+11Hz -0.0264409 -0.00246286
+ 2.376e+11Hz -0.026415 -0.00242394
+ 2.377e+11Hz -0.0263888 -0.00238526
+ 2.378e+11Hz -0.0263623 -0.00234684
+ 2.379e+11Hz -0.0263355 -0.00230868
+ 2.38e+11Hz -0.0263084 -0.00227078
+ 2.381e+11Hz -0.0262811 -0.00223314
+ 2.382e+11Hz -0.0262535 -0.00219577
+ 2.383e+11Hz -0.0262257 -0.00215867
+ 2.384e+11Hz -0.0261976 -0.00212184
+ 2.385e+11Hz -0.0261693 -0.00208528
+ 2.386e+11Hz -0.0261407 -0.00204901
+ 2.387e+11Hz -0.0261119 -0.00201301
+ 2.388e+11Hz -0.0260828 -0.0019773
+ 2.389e+11Hz -0.0260535 -0.00194187
+ 2.39e+11Hz -0.0260239 -0.00190674
+ 2.391e+11Hz -0.0259942 -0.00187189
+ 2.392e+11Hz -0.0259642 -0.00183734
+ 2.393e+11Hz -0.025934 -0.00180309
+ 2.394e+11Hz -0.0259036 -0.00176913
+ 2.395e+11Hz -0.0258729 -0.00173548
+ 2.396e+11Hz -0.0258421 -0.00170213
+ 2.397e+11Hz -0.0258111 -0.00166908
+ 2.398e+11Hz -0.0257798 -0.00163634
+ 2.399e+11Hz -0.0257484 -0.0016039
+ 2.4e+11Hz -0.0257168 -0.00157178
+ 2.401e+11Hz -0.025685 -0.00153997
+ 2.402e+11Hz -0.025653 -0.00150848
+ 2.403e+11Hz -0.0256209 -0.0014773
+ 2.404e+11Hz -0.0255886 -0.00144644
+ 2.405e+11Hz -0.0255561 -0.00141589
+ 2.406e+11Hz -0.0255234 -0.00138567
+ 2.407e+11Hz -0.0254906 -0.00135577
+ 2.408e+11Hz -0.0254577 -0.00132619
+ 2.409e+11Hz -0.0254246 -0.00129693
+ 2.41e+11Hz -0.0253913 -0.001268
+ 2.411e+11Hz -0.0253579 -0.0012394
+ 2.412e+11Hz -0.0253244 -0.00121112
+ 2.413e+11Hz -0.0252908 -0.00118317
+ 2.414e+11Hz -0.025257 -0.00115555
+ 2.415e+11Hz -0.0252231 -0.00112826
+ 2.416e+11Hz -0.0251891 -0.00110129
+ 2.417e+11Hz -0.025155 -0.00107466
+ 2.418e+11Hz -0.0251207 -0.00104836
+ 2.419e+11Hz -0.0250864 -0.00102239
+ 2.42e+11Hz -0.025052 -0.000996754
+ 2.421e+11Hz -0.0250174 -0.000971449
+ 2.422e+11Hz -0.0249828 -0.000946475
+ 2.423e+11Hz -0.0249481 -0.000921835
+ 2.424e+11Hz -0.0249134 -0.000897527
+ 2.425e+11Hz -0.0248785 -0.000873551
+ 2.426e+11Hz -0.0248436 -0.000849908
+ 2.427e+11Hz -0.0248086 -0.000826598
+ 2.428e+11Hz -0.0247735 -0.000803619
+ 2.429e+11Hz -0.0247384 -0.000780973
+ 2.43e+11Hz -0.0247033 -0.000758658
+ 2.431e+11Hz -0.0246681 -0.000736674
+ 2.432e+11Hz -0.0246328 -0.000715021
+ 2.433e+11Hz -0.0245975 -0.000693698
+ 2.434e+11Hz -0.0245622 -0.000672704
+ 2.435e+11Hz -0.0245268 -0.000652039
+ 2.436e+11Hz -0.0244914 -0.000631703
+ 2.437e+11Hz -0.024456 -0.000611694
+ 2.438e+11Hz -0.0244206 -0.000592011
+ 2.439e+11Hz -0.0243851 -0.000572654
+ 2.44e+11Hz -0.0243497 -0.000553621
+ 2.441e+11Hz -0.0243142 -0.000534912
+ 2.442e+11Hz -0.0242788 -0.000516525
+ 2.443e+11Hz -0.0242433 -0.000498459
+ 2.444e+11Hz -0.0242078 -0.000480714
+ 2.445e+11Hz -0.0241724 -0.000463287
+ 2.446e+11Hz -0.024137 -0.000446178
+ 2.447e+11Hz -0.0241015 -0.000429384
+ 2.448e+11Hz -0.0240662 -0.000412905
+ 2.449e+11Hz -0.0240308 -0.00039674
+ 2.45e+11Hz -0.0239955 -0.000380885
+ 2.451e+11Hz -0.0239601 -0.000365341
+ 2.452e+11Hz -0.0239249 -0.000350105
+ 2.453e+11Hz -0.0238897 -0.000335176
+ 2.454e+11Hz -0.0238545 -0.000320551
+ 2.455e+11Hz -0.0238193 -0.000306229
+ 2.456e+11Hz -0.0237843 -0.000292209
+ 2.457e+11Hz -0.0237492 -0.000278487
+ 2.458e+11Hz -0.0237143 -0.000265063
+ 2.459e+11Hz -0.0236794 -0.000251935
+ 2.46e+11Hz -0.0236445 -0.000239099
+ 2.461e+11Hz -0.0236097 -0.000226555
+ 2.462e+11Hz -0.023575 -0.0002143
+ 2.463e+11Hz -0.0235404 -0.000202332
+ 2.464e+11Hz -0.0235059 -0.000190649
+ 2.465e+11Hz -0.0234714 -0.000179248
+ 2.466e+11Hz -0.023437 -0.000168128
+ 2.467e+11Hz -0.0234027 -0.000157285
+ 2.468e+11Hz -0.0233685 -0.000146718
+ 2.469e+11Hz -0.0233344 -0.000136425
+ 2.47e+11Hz -0.0233004 -0.000126402
+ 2.471e+11Hz -0.0232665 -0.000116648
+ 2.472e+11Hz -0.0232327 -0.00010716
+ 2.473e+11Hz -0.023199 -9.7935e-05
+ 2.474e+11Hz -0.0231654 -8.89712e-05
+ 2.475e+11Hz -0.023132 -8.02658e-05
+ 2.476e+11Hz -0.0230986 -7.18163e-05
+ 2.477e+11Hz -0.0230653 -6.36199e-05
+ 2.478e+11Hz -0.0230322 -5.56742e-05
+ 2.479e+11Hz -0.0229992 -4.79764e-05
+ 2.48e+11Hz -0.0229663 -4.05238e-05
+ 2.481e+11Hz -0.0229336 -3.33139e-05
+ 2.482e+11Hz -0.0229009 -2.63438e-05
+ 2.483e+11Hz -0.0228684 -1.96108e-05
+ 2.484e+11Hz -0.0228361 -1.31123e-05
+ 2.485e+11Hz -0.0228038 -6.84528e-06
+ 2.486e+11Hz -0.0227717 -8.0713e-07
+ 2.487e+11Hz -0.0227398 5.005e-06
+ 2.488e+11Hz -0.022708 1.05939e-05
+ 2.489e+11Hz -0.0226763 1.59625e-05
+ 2.49e+11Hz -0.0226448 2.11135e-05
+ 2.491e+11Hz -0.0226134 2.60498e-05
+ 2.492e+11Hz -0.0225822 3.07743e-05
+ 2.493e+11Hz -0.0225511 3.52899e-05
+ 2.494e+11Hz -0.0225202 3.95994e-05
+ 2.495e+11Hz -0.0224894 4.37058e-05
+ 2.496e+11Hz -0.0224588 4.76118e-05
+ 2.497e+11Hz -0.0224284 5.13205e-05
+ 2.498e+11Hz -0.0223981 5.48347e-05
+ 2.499e+11Hz -0.0223679 5.81574e-05
+ 2.5e+11Hz -0.022338 6.12915e-05
+ 2.501e+11Hz -0.0223082 6.42398e-05
+ 2.502e+11Hz -0.0222785 6.70053e-05
+ 2.503e+11Hz -0.022249 6.9591e-05
+ 2.504e+11Hz -0.0222197 7.19997e-05
+ 2.505e+11Hz -0.0221906 7.42343e-05
+ 2.506e+11Hz -0.0221616 7.62979e-05
+ 2.507e+11Hz -0.0221328 7.81932e-05
+ 2.508e+11Hz -0.0221042 7.99233e-05
+ 2.509e+11Hz -0.0220758 8.1491e-05
+ 2.51e+11Hz -0.0220475 8.28993e-05
+ 2.511e+11Hz -0.0220194 8.4151e-05
+ 2.512e+11Hz -0.0219915 8.52491e-05
+ 2.513e+11Hz -0.0219637 8.61964e-05
+ 2.514e+11Hz -0.0219362 8.69958e-05
+ 2.515e+11Hz -0.0219088 8.76503e-05
+ 2.516e+11Hz -0.0218816 8.81626e-05
+ 2.517e+11Hz -0.0218545 8.85356e-05
+ 2.518e+11Hz -0.0218277 8.87723e-05
+ 2.519e+11Hz -0.021801 8.88754e-05
+ 2.52e+11Hz -0.0217745 8.88478e-05
+ 2.521e+11Hz -0.0217482 8.86923e-05
+ 2.522e+11Hz -0.0217221 8.84117e-05
+ 2.523e+11Hz -0.0216962 8.80088e-05
+ 2.524e+11Hz -0.0216704 8.74864e-05
+ 2.525e+11Hz -0.0216449 8.68474e-05
+ 2.526e+11Hz -0.0216195 8.60944e-05
+ 2.527e+11Hz -0.0215943 8.52302e-05
+ 2.528e+11Hz -0.0215693 8.42576e-05
+ 2.529e+11Hz -0.0215445 8.31793e-05
+ 2.53e+11Hz -0.0215198 8.1998e-05
+ 2.531e+11Hz -0.0214954 8.07164e-05
+ 2.532e+11Hz -0.0214711 7.93372e-05
+ 2.533e+11Hz -0.0214471 7.78631e-05
+ 2.534e+11Hz -0.0214232 7.62967e-05
+ 2.535e+11Hz -0.0213995 7.46407e-05
+ 2.536e+11Hz -0.021376 7.28978e-05
+ 2.537e+11Hz -0.0213526 7.10704e-05
+ 2.538e+11Hz -0.0213295 6.91612e-05
+ 2.539e+11Hz -0.0213066 6.71729e-05
+ 2.54e+11Hz -0.0212838 6.5108e-05
+ 2.541e+11Hz -0.0212612 6.29689e-05
+ 2.542e+11Hz -0.0212389 6.07584e-05
+ 2.543e+11Hz -0.0212167 5.84788e-05
+ 2.544e+11Hz -0.0211947 5.61327e-05
+ 2.545e+11Hz -0.0211728 5.37226e-05
+ 2.546e+11Hz -0.0211512 5.1251e-05
+ 2.547e+11Hz -0.0211298 4.87203e-05
+ 2.548e+11Hz -0.0211085 4.61329e-05
+ 2.549e+11Hz -0.0210874 4.34914e-05
+ 2.55e+11Hz -0.0210665 4.0798e-05
+ 2.551e+11Hz -0.0210458 3.80552e-05
+ 2.552e+11Hz -0.0210253 3.52655e-05
+ 2.553e+11Hz -0.021005 3.2431e-05
+ 2.554e+11Hz -0.0209849 2.95543e-05
+ 2.555e+11Hz -0.0209649 2.66376e-05
+ 2.556e+11Hz -0.0209451 2.36832e-05
+ 2.557e+11Hz -0.0209255 2.06935e-05
+ 2.558e+11Hz -0.0209061 1.76707e-05
+ 2.559e+11Hz -0.0208869 1.46172e-05
+ 2.56e+11Hz -0.0208679 1.15352e-05
+ 2.561e+11Hz -0.020849 8.42689e-06
+ 2.562e+11Hz -0.0208303 5.29458e-06
+ 2.563e+11Hz -0.0208119 2.14047e-06
+ 2.564e+11Hz -0.0207935 -1.03323e-06
+ 2.565e+11Hz -0.0207754 -4.22433e-06
+ 2.566e+11Hz -0.0207575 -7.43064e-06
+ 2.567e+11Hz -0.0207397 -1.065e-05
+ 2.568e+11Hz -0.0207221 -1.38802e-05
+ 2.569e+11Hz -0.0207047 -1.71192e-05
+ 2.57e+11Hz -0.0206875 -2.03647e-05
+ 2.571e+11Hz -0.0206704 -2.36147e-05
+ 2.572e+11Hz -0.0206535 -2.68671e-05
+ 2.573e+11Hz -0.0206368 -3.01198e-05
+ 2.574e+11Hz -0.0206203 -3.33706e-05
+ 2.575e+11Hz -0.020604 -3.66174e-05
+ 2.576e+11Hz -0.0205878 -3.98583e-05
+ 2.577e+11Hz -0.0205718 -4.30911e-05
+ 2.578e+11Hz -0.020556 -4.63138e-05
+ 2.579e+11Hz -0.0205403 -4.95243e-05
+ 2.58e+11Hz -0.0205248 -5.27206e-05
+ 2.581e+11Hz -0.0205095 -5.59006e-05
+ 2.582e+11Hz -0.0204944 -5.90624e-05
+ 2.583e+11Hz -0.0204794 -6.22039e-05
+ 2.584e+11Hz -0.0204646 -6.53231e-05
+ 2.585e+11Hz -0.02045 -6.8418e-05
+ 2.586e+11Hz -0.0204355 -7.14866e-05
+ 2.587e+11Hz -0.0204212 -7.45269e-05
+ 2.588e+11Hz -0.0204071 -7.75369e-05
+ 2.589e+11Hz -0.0203931 -8.05147e-05
+ 2.59e+11Hz -0.0203793 -8.34582e-05
+ 2.591e+11Hz -0.0203657 -8.63655e-05
+ 2.592e+11Hz -0.0203522 -8.92346e-05
+ 2.593e+11Hz -0.0203389 -9.20635e-05
+ 2.594e+11Hz -0.0203258 -9.48504e-05
+ 2.595e+11Hz -0.0203128 -9.75931e-05
+ 2.596e+11Hz -0.0203 -0.00010029
+ 2.597e+11Hz -0.0202874 -0.000102939
+ 2.598e+11Hz -0.0202749 -0.000105537
+ 2.599e+11Hz -0.0202625 -0.000108084
+ 2.6e+11Hz -0.0202503 -0.000110577
+ 2.601e+11Hz -0.0202383 -0.000113014
+ 2.602e+11Hz -0.0202264 -0.000115394
+ 2.603e+11Hz -0.0202147 -0.000117713
+ 2.604e+11Hz -0.0202032 -0.000119971
+ 2.605e+11Hz -0.0201917 -0.000122166
+ 2.606e+11Hz -0.0201805 -0.000124295
+ 2.607e+11Hz -0.0201694 -0.000126356
+ 2.608e+11Hz -0.0201584 -0.000128348
+ 2.609e+11Hz -0.0201476 -0.000130269
+ 2.61e+11Hz -0.020137 -0.000132116
+ 2.611e+11Hz -0.0201265 -0.000133888
+ 2.612e+11Hz -0.0201161 -0.000135583
+ 2.613e+11Hz -0.0201059 -0.000137198
+ 2.614e+11Hz -0.0200958 -0.000138732
+ 2.615e+11Hz -0.0200859 -0.000140183
+ 2.616e+11Hz -0.0200761 -0.00014155
+ 2.617e+11Hz -0.0200664 -0.000142829
+ 2.618e+11Hz -0.0200569 -0.000144019
+ 2.619e+11Hz -0.0200476 -0.000145118
+ 2.62e+11Hz -0.0200383 -0.000146124
+ 2.621e+11Hz -0.0200292 -0.000147035
+ 2.622e+11Hz -0.0200203 -0.000147849
+ 2.623e+11Hz -0.0200115 -0.000148565
+ 2.624e+11Hz -0.0200028 -0.000149179
+ 2.625e+11Hz -0.0199942 -0.000149691
+ 2.626e+11Hz -0.0199858 -0.000150098
+ 2.627e+11Hz -0.0199775 -0.000150399
+ 2.628e+11Hz -0.0199693 -0.00015059
+ 2.629e+11Hz -0.0199613 -0.000150671
+ 2.63e+11Hz -0.0199534 -0.00015064
+ 2.631e+11Hz -0.0199456 -0.000150493
+ 2.632e+11Hz -0.0199379 -0.00015023
+ 2.633e+11Hz -0.0199303 -0.000149848
+ 2.634e+11Hz -0.0199229 -0.000149346
+ 2.635e+11Hz -0.0199156 -0.000148721
+ 2.636e+11Hz -0.0199084 -0.000147972
+ 2.637e+11Hz -0.0199013 -0.000147096
+ 2.638e+11Hz -0.0198943 -0.000146091
+ 2.639e+11Hz -0.0198875 -0.000144956
+ 2.64e+11Hz -0.0198807 -0.000143689
+ 2.641e+11Hz -0.0198741 -0.000142287
+ 2.642e+11Hz -0.0198676 -0.000140749
+ 2.643e+11Hz -0.0198611 -0.000139072
+ 2.644e+11Hz -0.0198548 -0.000137255
+ 2.645e+11Hz -0.0198486 -0.000135296
+ 2.646e+11Hz -0.0198425 -0.000133192
+ 2.647e+11Hz -0.0198364 -0.000130943
+ 2.648e+11Hz -0.0198305 -0.000128545
+ 2.649e+11Hz -0.0198247 -0.000125997
+ 2.65e+11Hz -0.0198189 -0.000123297
+ 2.651e+11Hz -0.0198133 -0.000120444
+ 2.652e+11Hz -0.0198077 -0.000117434
+ 2.653e+11Hz -0.0198022 -0.000114267
+ 2.654e+11Hz -0.0197968 -0.00011094
+ 2.655e+11Hz -0.0197915 -0.000107452
+ 2.656e+11Hz -0.0197863 -0.0001038
+ 2.657e+11Hz -0.0197811 -9.99837e-05
+ 2.658e+11Hz -0.019776 -9.59999e-05
+ 2.659e+11Hz -0.019771 -9.18472e-05
+ 2.66e+11Hz -0.0197661 -8.75239e-05
+ 2.661e+11Hz -0.0197612 -8.30281e-05
+ 2.662e+11Hz -0.0197564 -7.83581e-05
+ 2.663e+11Hz -0.0197517 -7.3512e-05
+ 2.664e+11Hz -0.019747 -6.84882e-05
+ 2.665e+11Hz -0.0197424 -6.32849e-05
+ 2.666e+11Hz -0.0197378 -5.79003e-05
+ 2.667e+11Hz -0.0197333 -5.23329e-05
+ 2.668e+11Hz -0.0197288 -4.65809e-05
+ 2.669e+11Hz -0.0197244 -4.06428e-05
+ 2.67e+11Hz -0.01972 -3.45167e-05
+ 2.671e+11Hz -0.0197157 -2.82013e-05
+ 2.672e+11Hz -0.0197114 -2.16949e-05
+ 2.673e+11Hz -0.0197072 -1.49959e-05
+ 2.674e+11Hz -0.0197029 -8.10288e-06
+ 2.675e+11Hz -0.0196988 -1.0143e-06
+ 2.676e+11Hz -0.0196946 6.27128e-06
+ 2.677e+11Hz -0.0196905 1.37553e-05
+ 2.678e+11Hz -0.0196863 2.14392e-05
+ 2.679e+11Hz -0.0196822 2.93242e-05
+ 2.68e+11Hz -0.0196782 3.74118e-05
+ 2.681e+11Hz -0.0196741 4.57032e-05
+ 2.682e+11Hz -0.01967 5.41997e-05
+ 2.683e+11Hz -0.019666 6.29025e-05
+ 2.684e+11Hz -0.0196619 7.18128e-05
+ 2.685e+11Hz -0.0196579 8.09317e-05
+ 2.686e+11Hz -0.0196538 9.02604e-05
+ 2.687e+11Hz -0.0196498 9.97999e-05
+ 2.688e+11Hz -0.0196457 0.000109551
+ 2.689e+11Hz -0.0196416 0.000119515
+ 2.69e+11Hz -0.0196375 0.000129693
+ 2.691e+11Hz -0.0196334 0.000140086
+ 2.692e+11Hz -0.0196292 0.000150694
+ 2.693e+11Hz -0.019625 0.000161518
+ 2.694e+11Hz -0.0196208 0.000172559
+ 2.695e+11Hz -0.0196166 0.000183818
+ 2.696e+11Hz -0.0196123 0.000195295
+ 2.697e+11Hz -0.019608 0.000206992
+ 2.698e+11Hz -0.0196036 0.000218907
+ 2.699e+11Hz -0.0195992 0.000231043
+ 2.7e+11Hz -0.0195947 0.000243399
+ 2.701e+11Hz -0.0195901 0.000255975
+ 2.702e+11Hz -0.0195855 0.000268773
+ 2.703e+11Hz -0.0195808 0.000281792
+ 2.704e+11Hz -0.0195761 0.000295032
+ 2.705e+11Hz -0.0195713 0.000308494
+ 2.706e+11Hz -0.0195664 0.000322178
+ 2.707e+11Hz -0.0195614 0.000336083
+ 2.708e+11Hz -0.0195563 0.00035021
+ 2.709e+11Hz -0.0195511 0.000364558
+ 2.71e+11Hz -0.0195459 0.000379128
+ 2.711e+11Hz -0.0195405 0.000393918
+ 2.712e+11Hz -0.0195351 0.00040893
+ 2.713e+11Hz -0.0195295 0.000424161
+ 2.714e+11Hz -0.0195238 0.000439612
+ 2.715e+11Hz -0.019518 0.000455283
+ 2.716e+11Hz -0.0195121 0.000471172
+ 2.717e+11Hz -0.019506 0.000487279
+ 2.718e+11Hz -0.0194999 0.000503603
+ 2.719e+11Hz -0.0194936 0.000520144
+ 2.72e+11Hz -0.0194871 0.000536899
+ 2.721e+11Hz -0.0194805 0.00055387
+ 2.722e+11Hz -0.0194738 0.000571054
+ 2.723e+11Hz -0.0194669 0.000588449
+ 2.724e+11Hz -0.0194599 0.000606056
+ 2.725e+11Hz -0.0194527 0.000623873
+ 2.726e+11Hz -0.0194453 0.000641898
+ 2.727e+11Hz -0.0194378 0.00066013
+ 2.728e+11Hz -0.01943 0.000678567
+ 2.729e+11Hz -0.0194222 0.000697208
+ 2.73e+11Hz -0.0194141 0.00071605
+ 2.731e+11Hz -0.0194058 0.000735093
+ 2.732e+11Hz -0.0193974 0.000754334
+ 2.733e+11Hz -0.0193888 0.000773772
+ 2.734e+11Hz -0.0193799 0.000793404
+ 2.735e+11Hz -0.0193709 0.000813228
+ 2.736e+11Hz -0.0193616 0.000833242
+ 2.737e+11Hz -0.0193522 0.000853444
+ 2.738e+11Hz -0.0193425 0.000873831
+ 2.739e+11Hz -0.0193326 0.000894401
+ 2.74e+11Hz -0.0193225 0.000915151
+ 2.741e+11Hz -0.0193121 0.000936079
+ 2.742e+11Hz -0.0193016 0.000957182
+ 2.743e+11Hz -0.0192907 0.000978457
+ 2.744e+11Hz -0.0192797 0.000999901
+ 2.745e+11Hz -0.0192684 0.00102151
+ 2.746e+11Hz -0.0192568 0.00104328
+ 2.747e+11Hz -0.019245 0.00106522
+ 2.748e+11Hz -0.0192329 0.00108731
+ 2.749e+11Hz -0.0192206 0.00110955
+ 2.75e+11Hz -0.019208 0.00113195
+ 2.751e+11Hz -0.0191951 0.00115449
+ 2.752e+11Hz -0.019182 0.00117717
+ 2.753e+11Hz -0.0191686 0.0012
+ 2.754e+11Hz -0.0191549 0.00122295
+ 2.755e+11Hz -0.0191409 0.00124604
+ 2.756e+11Hz -0.0191266 0.00126926
+ 2.757e+11Hz -0.0191121 0.00129261
+ 2.758e+11Hz -0.0190972 0.00131607
+ 2.759e+11Hz -0.0190821 0.00133965
+ 2.76e+11Hz -0.0190666 0.00136333
+ 2.761e+11Hz -0.0190509 0.00138713
+ 2.762e+11Hz -0.0190348 0.00141103
+ 2.763e+11Hz -0.0190184 0.00143503
+ 2.764e+11Hz -0.0190017 0.00145912
+ 2.765e+11Hz -0.0189847 0.0014833
+ 2.766e+11Hz -0.0189674 0.00150756
+ 2.767e+11Hz -0.0189497 0.00153191
+ 2.768e+11Hz -0.0189317 0.00155633
+ 2.769e+11Hz -0.0189134 0.00158082
+ 2.77e+11Hz -0.0188947 0.00160537
+ 2.771e+11Hz -0.0188757 0.00162998
+ 2.772e+11Hz -0.0188564 0.00165465
+ 2.773e+11Hz -0.0188367 0.00167937
+ 2.774e+11Hz -0.0188167 0.00170413
+ 2.775e+11Hz -0.0187964 0.00172893
+ 2.776e+11Hz -0.0187757 0.00175376
+ 2.777e+11Hz -0.0187546 0.00177862
+ 2.778e+11Hz -0.0187332 0.00180351
+ 2.779e+11Hz -0.0187114 0.00182841
+ 2.78e+11Hz -0.0186893 0.00185332
+ 2.781e+11Hz -0.0186668 0.00187824
+ 2.782e+11Hz -0.018644 0.00190316
+ 2.783e+11Hz -0.0186208 0.00192807
+ 2.784e+11Hz -0.0185972 0.00195297
+ 2.785e+11Hz -0.0185733 0.00197785
+ 2.786e+11Hz -0.018549 0.00200271
+ 2.787e+11Hz -0.0185243 0.00202753
+ 2.788e+11Hz -0.0184993 0.00205232
+ 2.789e+11Hz -0.0184739 0.00207707
+ 2.79e+11Hz -0.0184482 0.00210178
+ 2.791e+11Hz -0.018422 0.00212642
+ 2.792e+11Hz -0.0183955 0.00215101
+ 2.793e+11Hz -0.0183686 0.00217553
+ 2.794e+11Hz -0.0183414 0.00219998
+ 2.795e+11Hz -0.0183137 0.00222435
+ 2.796e+11Hz -0.0182857 0.00224863
+ 2.797e+11Hz -0.0182574 0.00227282
+ 2.798e+11Hz -0.0182286 0.00229692
+ 2.799e+11Hz -0.0181995 0.0023209
+ 2.8e+11Hz -0.01817 0.00234478
+ 2.801e+11Hz -0.0181401 0.00236854
+ 2.802e+11Hz -0.0181099 0.00239218
+ 2.803e+11Hz -0.0180793 0.00241568
+ 2.804e+11Hz -0.0180483 0.00243905
+ 2.805e+11Hz -0.018017 0.00246227
+ 2.806e+11Hz -0.0179852 0.00248535
+ 2.807e+11Hz -0.0179531 0.00250826
+ 2.808e+11Hz -0.0179207 0.00253102
+ 2.809e+11Hz -0.0178879 0.00255361
+ 2.81e+11Hz -0.0178547 0.00257602
+ 2.811e+11Hz -0.0178211 0.00259824
+ 2.812e+11Hz -0.0177872 0.00262028
+ 2.813e+11Hz -0.017753 0.00264213
+ 2.814e+11Hz -0.0177183 0.00266377
+ 2.815e+11Hz -0.0176833 0.0026852
+ 2.816e+11Hz -0.017648 0.00270642
+ 2.817e+11Hz -0.0176123 0.00272742
+ 2.818e+11Hz -0.0175763 0.00274819
+ 2.819e+11Hz -0.0175399 0.00276873
+ 2.82e+11Hz -0.0175032 0.00278903
+ 2.821e+11Hz -0.0174661 0.00280908
+ 2.822e+11Hz -0.0174287 0.00282888
+ 2.823e+11Hz -0.017391 0.00284842
+ 2.824e+11Hz -0.0173529 0.00286769
+ 2.825e+11Hz -0.0173146 0.0028867
+ 2.826e+11Hz -0.0172758 0.00290543
+ 2.827e+11Hz -0.0172368 0.00292387
+ 2.828e+11Hz -0.0171975 0.00294203
+ 2.829e+11Hz -0.0171578 0.00295989
+ 2.83e+11Hz -0.0171178 0.00297745
+ 2.831e+11Hz -0.0170775 0.00299471
+ 2.832e+11Hz -0.0170369 0.00301165
+ 2.833e+11Hz -0.0169961 0.00302828
+ 2.834e+11Hz -0.0169549 0.00304458
+ 2.835e+11Hz -0.0169134 0.00306056
+ 2.836e+11Hz -0.0168717 0.0030762
+ 2.837e+11Hz -0.0168297 0.0030915
+ 2.838e+11Hz -0.0167874 0.00310645
+ 2.839e+11Hz -0.0167448 0.00312106
+ 2.84e+11Hz -0.016702 0.00313531
+ 2.841e+11Hz -0.0166589 0.0031492
+ 2.842e+11Hz -0.0166156 0.00316272
+ 2.843e+11Hz -0.016572 0.00317587
+ 2.844e+11Hz -0.0165281 0.00318865
+ 2.845e+11Hz -0.0164841 0.00320105
+ 2.846e+11Hz -0.0164398 0.00321307
+ 2.847e+11Hz -0.0163952 0.0032247
+ 2.848e+11Hz -0.0163505 0.00323593
+ 2.849e+11Hz -0.0163055 0.00324677
+ 2.85e+11Hz -0.0162604 0.0032572
+ 2.851e+11Hz -0.016215 0.00326723
+ 2.852e+11Hz -0.0161694 0.00327685
+ 2.853e+11Hz -0.0161237 0.00328606
+ 2.854e+11Hz -0.0160777 0.00329485
+ 2.855e+11Hz -0.0160316 0.00330322
+ 2.856e+11Hz -0.0159853 0.00331116
+ 2.857e+11Hz -0.0159389 0.00331868
+ 2.858e+11Hz -0.0158923 0.00332577
+ 2.859e+11Hz -0.0158455 0.00333242
+ 2.86e+11Hz -0.0157986 0.00333863
+ 2.861e+11Hz -0.0157516 0.00334441
+ 2.862e+11Hz -0.0157044 0.00334974
+ 2.863e+11Hz -0.0156571 0.00335463
+ 2.864e+11Hz -0.0156097 0.00335906
+ 2.865e+11Hz -0.0155622 0.00336305
+ 2.866e+11Hz -0.0155146 0.00336659
+ 2.867e+11Hz -0.0154669 0.00336967
+ 2.868e+11Hz -0.0154191 0.00337229
+ 2.869e+11Hz -0.0153712 0.00337446
+ 2.87e+11Hz -0.0153233 0.00337616
+ 2.871e+11Hz -0.0152753 0.00337741
+ 2.872e+11Hz -0.0152272 0.00337819
+ 2.873e+11Hz -0.0151791 0.0033785
+ 2.874e+11Hz -0.0151309 0.00337835
+ 2.875e+11Hz -0.0150827 0.00337774
+ 2.876e+11Hz -0.0150345 0.00337665
+ 2.877e+11Hz -0.0149863 0.0033751
+ 2.878e+11Hz -0.014938 0.00337308
+ 2.879e+11Hz -0.0148898 0.00337059
+ 2.88e+11Hz -0.0148415 0.00336763
+ 2.881e+11Hz -0.0147933 0.0033642
+ 2.882e+11Hz -0.0147451 0.0033603
+ 2.883e+11Hz -0.0146969 0.00335593
+ 2.884e+11Hz -0.0146487 0.00335109
+ 2.885e+11Hz -0.0146006 0.00334578
+ 2.886e+11Hz -0.0145525 0.00334001
+ 2.887e+11Hz -0.0145045 0.00333376
+ 2.888e+11Hz -0.0144566 0.00332705
+ 2.889e+11Hz -0.0144087 0.00331988
+ 2.89e+11Hz -0.0143609 0.00331224
+ 2.891e+11Hz -0.0143132 0.00330414
+ 2.892e+11Hz -0.0142656 0.00329557
+ 2.893e+11Hz -0.0142181 0.00328655
+ 2.894e+11Hz -0.0141707 0.00327707
+ 2.895e+11Hz -0.0141234 0.00326713
+ 2.896e+11Hz -0.0140763 0.00325674
+ 2.897e+11Hz -0.0140293 0.0032459
+ 2.898e+11Hz -0.0139824 0.00323461
+ 2.899e+11Hz -0.0139357 0.00322287
+ 2.9e+11Hz -0.0138891 0.00321068
+ 2.901e+11Hz -0.0138427 0.00319805
+ 2.902e+11Hz -0.0137964 0.00318499
+ 2.903e+11Hz -0.0137504 0.00317149
+ 2.904e+11Hz -0.0137045 0.00315756
+ 2.905e+11Hz -0.0136588 0.0031432
+ 2.906e+11Hz -0.0136133 0.00312841
+ 2.907e+11Hz -0.013568 0.0031132
+ 2.908e+11Hz -0.0135229 0.00309757
+ 2.909e+11Hz -0.013478 0.00308153
+ 2.91e+11Hz -0.0134334 0.00306507
+ 2.911e+11Hz -0.013389 0.00304821
+ 2.912e+11Hz -0.0133448 0.00303095
+ 2.913e+11Hz -0.0133009 0.00301329
+ 2.914e+11Hz -0.0132572 0.00299524
+ 2.915e+11Hz -0.0132138 0.0029768
+ 2.916e+11Hz -0.0131706 0.00295797
+ 2.917e+11Hz -0.0131277 0.00293877
+ 2.918e+11Hz -0.0130851 0.00291919
+ 2.919e+11Hz -0.0130427 0.00289924
+ 2.92e+11Hz -0.0130007 0.00287893
+ 2.921e+11Hz -0.0129589 0.00285826
+ 2.922e+11Hz -0.0129174 0.00283723
+ 2.923e+11Hz -0.0128763 0.00281586
+ 2.924e+11Hz -0.0128354 0.00279415
+ 2.925e+11Hz -0.0127949 0.0027721
+ 2.926e+11Hz -0.0127546 0.00274972
+ 2.927e+11Hz -0.0127147 0.00272701
+ 2.928e+11Hz -0.0126751 0.00270398
+ 2.929e+11Hz -0.0126359 0.00268065
+ 2.93e+11Hz -0.012597 0.002657
+ 2.931e+11Hz -0.0125584 0.00263305
+ 2.932e+11Hz -0.0125202 0.00260882
+ 2.933e+11Hz -0.0124823 0.00258429
+ 2.934e+11Hz -0.0124448 0.00255948
+ 2.935e+11Hz -0.0124076 0.0025344
+ 2.936e+11Hz -0.0123708 0.00250904
+ 2.937e+11Hz -0.0123344 0.00248343
+ 2.938e+11Hz -0.0122983 0.00245756
+ 2.939e+11Hz -0.0122626 0.00243145
+ 2.94e+11Hz -0.0122273 0.00240509
+ 2.941e+11Hz -0.0121923 0.0023785
+ 2.942e+11Hz -0.0121578 0.00235168
+ 2.943e+11Hz -0.0121236 0.00232464
+ 2.944e+11Hz -0.0120898 0.00229738
+ 2.945e+11Hz -0.0120564 0.00226993
+ 2.946e+11Hz -0.0120234 0.00224227
+ 2.947e+11Hz -0.0119908 0.00221442
+ 2.948e+11Hz -0.0119585 0.00218638
+ 2.949e+11Hz -0.0119267 0.00215817
+ 2.95e+11Hz -0.0118953 0.00212979
+ 2.951e+11Hz -0.0118642 0.00210124
+ 2.952e+11Hz -0.0118336 0.00207254
+ 2.953e+11Hz -0.0118034 0.00204369
+ 2.954e+11Hz -0.0117736 0.0020147
+ 2.955e+11Hz -0.0117442 0.00198558
+ 2.956e+11Hz -0.0117152 0.00195633
+ 2.957e+11Hz -0.0116866 0.00192696
+ 2.958e+11Hz -0.0116584 0.00189747
+ 2.959e+11Hz -0.0116306 0.00186789
+ 2.96e+11Hz -0.0116033 0.0018382
+ 2.961e+11Hz -0.0115763 0.00180843
+ 2.962e+11Hz -0.0115498 0.00177858
+ 2.963e+11Hz -0.0115237 0.00174865
+ 2.964e+11Hz -0.0114979 0.00171865
+ 2.965e+11Hz -0.0114726 0.00168859
+ 2.966e+11Hz -0.0114477 0.00165848
+ 2.967e+11Hz -0.0114232 0.00162832
+ 2.968e+11Hz -0.0113991 0.00159812
+ 2.969e+11Hz -0.0113754 0.00156789
+ 2.97e+11Hz -0.0113522 0.00153764
+ 2.971e+11Hz -0.0113293 0.00150737
+ 2.972e+11Hz -0.0113068 0.00147708
+ 2.973e+11Hz -0.0112848 0.0014468
+ 2.974e+11Hz -0.0112631 0.00141651
+ 2.975e+11Hz -0.0112418 0.00138624
+ 2.976e+11Hz -0.0112209 0.00135598
+ 2.977e+11Hz -0.0112004 0.00132575
+ 2.978e+11Hz -0.0111804 0.00129555
+ 2.979e+11Hz -0.0111607 0.00126538
+ 2.98e+11Hz -0.0111413 0.00123526
+ 2.981e+11Hz -0.0111224 0.00120519
+ 2.982e+11Hz -0.0111039 0.00117517
+ 2.983e+11Hz -0.0110857 0.00114522
+ 2.984e+11Hz -0.0110679 0.00111534
+ 2.985e+11Hz -0.0110505 0.00108553
+ 2.986e+11Hz -0.0110334 0.0010558
+ 2.987e+11Hz -0.0110167 0.00102616
+ 2.988e+11Hz -0.0110004 0.000996611
+ 2.989e+11Hz -0.0109844 0.000967163
+ 2.99e+11Hz -0.0109688 0.000937819
+ 2.991e+11Hz -0.0109536 0.000908586
+ 2.992e+11Hz -0.0109387 0.000879469
+ 2.993e+11Hz -0.0109241 0.000850473
+ 2.994e+11Hz -0.0109099 0.000821604
+ 2.995e+11Hz -0.010896 0.000792867
+ 2.996e+11Hz -0.0108824 0.000764267
+ 2.997e+11Hz -0.0108692 0.00073581
+ 2.998e+11Hz -0.0108563 0.000707499
+ 2.999e+11Hz -0.0108437 0.000679341
+ 3e+11Hz -0.0108314 0.00065134
+ ]

A12 %vd(20 3) %vd(12, 3) xfer2
.model xfer2 xfer R_I=true table=[
+ 0Hz 0.995436 0
+ 1e+08Hz 0.995435 -0.000814178
+ 2e+08Hz 0.995433 -0.00162834
+ 3e+08Hz 0.99543 -0.00244247
+ 4e+08Hz 0.995425 -0.00325656
+ 5e+08Hz 0.99542 -0.00407058
+ 6e+08Hz 0.995412 -0.00488452
+ 7e+08Hz 0.995404 -0.00569837
+ 8e+08Hz 0.995394 -0.00651211
+ 9e+08Hz 0.995383 -0.00732573
+ 1e+09Hz 0.995371 -0.0081392
+ 1.1e+09Hz 0.995358 -0.00895252
+ 1.2e+09Hz 0.995343 -0.00976567
+ 1.3e+09Hz 0.995327 -0.0105786
+ 1.4e+09Hz 0.99531 -0.0113914
+ 1.5e+09Hz 0.995291 -0.012204
+ 1.6e+09Hz 0.995271 -0.0130163
+ 1.7e+09Hz 0.99525 -0.0138284
+ 1.8e+09Hz 0.995228 -0.0146402
+ 1.9e+09Hz 0.995204 -0.0154517
+ 2e+09Hz 0.99518 -0.016263
+ 2.1e+09Hz 0.995154 -0.017074
+ 2.2e+09Hz 0.995126 -0.0178846
+ 2.3e+09Hz 0.995098 -0.0186949
+ 2.4e+09Hz 0.995068 -0.0195049
+ 2.5e+09Hz 0.995038 -0.0203146
+ 2.6e+09Hz 0.995006 -0.0211238
+ 2.7e+09Hz 0.994973 -0.0219327
+ 2.8e+09Hz 0.994938 -0.0227412
+ 2.9e+09Hz 0.994903 -0.0235493
+ 3e+09Hz 0.994866 -0.024357
+ 3.1e+09Hz 0.994829 -0.0251643
+ 3.2e+09Hz 0.99479 -0.0259711
+ 3.3e+09Hz 0.99475 -0.0267775
+ 3.4e+09Hz 0.994709 -0.0275834
+ 3.5e+09Hz 0.994667 -0.0283889
+ 3.6e+09Hz 0.994624 -0.0291939
+ 3.7e+09Hz 0.994579 -0.0299984
+ 3.8e+09Hz 0.994534 -0.0308024
+ 3.9e+09Hz 0.994488 -0.031606
+ 4e+09Hz 0.994441 -0.032409
+ 4.1e+09Hz 0.994392 -0.0332114
+ 4.2e+09Hz 0.994343 -0.0340134
+ 4.3e+09Hz 0.994292 -0.0348148
+ 4.4e+09Hz 0.994241 -0.0356157
+ 4.5e+09Hz 0.994189 -0.036416
+ 4.6e+09Hz 0.994136 -0.0372158
+ 4.7e+09Hz 0.994081 -0.038015
+ 4.8e+09Hz 0.994026 -0.0388137
+ 4.9e+09Hz 0.99397 -0.0396118
+ 5e+09Hz 0.993913 -0.0404093
+ 5.1e+09Hz 0.993856 -0.0412062
+ 5.2e+09Hz 0.993797 -0.0420026
+ 5.3e+09Hz 0.993737 -0.0427983
+ 5.4e+09Hz 0.993677 -0.0435935
+ 5.5e+09Hz 0.993616 -0.044388
+ 5.6e+09Hz 0.993554 -0.045182
+ 5.7e+09Hz 0.993491 -0.0459753
+ 5.8e+09Hz 0.993427 -0.0467681
+ 5.9e+09Hz 0.993363 -0.0475602
+ 6e+09Hz 0.993298 -0.0483518
+ 6.1e+09Hz 0.993232 -0.0491427
+ 6.2e+09Hz 0.993165 -0.049933
+ 6.3e+09Hz 0.993098 -0.0507227
+ 6.4e+09Hz 0.99303 -0.0515118
+ 6.5e+09Hz 0.992961 -0.0523003
+ 6.6e+09Hz 0.992892 -0.0530882
+ 6.7e+09Hz 0.992821 -0.0538755
+ 6.8e+09Hz 0.992751 -0.0546622
+ 6.9e+09Hz 0.992679 -0.0554482
+ 7e+09Hz 0.992607 -0.0562337
+ 7.1e+09Hz 0.992535 -0.0570185
+ 7.2e+09Hz 0.992461 -0.0578028
+ 7.3e+09Hz 0.992387 -0.0585865
+ 7.4e+09Hz 0.992313 -0.0593695
+ 7.5e+09Hz 0.992238 -0.060152
+ 7.6e+09Hz 0.992162 -0.0609339
+ 7.7e+09Hz 0.992086 -0.0617152
+ 7.8e+09Hz 0.99201 -0.062496
+ 7.9e+09Hz 0.991933 -0.0632762
+ 8e+09Hz 0.991855 -0.0640558
+ 8.1e+09Hz 0.991777 -0.0648348
+ 8.2e+09Hz 0.991698 -0.0656133
+ 8.3e+09Hz 0.991619 -0.0663912
+ 8.4e+09Hz 0.99154 -0.0671686
+ 8.5e+09Hz 0.991459 -0.0679455
+ 8.6e+09Hz 0.991379 -0.0687218
+ 8.7e+09Hz 0.991298 -0.0694976
+ 8.8e+09Hz 0.991217 -0.0702728
+ 8.9e+09Hz 0.991135 -0.0710476
+ 9e+09Hz 0.991053 -0.0718218
+ 9.1e+09Hz 0.99097 -0.0725956
+ 9.2e+09Hz 0.990888 -0.0733689
+ 9.3e+09Hz 0.990804 -0.0741417
+ 9.4e+09Hz 0.990721 -0.074914
+ 9.5e+09Hz 0.990637 -0.0756858
+ 9.6e+09Hz 0.990552 -0.0764572
+ 9.7e+09Hz 0.990467 -0.0772282
+ 9.8e+09Hz 0.990382 -0.0779987
+ 9.9e+09Hz 0.990297 -0.0787687
+ 1e+10Hz 0.990211 -0.0795384
+ 1.01e+10Hz 0.990125 -0.0803076
+ 1.02e+10Hz 0.990039 -0.0810764
+ 1.03e+10Hz 0.989952 -0.0818449
+ 1.04e+10Hz 0.989865 -0.0826129
+ 1.05e+10Hz 0.989778 -0.0833806
+ 1.06e+10Hz 0.98969 -0.0841479
+ 1.07e+10Hz 0.989603 -0.0849148
+ 1.08e+10Hz 0.989514 -0.0856814
+ 1.09e+10Hz 0.989426 -0.0864477
+ 1.1e+10Hz 0.989337 -0.0872136
+ 1.11e+10Hz 0.989248 -0.0879793
+ 1.12e+10Hz 0.989159 -0.0887446
+ 1.13e+10Hz 0.98907 -0.0895096
+ 1.14e+10Hz 0.98898 -0.0902743
+ 1.15e+10Hz 0.98889 -0.0910387
+ 1.16e+10Hz 0.9888 -0.0918029
+ 1.17e+10Hz 0.988709 -0.0925668
+ 1.18e+10Hz 0.988618 -0.0933304
+ 1.19e+10Hz 0.988527 -0.0940938
+ 1.2e+10Hz 0.988436 -0.094857
+ 1.21e+10Hz 0.988344 -0.09562
+ 1.22e+10Hz 0.988253 -0.0963827
+ 1.23e+10Hz 0.988161 -0.0971453
+ 1.24e+10Hz 0.988068 -0.0979076
+ 1.25e+10Hz 0.987976 -0.0986698
+ 1.26e+10Hz 0.987883 -0.0994318
+ 1.27e+10Hz 0.98779 -0.100194
+ 1.28e+10Hz 0.987697 -0.100955
+ 1.29e+10Hz 0.987603 -0.101717
+ 1.3e+10Hz 0.987509 -0.102478
+ 1.31e+10Hz 0.987415 -0.10324
+ 1.32e+10Hz 0.987321 -0.104001
+ 1.33e+10Hz 0.987226 -0.104762
+ 1.34e+10Hz 0.987131 -0.105523
+ 1.35e+10Hz 0.987036 -0.106283
+ 1.36e+10Hz 0.986941 -0.107044
+ 1.37e+10Hz 0.986845 -0.107805
+ 1.38e+10Hz 0.986749 -0.108566
+ 1.39e+10Hz 0.986653 -0.109326
+ 1.4e+10Hz 0.986556 -0.110087
+ 1.41e+10Hz 0.986459 -0.110847
+ 1.42e+10Hz 0.986362 -0.111607
+ 1.43e+10Hz 0.986265 -0.112368
+ 1.44e+10Hz 0.986167 -0.113128
+ 1.45e+10Hz 0.986069 -0.113888
+ 1.46e+10Hz 0.985971 -0.114649
+ 1.47e+10Hz 0.985872 -0.115409
+ 1.48e+10Hz 0.985773 -0.116169
+ 1.49e+10Hz 0.985673 -0.11693
+ 1.5e+10Hz 0.985574 -0.11769
+ 1.51e+10Hz 0.985474 -0.11845
+ 1.52e+10Hz 0.985373 -0.119211
+ 1.53e+10Hz 0.985273 -0.119971
+ 1.54e+10Hz 0.985172 -0.120732
+ 1.55e+10Hz 0.98507 -0.121492
+ 1.56e+10Hz 0.984968 -0.122253
+ 1.57e+10Hz 0.984866 -0.123013
+ 1.58e+10Hz 0.984763 -0.123774
+ 1.59e+10Hz 0.98466 -0.124535
+ 1.6e+10Hz 0.984557 -0.125295
+ 1.61e+10Hz 0.984453 -0.126056
+ 1.62e+10Hz 0.984349 -0.126817
+ 1.63e+10Hz 0.984244 -0.127578
+ 1.64e+10Hz 0.984139 -0.128339
+ 1.65e+10Hz 0.984034 -0.1291
+ 1.66e+10Hz 0.983928 -0.129861
+ 1.67e+10Hz 0.983822 -0.130623
+ 1.68e+10Hz 0.983715 -0.131384
+ 1.69e+10Hz 0.983607 -0.132145
+ 1.7e+10Hz 0.9835 -0.132907
+ 1.71e+10Hz 0.983391 -0.133669
+ 1.72e+10Hz 0.983283 -0.13443
+ 1.73e+10Hz 0.983174 -0.135192
+ 1.74e+10Hz 0.983064 -0.135954
+ 1.75e+10Hz 0.982954 -0.136716
+ 1.76e+10Hz 0.982843 -0.137478
+ 1.77e+10Hz 0.982732 -0.13824
+ 1.78e+10Hz 0.98262 -0.139002
+ 1.79e+10Hz 0.982508 -0.139765
+ 1.8e+10Hz 0.982395 -0.140527
+ 1.81e+10Hz 0.982281 -0.14129
+ 1.82e+10Hz 0.982167 -0.142052
+ 1.83e+10Hz 0.982053 -0.142815
+ 1.84e+10Hz 0.981938 -0.143578
+ 1.85e+10Hz 0.981822 -0.14434
+ 1.86e+10Hz 0.981706 -0.145103
+ 1.87e+10Hz 0.981589 -0.145866
+ 1.88e+10Hz 0.981472 -0.146629
+ 1.89e+10Hz 0.981354 -0.147393
+ 1.9e+10Hz 0.981235 -0.148156
+ 1.91e+10Hz 0.981116 -0.148919
+ 1.92e+10Hz 0.980996 -0.149682
+ 1.93e+10Hz 0.980876 -0.150446
+ 1.94e+10Hz 0.980754 -0.151209
+ 1.95e+10Hz 0.980633 -0.151973
+ 1.96e+10Hz 0.98051 -0.152736
+ 1.97e+10Hz 0.980387 -0.1535
+ 1.98e+10Hz 0.980264 -0.154264
+ 1.99e+10Hz 0.980139 -0.155027
+ 2e+10Hz 0.980014 -0.155791
+ 2.01e+10Hz 0.979889 -0.156555
+ 2.02e+10Hz 0.979762 -0.157319
+ 2.03e+10Hz 0.979635 -0.158083
+ 2.04e+10Hz 0.979508 -0.158846
+ 2.05e+10Hz 0.979379 -0.15961
+ 2.06e+10Hz 0.97925 -0.160374
+ 2.07e+10Hz 0.979121 -0.161138
+ 2.08e+10Hz 0.97899 -0.161902
+ 2.09e+10Hz 0.978859 -0.162666
+ 2.1e+10Hz 0.978727 -0.16343
+ 2.11e+10Hz 0.978595 -0.164193
+ 2.12e+10Hz 0.978461 -0.164957
+ 2.13e+10Hz 0.978327 -0.165721
+ 2.14e+10Hz 0.978193 -0.166485
+ 2.15e+10Hz 0.978057 -0.167249
+ 2.16e+10Hz 0.977921 -0.168012
+ 2.17e+10Hz 0.977785 -0.168776
+ 2.18e+10Hz 0.977647 -0.169539
+ 2.19e+10Hz 0.977509 -0.170303
+ 2.2e+10Hz 0.97737 -0.171066
+ 2.21e+10Hz 0.97723 -0.17183
+ 2.22e+10Hz 0.97709 -0.172593
+ 2.23e+10Hz 0.976948 -0.173356
+ 2.24e+10Hz 0.976807 -0.174119
+ 2.25e+10Hz 0.976664 -0.174882
+ 2.26e+10Hz 0.976521 -0.175645
+ 2.27e+10Hz 0.976377 -0.176408
+ 2.28e+10Hz 0.976232 -0.17717
+ 2.29e+10Hz 0.976086 -0.177933
+ 2.3e+10Hz 0.97594 -0.178695
+ 2.31e+10Hz 0.975793 -0.179458
+ 2.32e+10Hz 0.975645 -0.18022
+ 2.33e+10Hz 0.975497 -0.180982
+ 2.34e+10Hz 0.975348 -0.181743
+ 2.35e+10Hz 0.975198 -0.182505
+ 2.36e+10Hz 0.975047 -0.183267
+ 2.37e+10Hz 0.974896 -0.184028
+ 2.38e+10Hz 0.974744 -0.184789
+ 2.39e+10Hz 0.974591 -0.18555
+ 2.4e+10Hz 0.974438 -0.186311
+ 2.41e+10Hz 0.974284 -0.187072
+ 2.42e+10Hz 0.974129 -0.187832
+ 2.43e+10Hz 0.973973 -0.188592
+ 2.44e+10Hz 0.973817 -0.189352
+ 2.45e+10Hz 0.97366 -0.190112
+ 2.46e+10Hz 0.973502 -0.190872
+ 2.47e+10Hz 0.973344 -0.191631
+ 2.48e+10Hz 0.973185 -0.19239
+ 2.49e+10Hz 0.973025 -0.193149
+ 2.5e+10Hz 0.972864 -0.193908
+ 2.51e+10Hz 0.972703 -0.194667
+ 2.52e+10Hz 0.972541 -0.195425
+ 2.53e+10Hz 0.972379 -0.196183
+ 2.54e+10Hz 0.972216 -0.196941
+ 2.55e+10Hz 0.972052 -0.197698
+ 2.56e+10Hz 0.971887 -0.198455
+ 2.57e+10Hz 0.971722 -0.199212
+ 2.58e+10Hz 0.971556 -0.199969
+ 2.59e+10Hz 0.97139 -0.200726
+ 2.6e+10Hz 0.971223 -0.201482
+ 2.61e+10Hz 0.971055 -0.202238
+ 2.62e+10Hz 0.970886 -0.202994
+ 2.63e+10Hz 0.970717 -0.203749
+ 2.64e+10Hz 0.970548 -0.204504
+ 2.65e+10Hz 0.970377 -0.205259
+ 2.66e+10Hz 0.970206 -0.206014
+ 2.67e+10Hz 0.970035 -0.206768
+ 2.68e+10Hz 0.969863 -0.207522
+ 2.69e+10Hz 0.96969 -0.208276
+ 2.7e+10Hz 0.969516 -0.209029
+ 2.71e+10Hz 0.969342 -0.209782
+ 2.72e+10Hz 0.969168 -0.210535
+ 2.73e+10Hz 0.968993 -0.211288
+ 2.74e+10Hz 0.968817 -0.21204
+ 2.75e+10Hz 0.968641 -0.212792
+ 2.76e+10Hz 0.968464 -0.213544
+ 2.77e+10Hz 0.968286 -0.214296
+ 2.78e+10Hz 0.968108 -0.215047
+ 2.79e+10Hz 0.96793 -0.215798
+ 2.8e+10Hz 0.96775 -0.216548
+ 2.81e+10Hz 0.967571 -0.217298
+ 2.82e+10Hz 0.96739 -0.218048
+ 2.83e+10Hz 0.96721 -0.218798
+ 2.84e+10Hz 0.967028 -0.219548
+ 2.85e+10Hz 0.966846 -0.220297
+ 2.86e+10Hz 0.966664 -0.221046
+ 2.87e+10Hz 0.966481 -0.221794
+ 2.88e+10Hz 0.966298 -0.222542
+ 2.89e+10Hz 0.966114 -0.22329
+ 2.9e+10Hz 0.965929 -0.224038
+ 2.91e+10Hz 0.965744 -0.224785
+ 2.92e+10Hz 0.965559 -0.225533
+ 2.93e+10Hz 0.965373 -0.22628
+ 2.94e+10Hz 0.965186 -0.227026
+ 2.95e+10Hz 0.964999 -0.227772
+ 2.96e+10Hz 0.964812 -0.228519
+ 2.97e+10Hz 0.964624 -0.229264
+ 2.98e+10Hz 0.964435 -0.23001
+ 2.99e+10Hz 0.964246 -0.230755
+ 3e+10Hz 0.964057 -0.2315
+ 3.01e+10Hz 0.963867 -0.232245
+ 3.02e+10Hz 0.963677 -0.232989
+ 3.03e+10Hz 0.963486 -0.233734
+ 3.04e+10Hz 0.963295 -0.234478
+ 3.05e+10Hz 0.963103 -0.235221
+ 3.06e+10Hz 0.962911 -0.235965
+ 3.07e+10Hz 0.962718 -0.236708
+ 3.08e+10Hz 0.962525 -0.237451
+ 3.09e+10Hz 0.962332 -0.238194
+ 3.1e+10Hz 0.962138 -0.238936
+ 3.11e+10Hz 0.961943 -0.239679
+ 3.12e+10Hz 0.961748 -0.240421
+ 3.13e+10Hz 0.961553 -0.241163
+ 3.14e+10Hz 0.961357 -0.241905
+ 3.15e+10Hz 0.961161 -0.242646
+ 3.16e+10Hz 0.960964 -0.243387
+ 3.17e+10Hz 0.960767 -0.244128
+ 3.18e+10Hz 0.96057 -0.244869
+ 3.19e+10Hz 0.960372 -0.24561
+ 3.2e+10Hz 0.960174 -0.24635
+ 3.21e+10Hz 0.959975 -0.247091
+ 3.22e+10Hz 0.959775 -0.247831
+ 3.23e+10Hz 0.959576 -0.248571
+ 3.24e+10Hz 0.959376 -0.24931
+ 3.25e+10Hz 0.959175 -0.25005
+ 3.26e+10Hz 0.958974 -0.250789
+ 3.27e+10Hz 0.958773 -0.251528
+ 3.28e+10Hz 0.958571 -0.252267
+ 3.29e+10Hz 0.958369 -0.253006
+ 3.3e+10Hz 0.958166 -0.253745
+ 3.31e+10Hz 0.957963 -0.254484
+ 3.32e+10Hz 0.95776 -0.255222
+ 3.33e+10Hz 0.957556 -0.25596
+ 3.34e+10Hz 0.957351 -0.256698
+ 3.35e+10Hz 0.957146 -0.257436
+ 3.36e+10Hz 0.956941 -0.258174
+ 3.37e+10Hz 0.956735 -0.258912
+ 3.38e+10Hz 0.956529 -0.25965
+ 3.39e+10Hz 0.956323 -0.260387
+ 3.4e+10Hz 0.956116 -0.261125
+ 3.41e+10Hz 0.955908 -0.261862
+ 3.42e+10Hz 0.9557 -0.262599
+ 3.43e+10Hz 0.955492 -0.263336
+ 3.44e+10Hz 0.955283 -0.264073
+ 3.45e+10Hz 0.955074 -0.26481
+ 3.46e+10Hz 0.954864 -0.265546
+ 3.47e+10Hz 0.954654 -0.266283
+ 3.48e+10Hz 0.954443 -0.26702
+ 3.49e+10Hz 0.954232 -0.267756
+ 3.5e+10Hz 0.954021 -0.268492
+ 3.51e+10Hz 0.953809 -0.269228
+ 3.52e+10Hz 0.953596 -0.269965
+ 3.53e+10Hz 0.953383 -0.270701
+ 3.54e+10Hz 0.95317 -0.271437
+ 3.55e+10Hz 0.952956 -0.272173
+ 3.56e+10Hz 0.952742 -0.272908
+ 3.57e+10Hz 0.952527 -0.273644
+ 3.58e+10Hz 0.952312 -0.27438
+ 3.59e+10Hz 0.952096 -0.275115
+ 3.6e+10Hz 0.951879 -0.275851
+ 3.61e+10Hz 0.951663 -0.276586
+ 3.62e+10Hz 0.951445 -0.277322
+ 3.63e+10Hz 0.951227 -0.278057
+ 3.64e+10Hz 0.951009 -0.278792
+ 3.65e+10Hz 0.95079 -0.279528
+ 3.66e+10Hz 0.950571 -0.280263
+ 3.67e+10Hz 0.950351 -0.280998
+ 3.68e+10Hz 0.950131 -0.281733
+ 3.69e+10Hz 0.94991 -0.282468
+ 3.7e+10Hz 0.949689 -0.283203
+ 3.71e+10Hz 0.949467 -0.283938
+ 3.72e+10Hz 0.949244 -0.284672
+ 3.73e+10Hz 0.949021 -0.285407
+ 3.74e+10Hz 0.948798 -0.286142
+ 3.75e+10Hz 0.948574 -0.286876
+ 3.76e+10Hz 0.948349 -0.287611
+ 3.77e+10Hz 0.948124 -0.288345
+ 3.78e+10Hz 0.947898 -0.28908
+ 3.79e+10Hz 0.947672 -0.289814
+ 3.8e+10Hz 0.947445 -0.290549
+ 3.81e+10Hz 0.947218 -0.291283
+ 3.82e+10Hz 0.94699 -0.292017
+ 3.83e+10Hz 0.946761 -0.292751
+ 3.84e+10Hz 0.946532 -0.293485
+ 3.85e+10Hz 0.946302 -0.294219
+ 3.86e+10Hz 0.946072 -0.294953
+ 3.87e+10Hz 0.945841 -0.295687
+ 3.88e+10Hz 0.94561 -0.296421
+ 3.89e+10Hz 0.945377 -0.297154
+ 3.9e+10Hz 0.945145 -0.297888
+ 3.91e+10Hz 0.944912 -0.298622
+ 3.92e+10Hz 0.944678 -0.299355
+ 3.93e+10Hz 0.944443 -0.300088
+ 3.94e+10Hz 0.944208 -0.300822
+ 3.95e+10Hz 0.943972 -0.301555
+ 3.96e+10Hz 0.943736 -0.302288
+ 3.97e+10Hz 0.943499 -0.303021
+ 3.98e+10Hz 0.943262 -0.303754
+ 3.99e+10Hz 0.943023 -0.304487
+ 4e+10Hz 0.942785 -0.30522
+ 4.01e+10Hz 0.942545 -0.305953
+ 4.02e+10Hz 0.942305 -0.306685
+ 4.03e+10Hz 0.942065 -0.307418
+ 4.04e+10Hz 0.941823 -0.30815
+ 4.05e+10Hz 0.941581 -0.308882
+ 4.06e+10Hz 0.941339 -0.309615
+ 4.07e+10Hz 0.941095 -0.310347
+ 4.08e+10Hz 0.940851 -0.311079
+ 4.09e+10Hz 0.940607 -0.31181
+ 4.1e+10Hz 0.940362 -0.312542
+ 4.11e+10Hz 0.940116 -0.313274
+ 4.12e+10Hz 0.939869 -0.314005
+ 4.13e+10Hz 0.939622 -0.314736
+ 4.14e+10Hz 0.939374 -0.315468
+ 4.15e+10Hz 0.939126 -0.316199
+ 4.16e+10Hz 0.938877 -0.316929
+ 4.17e+10Hz 0.938627 -0.31766
+ 4.18e+10Hz 0.938377 -0.318391
+ 4.19e+10Hz 0.938126 -0.319121
+ 4.2e+10Hz 0.937874 -0.319851
+ 4.21e+10Hz 0.937621 -0.320581
+ 4.22e+10Hz 0.937368 -0.321311
+ 4.23e+10Hz 0.937114 -0.322041
+ 4.24e+10Hz 0.93686 -0.322771
+ 4.25e+10Hz 0.936605 -0.3235
+ 4.26e+10Hz 0.936349 -0.324229
+ 4.27e+10Hz 0.936093 -0.324958
+ 4.28e+10Hz 0.935836 -0.325687
+ 4.29e+10Hz 0.935578 -0.326416
+ 4.3e+10Hz 0.935319 -0.327144
+ 4.31e+10Hz 0.93506 -0.327872
+ 4.32e+10Hz 0.934801 -0.328601
+ 4.33e+10Hz 0.93454 -0.329328
+ 4.34e+10Hz 0.934279 -0.330056
+ 4.35e+10Hz 0.934017 -0.330783
+ 4.36e+10Hz 0.933755 -0.331511
+ 4.37e+10Hz 0.933492 -0.332238
+ 4.38e+10Hz 0.933228 -0.332964
+ 4.39e+10Hz 0.932964 -0.333691
+ 4.4e+10Hz 0.932698 -0.334417
+ 4.41e+10Hz 0.932433 -0.335143
+ 4.42e+10Hz 0.932166 -0.335869
+ 4.43e+10Hz 0.931899 -0.336594
+ 4.44e+10Hz 0.931632 -0.33732
+ 4.45e+10Hz 0.931363 -0.338045
+ 4.46e+10Hz 0.931094 -0.338769
+ 4.47e+10Hz 0.930825 -0.339494
+ 4.48e+10Hz 0.930554 -0.340218
+ 4.49e+10Hz 0.930283 -0.340942
+ 4.5e+10Hz 0.930012 -0.341666
+ 4.51e+10Hz 0.929739 -0.342389
+ 4.52e+10Hz 0.929467 -0.343113
+ 4.53e+10Hz 0.929193 -0.343836
+ 4.54e+10Hz 0.928919 -0.344558
+ 4.55e+10Hz 0.928644 -0.345281
+ 4.56e+10Hz 0.928369 -0.346003
+ 4.57e+10Hz 0.928093 -0.346724
+ 4.58e+10Hz 0.927816 -0.347446
+ 4.59e+10Hz 0.927539 -0.348167
+ 4.6e+10Hz 0.927261 -0.348888
+ 4.61e+10Hz 0.926982 -0.349609
+ 4.62e+10Hz 0.926703 -0.350329
+ 4.63e+10Hz 0.926423 -0.351049
+ 4.64e+10Hz 0.926143 -0.351769
+ 4.65e+10Hz 0.925862 -0.352488
+ 4.66e+10Hz 0.92558 -0.353207
+ 4.67e+10Hz 0.925298 -0.353926
+ 4.68e+10Hz 0.925015 -0.354644
+ 4.69e+10Hz 0.924732 -0.355362
+ 4.7e+10Hz 0.924448 -0.35608
+ 4.71e+10Hz 0.924163 -0.356798
+ 4.72e+10Hz 0.923878 -0.357515
+ 4.73e+10Hz 0.923592 -0.358232
+ 4.74e+10Hz 0.923306 -0.358949
+ 4.75e+10Hz 0.923019 -0.359665
+ 4.76e+10Hz 0.922732 -0.360381
+ 4.77e+10Hz 0.922444 -0.361096
+ 4.78e+10Hz 0.922155 -0.361812
+ 4.79e+10Hz 0.921866 -0.362527
+ 4.8e+10Hz 0.921576 -0.363241
+ 4.81e+10Hz 0.921286 -0.363955
+ 4.82e+10Hz 0.920995 -0.364669
+ 4.83e+10Hz 0.920704 -0.365383
+ 4.84e+10Hz 0.920412 -0.366096
+ 4.85e+10Hz 0.920119 -0.366809
+ 4.86e+10Hz 0.919826 -0.367522
+ 4.87e+10Hz 0.919532 -0.368234
+ 4.88e+10Hz 0.919238 -0.368946
+ 4.89e+10Hz 0.918944 -0.369658
+ 4.9e+10Hz 0.918649 -0.37037
+ 4.91e+10Hz 0.918353 -0.371081
+ 4.92e+10Hz 0.918057 -0.371791
+ 4.93e+10Hz 0.91776 -0.372502
+ 4.94e+10Hz 0.917463 -0.373212
+ 4.95e+10Hz 0.917165 -0.373922
+ 4.96e+10Hz 0.916866 -0.374631
+ 4.97e+10Hz 0.916568 -0.37534
+ 4.98e+10Hz 0.916268 -0.376049
+ 4.99e+10Hz 0.915969 -0.376757
+ 5e+10Hz 0.915668 -0.377465
+ 5.01e+10Hz 0.915367 -0.378173
+ 5.02e+10Hz 0.915066 -0.378881
+ 5.03e+10Hz 0.914764 -0.379588
+ 5.04e+10Hz 0.914462 -0.380295
+ 5.05e+10Hz 0.914159 -0.381002
+ 5.06e+10Hz 0.913856 -0.381708
+ 5.07e+10Hz 0.913552 -0.382414
+ 5.08e+10Hz 0.913248 -0.383119
+ 5.09e+10Hz 0.912943 -0.383825
+ 5.1e+10Hz 0.912638 -0.38453
+ 5.11e+10Hz 0.912332 -0.385234
+ 5.12e+10Hz 0.912026 -0.385939
+ 5.13e+10Hz 0.91172 -0.386643
+ 5.14e+10Hz 0.911412 -0.387347
+ 5.15e+10Hz 0.911105 -0.38805
+ 5.16e+10Hz 0.910797 -0.388754
+ 5.17e+10Hz 0.910488 -0.389457
+ 5.18e+10Hz 0.910179 -0.390159
+ 5.19e+10Hz 0.90987 -0.390862
+ 5.2e+10Hz 0.90956 -0.391564
+ 5.21e+10Hz 0.90925 -0.392266
+ 5.22e+10Hz 0.908939 -0.392967
+ 5.23e+10Hz 0.908628 -0.393668
+ 5.24e+10Hz 0.908316 -0.394369
+ 5.25e+10Hz 0.908004 -0.39507
+ 5.26e+10Hz 0.907691 -0.395771
+ 5.27e+10Hz 0.907378 -0.396471
+ 5.28e+10Hz 0.907065 -0.397171
+ 5.29e+10Hz 0.906751 -0.39787
+ 5.3e+10Hz 0.906436 -0.39857
+ 5.31e+10Hz 0.906121 -0.399269
+ 5.32e+10Hz 0.905806 -0.399968
+ 5.33e+10Hz 0.90549 -0.400666
+ 5.34e+10Hz 0.905174 -0.401365
+ 5.35e+10Hz 0.904857 -0.402063
+ 5.36e+10Hz 0.90454 -0.402761
+ 5.37e+10Hz 0.904223 -0.403458
+ 5.38e+10Hz 0.903905 -0.404156
+ 5.39e+10Hz 0.903586 -0.404853
+ 5.4e+10Hz 0.903267 -0.40555
+ 5.41e+10Hz 0.902948 -0.406246
+ 5.42e+10Hz 0.902628 -0.406943
+ 5.43e+10Hz 0.902308 -0.407639
+ 5.44e+10Hz 0.901987 -0.408335
+ 5.45e+10Hz 0.901666 -0.409031
+ 5.46e+10Hz 0.901344 -0.409726
+ 5.47e+10Hz 0.901022 -0.410421
+ 5.48e+10Hz 0.9007 -0.411116
+ 5.49e+10Hz 0.900377 -0.411811
+ 5.5e+10Hz 0.900053 -0.412506
+ 5.51e+10Hz 0.899729 -0.4132
+ 5.52e+10Hz 0.899405 -0.413894
+ 5.53e+10Hz 0.89908 -0.414588
+ 5.54e+10Hz 0.898755 -0.415282
+ 5.55e+10Hz 0.898429 -0.415976
+ 5.56e+10Hz 0.898103 -0.416669
+ 5.57e+10Hz 0.897776 -0.417362
+ 5.58e+10Hz 0.897449 -0.418055
+ 5.59e+10Hz 0.897121 -0.418748
+ 5.6e+10Hz 0.896793 -0.41944
+ 5.61e+10Hz 0.896465 -0.420133
+ 5.62e+10Hz 0.896135 -0.420825
+ 5.63e+10Hz 0.895806 -0.421517
+ 5.64e+10Hz 0.895476 -0.422209
+ 5.65e+10Hz 0.895145 -0.4229
+ 5.66e+10Hz 0.894814 -0.423592
+ 5.67e+10Hz 0.894483 -0.424283
+ 5.68e+10Hz 0.894151 -0.424974
+ 5.69e+10Hz 0.893819 -0.425665
+ 5.7e+10Hz 0.893486 -0.426355
+ 5.71e+10Hz 0.893152 -0.427046
+ 5.72e+10Hz 0.892818 -0.427736
+ 5.73e+10Hz 0.892484 -0.428426
+ 5.74e+10Hz 0.892149 -0.429116
+ 5.75e+10Hz 0.891814 -0.429805
+ 5.76e+10Hz 0.891478 -0.430495
+ 5.77e+10Hz 0.891141 -0.431184
+ 5.78e+10Hz 0.890805 -0.431873
+ 5.79e+10Hz 0.890467 -0.432562
+ 5.8e+10Hz 0.890129 -0.433251
+ 5.81e+10Hz 0.889791 -0.433939
+ 5.82e+10Hz 0.889452 -0.434628
+ 5.83e+10Hz 0.889112 -0.435316
+ 5.84e+10Hz 0.888772 -0.436004
+ 5.85e+10Hz 0.888432 -0.436692
+ 5.86e+10Hz 0.888091 -0.43738
+ 5.87e+10Hz 0.887749 -0.438067
+ 5.88e+10Hz 0.887407 -0.438754
+ 5.89e+10Hz 0.887064 -0.439441
+ 5.9e+10Hz 0.886721 -0.440128
+ 5.91e+10Hz 0.886378 -0.440815
+ 5.92e+10Hz 0.886033 -0.441501
+ 5.93e+10Hz 0.885689 -0.442188
+ 5.94e+10Hz 0.885343 -0.442874
+ 5.95e+10Hz 0.884997 -0.44356
+ 5.96e+10Hz 0.884651 -0.444246
+ 5.97e+10Hz 0.884304 -0.444931
+ 5.98e+10Hz 0.883956 -0.445617
+ 5.99e+10Hz 0.883608 -0.446302
+ 6e+10Hz 0.88326 -0.446987
+ 6.01e+10Hz 0.882911 -0.447671
+ 6.02e+10Hz 0.882561 -0.448356
+ 6.03e+10Hz 0.88221 -0.44904
+ 6.04e+10Hz 0.88186 -0.449725
+ 6.05e+10Hz 0.881508 -0.450409
+ 6.06e+10Hz 0.881156 -0.451092
+ 6.07e+10Hz 0.880804 -0.451776
+ 6.08e+10Hz 0.88045 -0.452459
+ 6.09e+10Hz 0.880097 -0.453142
+ 6.1e+10Hz 0.879742 -0.453825
+ 6.11e+10Hz 0.879388 -0.454508
+ 6.12e+10Hz 0.879032 -0.45519
+ 6.13e+10Hz 0.878676 -0.455873
+ 6.14e+10Hz 0.87832 -0.456555
+ 6.15e+10Hz 0.877962 -0.457237
+ 6.16e+10Hz 0.877605 -0.457918
+ 6.17e+10Hz 0.877246 -0.458599
+ 6.18e+10Hz 0.876887 -0.459281
+ 6.19e+10Hz 0.876528 -0.459962
+ 6.2e+10Hz 0.876168 -0.460642
+ 6.21e+10Hz 0.875807 -0.461323
+ 6.22e+10Hz 0.875446 -0.462003
+ 6.23e+10Hz 0.875084 -0.462683
+ 6.24e+10Hz 0.874721 -0.463362
+ 6.25e+10Hz 0.874358 -0.464042
+ 6.26e+10Hz 0.873995 -0.464721
+ 6.27e+10Hz 0.87363 -0.4654
+ 6.28e+10Hz 0.873265 -0.466079
+ 6.29e+10Hz 0.8729 -0.466757
+ 6.3e+10Hz 0.872534 -0.467435
+ 6.31e+10Hz 0.872167 -0.468113
+ 6.32e+10Hz 0.8718 -0.468791
+ 6.33e+10Hz 0.871432 -0.469468
+ 6.34e+10Hz 0.871064 -0.470146
+ 6.35e+10Hz 0.870695 -0.470822
+ 6.36e+10Hz 0.870325 -0.471499
+ 6.37e+10Hz 0.869955 -0.472175
+ 6.38e+10Hz 0.869584 -0.472851
+ 6.39e+10Hz 0.869213 -0.473527
+ 6.4e+10Hz 0.868841 -0.474202
+ 6.41e+10Hz 0.868468 -0.474878
+ 6.42e+10Hz 0.868095 -0.475552
+ 6.43e+10Hz 0.867721 -0.476227
+ 6.44e+10Hz 0.867347 -0.476901
+ 6.45e+10Hz 0.866972 -0.477575
+ 6.46e+10Hz 0.866596 -0.478249
+ 6.47e+10Hz 0.86622 -0.478922
+ 6.48e+10Hz 0.865843 -0.479595
+ 6.49e+10Hz 0.865466 -0.480268
+ 6.5e+10Hz 0.865088 -0.480941
+ 6.51e+10Hz 0.864709 -0.481613
+ 6.52e+10Hz 0.86433 -0.482284
+ 6.53e+10Hz 0.863951 -0.482956
+ 6.54e+10Hz 0.86357 -0.483627
+ 6.55e+10Hz 0.863189 -0.484298
+ 6.56e+10Hz 0.862808 -0.484969
+ 6.57e+10Hz 0.862426 -0.485639
+ 6.58e+10Hz 0.862043 -0.486309
+ 6.59e+10Hz 0.86166 -0.486978
+ 6.6e+10Hz 0.861276 -0.487647
+ 6.61e+10Hz 0.860892 -0.488316
+ 6.62e+10Hz 0.860507 -0.488985
+ 6.63e+10Hz 0.860121 -0.489653
+ 6.64e+10Hz 0.859735 -0.490321
+ 6.65e+10Hz 0.859349 -0.490988
+ 6.66e+10Hz 0.858961 -0.491655
+ 6.67e+10Hz 0.858573 -0.492322
+ 6.68e+10Hz 0.858185 -0.492988
+ 6.69e+10Hz 0.857796 -0.493655
+ 6.7e+10Hz 0.857407 -0.49432
+ 6.71e+10Hz 0.857017 -0.494986
+ 6.72e+10Hz 0.856626 -0.495651
+ 6.73e+10Hz 0.856235 -0.496315
+ 6.74e+10Hz 0.855843 -0.49698
+ 6.75e+10Hz 0.855451 -0.497643
+ 6.76e+10Hz 0.855058 -0.498307
+ 6.77e+10Hz 0.854665 -0.49897
+ 6.78e+10Hz 0.854271 -0.499633
+ 6.79e+10Hz 0.853876 -0.500295
+ 6.8e+10Hz 0.853481 -0.500958
+ 6.81e+10Hz 0.853085 -0.501619
+ 6.82e+10Hz 0.852689 -0.502281
+ 6.83e+10Hz 0.852293 -0.502942
+ 6.84e+10Hz 0.851896 -0.503602
+ 6.85e+10Hz 0.851498 -0.504262
+ 6.86e+10Hz 0.8511 -0.504922
+ 6.87e+10Hz 0.850701 -0.505582
+ 6.88e+10Hz 0.850302 -0.506241
+ 6.89e+10Hz 0.849902 -0.506899
+ 6.9e+10Hz 0.849501 -0.507558
+ 6.91e+10Hz 0.849101 -0.508216
+ 6.92e+10Hz 0.848699 -0.508873
+ 6.93e+10Hz 0.848297 -0.509531
+ 6.94e+10Hz 0.847895 -0.510187
+ 6.95e+10Hz 0.847492 -0.510844
+ 6.96e+10Hz 0.847089 -0.5115
+ 6.97e+10Hz 0.846685 -0.512156
+ 6.98e+10Hz 0.84628 -0.512811
+ 6.99e+10Hz 0.845875 -0.513466
+ 7e+10Hz 0.84547 -0.51412
+ 7.01e+10Hz 0.845064 -0.514774
+ 7.02e+10Hz 0.844658 -0.515428
+ 7.03e+10Hz 0.844251 -0.516082
+ 7.04e+10Hz 0.843843 -0.516735
+ 7.05e+10Hz 0.843436 -0.517387
+ 7.06e+10Hz 0.843027 -0.518039
+ 7.07e+10Hz 0.842618 -0.518691
+ 7.08e+10Hz 0.842209 -0.519343
+ 7.09e+10Hz 0.841799 -0.519994
+ 7.1e+10Hz 0.841389 -0.520645
+ 7.11e+10Hz 0.840978 -0.521295
+ 7.12e+10Hz 0.840567 -0.521945
+ 7.13e+10Hz 0.840155 -0.522595
+ 7.14e+10Hz 0.839743 -0.523244
+ 7.15e+10Hz 0.839331 -0.523893
+ 7.16e+10Hz 0.838918 -0.524541
+ 7.17e+10Hz 0.838504 -0.525189
+ 7.18e+10Hz 0.83809 -0.525837
+ 7.19e+10Hz 0.837676 -0.526484
+ 7.2e+10Hz 0.837261 -0.527131
+ 7.21e+10Hz 0.836845 -0.527778
+ 7.22e+10Hz 0.836429 -0.528424
+ 7.23e+10Hz 0.836013 -0.52907
+ 7.24e+10Hz 0.835596 -0.529716
+ 7.25e+10Hz 0.835179 -0.530361
+ 7.26e+10Hz 0.834762 -0.531005
+ 7.27e+10Hz 0.834343 -0.53165
+ 7.28e+10Hz 0.833925 -0.532294
+ 7.29e+10Hz 0.833506 -0.532938
+ 7.3e+10Hz 0.833087 -0.533581
+ 7.31e+10Hz 0.832667 -0.534224
+ 7.32e+10Hz 0.832246 -0.534867
+ 7.33e+10Hz 0.831826 -0.535509
+ 7.34e+10Hz 0.831404 -0.536151
+ 7.35e+10Hz 0.830983 -0.536792
+ 7.36e+10Hz 0.830561 -0.537434
+ 7.37e+10Hz 0.830138 -0.538075
+ 7.38e+10Hz 0.829715 -0.538715
+ 7.39e+10Hz 0.829292 -0.539355
+ 7.4e+10Hz 0.828868 -0.539995
+ 7.41e+10Hz 0.828444 -0.540635
+ 7.42e+10Hz 0.828019 -0.541274
+ 7.43e+10Hz 0.827594 -0.541913
+ 7.44e+10Hz 0.827168 -0.542551
+ 7.45e+10Hz 0.826742 -0.543189
+ 7.46e+10Hz 0.826316 -0.543827
+ 7.47e+10Hz 0.825889 -0.544465
+ 7.48e+10Hz 0.825462 -0.545102
+ 7.49e+10Hz 0.825034 -0.545739
+ 7.5e+10Hz 0.824606 -0.546375
+ 7.51e+10Hz 0.824177 -0.547011
+ 7.52e+10Hz 0.823748 -0.547647
+ 7.53e+10Hz 0.823318 -0.548283
+ 7.54e+10Hz 0.822888 -0.548918
+ 7.55e+10Hz 0.822458 -0.549553
+ 7.56e+10Hz 0.822027 -0.550187
+ 7.57e+10Hz 0.821596 -0.550821
+ 7.58e+10Hz 0.821164 -0.551455
+ 7.59e+10Hz 0.820732 -0.552089
+ 7.6e+10Hz 0.8203 -0.552722
+ 7.61e+10Hz 0.819867 -0.553355
+ 7.62e+10Hz 0.819433 -0.553988
+ 7.63e+10Hz 0.819 -0.55462
+ 7.64e+10Hz 0.818565 -0.555252
+ 7.65e+10Hz 0.818131 -0.555884
+ 7.66e+10Hz 0.817695 -0.556515
+ 7.67e+10Hz 0.81726 -0.557146
+ 7.68e+10Hz 0.816824 -0.557777
+ 7.69e+10Hz 0.816387 -0.558408
+ 7.7e+10Hz 0.81595 -0.559038
+ 7.71e+10Hz 0.815513 -0.559668
+ 7.72e+10Hz 0.815075 -0.560297
+ 7.73e+10Hz 0.814637 -0.560926
+ 7.74e+10Hz 0.814198 -0.561555
+ 7.75e+10Hz 0.813759 -0.562184
+ 7.76e+10Hz 0.813319 -0.562812
+ 7.77e+10Hz 0.812879 -0.563441
+ 7.78e+10Hz 0.812439 -0.564068
+ 7.79e+10Hz 0.811998 -0.564696
+ 7.8e+10Hz 0.811556 -0.565323
+ 7.81e+10Hz 0.811114 -0.56595
+ 7.82e+10Hz 0.810672 -0.566576
+ 7.83e+10Hz 0.810229 -0.567203
+ 7.84e+10Hz 0.809786 -0.567829
+ 7.85e+10Hz 0.809342 -0.568454
+ 7.86e+10Hz 0.808898 -0.56908
+ 7.87e+10Hz 0.808453 -0.569705
+ 7.88e+10Hz 0.808008 -0.57033
+ 7.89e+10Hz 0.807563 -0.570954
+ 7.9e+10Hz 0.807117 -0.571579
+ 7.91e+10Hz 0.80667 -0.572202
+ 7.92e+10Hz 0.806223 -0.572826
+ 7.93e+10Hz 0.805776 -0.573449
+ 7.94e+10Hz 0.805328 -0.574072
+ 7.95e+10Hz 0.804879 -0.574695
+ 7.96e+10Hz 0.804431 -0.575318
+ 7.97e+10Hz 0.803981 -0.57594
+ 7.98e+10Hz 0.803531 -0.576562
+ 7.99e+10Hz 0.803081 -0.577183
+ 8e+10Hz 0.80263 -0.577805
+ 8.01e+10Hz 0.802179 -0.578426
+ 8.02e+10Hz 0.801727 -0.579046
+ 8.03e+10Hz 0.801275 -0.579667
+ 8.04e+10Hz 0.800822 -0.580287
+ 8.05e+10Hz 0.800369 -0.580907
+ 8.06e+10Hz 0.799915 -0.581526
+ 8.07e+10Hz 0.799461 -0.582145
+ 8.08e+10Hz 0.799006 -0.582764
+ 8.09e+10Hz 0.798551 -0.583383
+ 8.1e+10Hz 0.798095 -0.584001
+ 8.11e+10Hz 0.797639 -0.584619
+ 8.12e+10Hz 0.797182 -0.585237
+ 8.13e+10Hz 0.796725 -0.585854
+ 8.14e+10Hz 0.796267 -0.586471
+ 8.15e+10Hz 0.795809 -0.587088
+ 8.16e+10Hz 0.795351 -0.587704
+ 8.17e+10Hz 0.794891 -0.58832
+ 8.18e+10Hz 0.794432 -0.588936
+ 8.19e+10Hz 0.793971 -0.589552
+ 8.2e+10Hz 0.793511 -0.590167
+ 8.21e+10Hz 0.793049 -0.590782
+ 8.22e+10Hz 0.792588 -0.591396
+ 8.23e+10Hz 0.792125 -0.592011
+ 8.24e+10Hz 0.791663 -0.592625
+ 8.25e+10Hz 0.791199 -0.593238
+ 8.26e+10Hz 0.790736 -0.593852
+ 8.27e+10Hz 0.790271 -0.594464
+ 8.28e+10Hz 0.789806 -0.595077
+ 8.29e+10Hz 0.789341 -0.595689
+ 8.3e+10Hz 0.788875 -0.596301
+ 8.31e+10Hz 0.788409 -0.596913
+ 8.32e+10Hz 0.787942 -0.597524
+ 8.33e+10Hz 0.787475 -0.598135
+ 8.34e+10Hz 0.787007 -0.598746
+ 8.35e+10Hz 0.786538 -0.599356
+ 8.36e+10Hz 0.786069 -0.599966
+ 8.37e+10Hz 0.7856 -0.600576
+ 8.38e+10Hz 0.78513 -0.601185
+ 8.39e+10Hz 0.784659 -0.601794
+ 8.4e+10Hz 0.784188 -0.602403
+ 8.41e+10Hz 0.783716 -0.603011
+ 8.42e+10Hz 0.783244 -0.603619
+ 8.43e+10Hz 0.782772 -0.604226
+ 8.44e+10Hz 0.782299 -0.604833
+ 8.45e+10Hz 0.781825 -0.60544
+ 8.46e+10Hz 0.781351 -0.606047
+ 8.47e+10Hz 0.780876 -0.606653
+ 8.48e+10Hz 0.780401 -0.607259
+ 8.49e+10Hz 0.779925 -0.607864
+ 8.5e+10Hz 0.779449 -0.608469
+ 8.51e+10Hz 0.778972 -0.609074
+ 8.52e+10Hz 0.778495 -0.609678
+ 8.53e+10Hz 0.778017 -0.610282
+ 8.54e+10Hz 0.777539 -0.610885
+ 8.55e+10Hz 0.77706 -0.611488
+ 8.56e+10Hz 0.77658 -0.612091
+ 8.57e+10Hz 0.7761 -0.612693
+ 8.58e+10Hz 0.77562 -0.613295
+ 8.59e+10Hz 0.775139 -0.613897
+ 8.6e+10Hz 0.774657 -0.614498
+ 8.61e+10Hz 0.774176 -0.615099
+ 8.62e+10Hz 0.773693 -0.6157
+ 8.63e+10Hz 0.77321 -0.6163
+ 8.64e+10Hz 0.772726 -0.616899
+ 8.65e+10Hz 0.772242 -0.617499
+ 8.66e+10Hz 0.771758 -0.618098
+ 8.67e+10Hz 0.771273 -0.618696
+ 8.68e+10Hz 0.770787 -0.619294
+ 8.69e+10Hz 0.770301 -0.619892
+ 8.7e+10Hz 0.769815 -0.620489
+ 8.71e+10Hz 0.769327 -0.621086
+ 8.72e+10Hz 0.76884 -0.621682
+ 8.73e+10Hz 0.768352 -0.622278
+ 8.74e+10Hz 0.767863 -0.622874
+ 8.75e+10Hz 0.767374 -0.623469
+ 8.76e+10Hz 0.766884 -0.624064
+ 8.77e+10Hz 0.766394 -0.624659
+ 8.78e+10Hz 0.765904 -0.625253
+ 8.79e+10Hz 0.765413 -0.625846
+ 8.8e+10Hz 0.764921 -0.626439
+ 8.81e+10Hz 0.764429 -0.627032
+ 8.82e+10Hz 0.763936 -0.627624
+ 8.83e+10Hz 0.763443 -0.628216
+ 8.84e+10Hz 0.76295 -0.628808
+ 8.85e+10Hz 0.762456 -0.629399
+ 8.86e+10Hz 0.761961 -0.629989
+ 8.87e+10Hz 0.761466 -0.63058
+ 8.88e+10Hz 0.760971 -0.631169
+ 8.89e+10Hz 0.760475 -0.631759
+ 8.9e+10Hz 0.759978 -0.632348
+ 8.91e+10Hz 0.759481 -0.632936
+ 8.92e+10Hz 0.758984 -0.633524
+ 8.93e+10Hz 0.758486 -0.634112
+ 8.94e+10Hz 0.757987 -0.634699
+ 8.95e+10Hz 0.757489 -0.635286
+ 8.96e+10Hz 0.756989 -0.635872
+ 8.97e+10Hz 0.756489 -0.636458
+ 8.98e+10Hz 0.755989 -0.637043
+ 8.99e+10Hz 0.755489 -0.637628
+ 9e+10Hz 0.754987 -0.638213
+ 9.01e+10Hz 0.754486 -0.638797
+ 9.02e+10Hz 0.753984 -0.639381
+ 9.03e+10Hz 0.753481 -0.639964
+ 9.04e+10Hz 0.752978 -0.640547
+ 9.05e+10Hz 0.752475 -0.641129
+ 9.06e+10Hz 0.751971 -0.641711
+ 9.07e+10Hz 0.751466 -0.642292
+ 9.08e+10Hz 0.750961 -0.642873
+ 9.09e+10Hz 0.750456 -0.643454
+ 9.1e+10Hz 0.749951 -0.644034
+ 9.11e+10Hz 0.749444 -0.644614
+ 9.12e+10Hz 0.748938 -0.645193
+ 9.13e+10Hz 0.748431 -0.645772
+ 9.14e+10Hz 0.747923 -0.646351
+ 9.15e+10Hz 0.747415 -0.646928
+ 9.16e+10Hz 0.746907 -0.647506
+ 9.17e+10Hz 0.746398 -0.648083
+ 9.18e+10Hz 0.745889 -0.64866
+ 9.19e+10Hz 0.745379 -0.649236
+ 9.2e+10Hz 0.744869 -0.649812
+ 9.21e+10Hz 0.744359 -0.650387
+ 9.22e+10Hz 0.743848 -0.650962
+ 9.23e+10Hz 0.743337 -0.651536
+ 9.24e+10Hz 0.742825 -0.65211
+ 9.25e+10Hz 0.742313 -0.652684
+ 9.26e+10Hz 0.7418 -0.653257
+ 9.27e+10Hz 0.741287 -0.65383
+ 9.28e+10Hz 0.740774 -0.654402
+ 9.29e+10Hz 0.74026 -0.654974
+ 9.3e+10Hz 0.739745 -0.655545
+ 9.31e+10Hz 0.739231 -0.656116
+ 9.32e+10Hz 0.738716 -0.656687
+ 9.33e+10Hz 0.7382 -0.657257
+ 9.34e+10Hz 0.737684 -0.657827
+ 9.35e+10Hz 0.737168 -0.658396
+ 9.36e+10Hz 0.736651 -0.658965
+ 9.37e+10Hz 0.736134 -0.659533
+ 9.38e+10Hz 0.735617 -0.660101
+ 9.39e+10Hz 0.735099 -0.660668
+ 9.4e+10Hz 0.73458 -0.661235
+ 9.41e+10Hz 0.734062 -0.661802
+ 9.42e+10Hz 0.733542 -0.662368
+ 9.43e+10Hz 0.733023 -0.662934
+ 9.44e+10Hz 0.732503 -0.6635
+ 9.45e+10Hz 0.731983 -0.664065
+ 9.46e+10Hz 0.731462 -0.664629
+ 9.47e+10Hz 0.730941 -0.665193
+ 9.48e+10Hz 0.730419 -0.665757
+ 9.49e+10Hz 0.729897 -0.66632
+ 9.5e+10Hz 0.729375 -0.666883
+ 9.51e+10Hz 0.728852 -0.667446
+ 9.52e+10Hz 0.728329 -0.668008
+ 9.53e+10Hz 0.727806 -0.668569
+ 9.54e+10Hz 0.727282 -0.669131
+ 9.55e+10Hz 0.726758 -0.669691
+ 9.56e+10Hz 0.726233 -0.670252
+ 9.57e+10Hz 0.725708 -0.670812
+ 9.58e+10Hz 0.725182 -0.671371
+ 9.59e+10Hz 0.724657 -0.671931
+ 9.6e+10Hz 0.72413 -0.672489
+ 9.61e+10Hz 0.723604 -0.673048
+ 9.62e+10Hz 0.723077 -0.673606
+ 9.63e+10Hz 0.722549 -0.674163
+ 9.64e+10Hz 0.722022 -0.67472
+ 9.65e+10Hz 0.721493 -0.675277
+ 9.66e+10Hz 0.720965 -0.675833
+ 9.67e+10Hz 0.720436 -0.676389
+ 9.68e+10Hz 0.719906 -0.676945
+ 9.69e+10Hz 0.719377 -0.6775
+ 9.7e+10Hz 0.718847 -0.678055
+ 9.71e+10Hz 0.718316 -0.678609
+ 9.72e+10Hz 0.717785 -0.679163
+ 9.73e+10Hz 0.717254 -0.679717
+ 9.74e+10Hz 0.716722 -0.68027
+ 9.75e+10Hz 0.71619 -0.680823
+ 9.76e+10Hz 0.715658 -0.681375
+ 9.77e+10Hz 0.715125 -0.681927
+ 9.78e+10Hz 0.714591 -0.682479
+ 9.79e+10Hz 0.714058 -0.68303
+ 9.8e+10Hz 0.713524 -0.683581
+ 9.81e+10Hz 0.712989 -0.684132
+ 9.82e+10Hz 0.712454 -0.684682
+ 9.83e+10Hz 0.711919 -0.685231
+ 9.84e+10Hz 0.711383 -0.685781
+ 9.85e+10Hz 0.710847 -0.68633
+ 9.86e+10Hz 0.710311 -0.686878
+ 9.87e+10Hz 0.709774 -0.687426
+ 9.88e+10Hz 0.709237 -0.687974
+ 9.89e+10Hz 0.708699 -0.688521
+ 9.9e+10Hz 0.708161 -0.689068
+ 9.91e+10Hz 0.707623 -0.689615
+ 9.92e+10Hz 0.707084 -0.690161
+ 9.93e+10Hz 0.706545 -0.690707
+ 9.94e+10Hz 0.706005 -0.691253
+ 9.95e+10Hz 0.705465 -0.691798
+ 9.96e+10Hz 0.704924 -0.692343
+ 9.97e+10Hz 0.704383 -0.692887
+ 9.98e+10Hz 0.703842 -0.693431
+ 9.99e+10Hz 0.7033 -0.693975
+ 1e+11Hz 0.702758 -0.694518
+ 1.001e+11Hz 0.702216 -0.695061
+ 1.002e+11Hz 0.701673 -0.695603
+ 1.003e+11Hz 0.70113 -0.696145
+ 1.004e+11Hz 0.700586 -0.696687
+ 1.005e+11Hz 0.700042 -0.697228
+ 1.006e+11Hz 0.699497 -0.697769
+ 1.007e+11Hz 0.698952 -0.69831
+ 1.008e+11Hz 0.698407 -0.69885
+ 1.009e+11Hz 0.697861 -0.69939
+ 1.01e+11Hz 0.697314 -0.699929
+ 1.011e+11Hz 0.696768 -0.700468
+ 1.012e+11Hz 0.696221 -0.701007
+ 1.013e+11Hz 0.695673 -0.701545
+ 1.014e+11Hz 0.695125 -0.702083
+ 1.015e+11Hz 0.694577 -0.702621
+ 1.016e+11Hz 0.694028 -0.703158
+ 1.017e+11Hz 0.693479 -0.703694
+ 1.018e+11Hz 0.692929 -0.704231
+ 1.019e+11Hz 0.692379 -0.704767
+ 1.02e+11Hz 0.691828 -0.705302
+ 1.021e+11Hz 0.691277 -0.705838
+ 1.022e+11Hz 0.690726 -0.706373
+ 1.023e+11Hz 0.690174 -0.706907
+ 1.024e+11Hz 0.689622 -0.707441
+ 1.025e+11Hz 0.689069 -0.707975
+ 1.026e+11Hz 0.688516 -0.708508
+ 1.027e+11Hz 0.687962 -0.709041
+ 1.028e+11Hz 0.687408 -0.709573
+ 1.029e+11Hz 0.686854 -0.710106
+ 1.03e+11Hz 0.686299 -0.710637
+ 1.031e+11Hz 0.685743 -0.711169
+ 1.032e+11Hz 0.685188 -0.711699
+ 1.033e+11Hz 0.684631 -0.71223
+ 1.034e+11Hz 0.684075 -0.71276
+ 1.035e+11Hz 0.683518 -0.71329
+ 1.036e+11Hz 0.68296 -0.713819
+ 1.037e+11Hz 0.682402 -0.714348
+ 1.038e+11Hz 0.681844 -0.714877
+ 1.039e+11Hz 0.681285 -0.715405
+ 1.04e+11Hz 0.680725 -0.715932
+ 1.041e+11Hz 0.680165 -0.71646
+ 1.042e+11Hz 0.679605 -0.716987
+ 1.043e+11Hz 0.679044 -0.717513
+ 1.044e+11Hz 0.678483 -0.718039
+ 1.045e+11Hz 0.677922 -0.718565
+ 1.046e+11Hz 0.67736 -0.71909
+ 1.047e+11Hz 0.676797 -0.719615
+ 1.048e+11Hz 0.676234 -0.720139
+ 1.049e+11Hz 0.675671 -0.720663
+ 1.05e+11Hz 0.675107 -0.721187
+ 1.051e+11Hz 0.674543 -0.72171
+ 1.052e+11Hz 0.673978 -0.722233
+ 1.053e+11Hz 0.673413 -0.722755
+ 1.054e+11Hz 0.672847 -0.723277
+ 1.055e+11Hz 0.672281 -0.723799
+ 1.056e+11Hz 0.671714 -0.72432
+ 1.057e+11Hz 0.671147 -0.72484
+ 1.058e+11Hz 0.67058 -0.72536
+ 1.059e+11Hz 0.670012 -0.72588
+ 1.06e+11Hz 0.669444 -0.7264
+ 1.061e+11Hz 0.668875 -0.726918
+ 1.062e+11Hz 0.668305 -0.727437
+ 1.063e+11Hz 0.667736 -0.727955
+ 1.064e+11Hz 0.667166 -0.728472
+ 1.065e+11Hz 0.666595 -0.728989
+ 1.066e+11Hz 0.666024 -0.729506
+ 1.067e+11Hz 0.665452 -0.730022
+ 1.068e+11Hz 0.66488 -0.730538
+ 1.069e+11Hz 0.664308 -0.731053
+ 1.07e+11Hz 0.663735 -0.731568
+ 1.071e+11Hz 0.663162 -0.732083
+ 1.072e+11Hz 0.662588 -0.732597
+ 1.073e+11Hz 0.662014 -0.73311
+ 1.074e+11Hz 0.661439 -0.733623
+ 1.075e+11Hz 0.660864 -0.734136
+ 1.076e+11Hz 0.660288 -0.734648
+ 1.077e+11Hz 0.659712 -0.73516
+ 1.078e+11Hz 0.659136 -0.735671
+ 1.079e+11Hz 0.658559 -0.736182
+ 1.08e+11Hz 0.657982 -0.736692
+ 1.081e+11Hz 0.657404 -0.737202
+ 1.082e+11Hz 0.656826 -0.737711
+ 1.083e+11Hz 0.656247 -0.73822
+ 1.084e+11Hz 0.655668 -0.738728
+ 1.085e+11Hz 0.655088 -0.739236
+ 1.086e+11Hz 0.654508 -0.739744
+ 1.087e+11Hz 0.653928 -0.740251
+ 1.088e+11Hz 0.653347 -0.740757
+ 1.089e+11Hz 0.652766 -0.741263
+ 1.09e+11Hz 0.652184 -0.741769
+ 1.091e+11Hz 0.651602 -0.742274
+ 1.092e+11Hz 0.65102 -0.742778
+ 1.093e+11Hz 0.650437 -0.743282
+ 1.094e+11Hz 0.649853 -0.743786
+ 1.095e+11Hz 0.649269 -0.744289
+ 1.096e+11Hz 0.648685 -0.744792
+ 1.097e+11Hz 0.6481 -0.745294
+ 1.098e+11Hz 0.647515 -0.745796
+ 1.099e+11Hz 0.64693 -0.746297
+ 1.1e+11Hz 0.646344 -0.746797
+ 1.101e+11Hz 0.645757 -0.747298
+ 1.102e+11Hz 0.645171 -0.747797
+ 1.103e+11Hz 0.644583 -0.748297
+ 1.104e+11Hz 0.643996 -0.748795
+ 1.105e+11Hz 0.643408 -0.749293
+ 1.106e+11Hz 0.642819 -0.749791
+ 1.107e+11Hz 0.642231 -0.750288
+ 1.108e+11Hz 0.641641 -0.750785
+ 1.109e+11Hz 0.641052 -0.751281
+ 1.11e+11Hz 0.640462 -0.751777
+ 1.111e+11Hz 0.639871 -0.752272
+ 1.112e+11Hz 0.63928 -0.752767
+ 1.113e+11Hz 0.638689 -0.753261
+ 1.114e+11Hz 0.638097 -0.753755
+ 1.115e+11Hz 0.637505 -0.754248
+ 1.116e+11Hz 0.636913 -0.754741
+ 1.117e+11Hz 0.63632 -0.755233
+ 1.118e+11Hz 0.635727 -0.755725
+ 1.119e+11Hz 0.635133 -0.756216
+ 1.12e+11Hz 0.634539 -0.756707
+ 1.121e+11Hz 0.633944 -0.757197
+ 1.122e+11Hz 0.63335 -0.757687
+ 1.123e+11Hz 0.632754 -0.758176
+ 1.124e+11Hz 0.632159 -0.758665
+ 1.125e+11Hz 0.631563 -0.759153
+ 1.126e+11Hz 0.630966 -0.75964
+ 1.127e+11Hz 0.63037 -0.760128
+ 1.128e+11Hz 0.629773 -0.760614
+ 1.129e+11Hz 0.629175 -0.761101
+ 1.13e+11Hz 0.628577 -0.761586
+ 1.131e+11Hz 0.627979 -0.762071
+ 1.132e+11Hz 0.62738 -0.762556
+ 1.133e+11Hz 0.626781 -0.76304
+ 1.134e+11Hz 0.626182 -0.763524
+ 1.135e+11Hz 0.625582 -0.764007
+ 1.136e+11Hz 0.624982 -0.76449
+ 1.137e+11Hz 0.624382 -0.764972
+ 1.138e+11Hz 0.623781 -0.765453
+ 1.139e+11Hz 0.62318 -0.765935
+ 1.14e+11Hz 0.622578 -0.766415
+ 1.141e+11Hz 0.621976 -0.766895
+ 1.142e+11Hz 0.621374 -0.767375
+ 1.143e+11Hz 0.620771 -0.767854
+ 1.144e+11Hz 0.620168 -0.768333
+ 1.145e+11Hz 0.619565 -0.768811
+ 1.146e+11Hz 0.618961 -0.769288
+ 1.147e+11Hz 0.618357 -0.769766
+ 1.148e+11Hz 0.617753 -0.770242
+ 1.149e+11Hz 0.617148 -0.770718
+ 1.15e+11Hz 0.616543 -0.771194
+ 1.151e+11Hz 0.615938 -0.771669
+ 1.152e+11Hz 0.615332 -0.772144
+ 1.153e+11Hz 0.614726 -0.772618
+ 1.154e+11Hz 0.614119 -0.773091
+ 1.155e+11Hz 0.613512 -0.773565
+ 1.156e+11Hz 0.612905 -0.774037
+ 1.157e+11Hz 0.612298 -0.774509
+ 1.158e+11Hz 0.61169 -0.774981
+ 1.159e+11Hz 0.611081 -0.775452
+ 1.16e+11Hz 0.610473 -0.775923
+ 1.161e+11Hz 0.609864 -0.776393
+ 1.162e+11Hz 0.609255 -0.776863
+ 1.163e+11Hz 0.608645 -0.777332
+ 1.164e+11Hz 0.608035 -0.777801
+ 1.165e+11Hz 0.607425 -0.778269
+ 1.166e+11Hz 0.606814 -0.778737
+ 1.167e+11Hz 0.606203 -0.779204
+ 1.168e+11Hz 0.605592 -0.779671
+ 1.169e+11Hz 0.60498 -0.780137
+ 1.17e+11Hz 0.604368 -0.780603
+ 1.171e+11Hz 0.603756 -0.781068
+ 1.172e+11Hz 0.603144 -0.781533
+ 1.173e+11Hz 0.602531 -0.781997
+ 1.174e+11Hz 0.601917 -0.782461
+ 1.175e+11Hz 0.601304 -0.782925
+ 1.176e+11Hz 0.60069 -0.783388
+ 1.177e+11Hz 0.600075 -0.78385
+ 1.178e+11Hz 0.599461 -0.784312
+ 1.179e+11Hz 0.598846 -0.784774
+ 1.18e+11Hz 0.59823 -0.785235
+ 1.181e+11Hz 0.597615 -0.785695
+ 1.182e+11Hz 0.596999 -0.786155
+ 1.183e+11Hz 0.596382 -0.786615
+ 1.184e+11Hz 0.595766 -0.787074
+ 1.185e+11Hz 0.595149 -0.787533
+ 1.186e+11Hz 0.594531 -0.787991
+ 1.187e+11Hz 0.593914 -0.788448
+ 1.188e+11Hz 0.593296 -0.788906
+ 1.189e+11Hz 0.592677 -0.789362
+ 1.19e+11Hz 0.592059 -0.789819
+ 1.191e+11Hz 0.59144 -0.790274
+ 1.192e+11Hz 0.59082 -0.79073
+ 1.193e+11Hz 0.590201 -0.791185
+ 1.194e+11Hz 0.589581 -0.791639
+ 1.195e+11Hz 0.58896 -0.792093
+ 1.196e+11Hz 0.58834 -0.792547
+ 1.197e+11Hz 0.587719 -0.793
+ 1.198e+11Hz 0.587097 -0.793452
+ 1.199e+11Hz 0.586475 -0.793904
+ 1.2e+11Hz 0.585853 -0.794356
+ 1.201e+11Hz 0.585231 -0.794807
+ 1.202e+11Hz 0.584608 -0.795258
+ 1.203e+11Hz 0.583985 -0.795708
+ 1.204e+11Hz 0.583362 -0.796158
+ 1.205e+11Hz 0.582738 -0.796607
+ 1.206e+11Hz 0.582114 -0.797056
+ 1.207e+11Hz 0.58149 -0.797504
+ 1.208e+11Hz 0.580865 -0.797952
+ 1.209e+11Hz 0.58024 -0.798399
+ 1.21e+11Hz 0.579614 -0.798846
+ 1.211e+11Hz 0.578988 -0.799293
+ 1.212e+11Hz 0.578362 -0.799739
+ 1.213e+11Hz 0.577736 -0.800185
+ 1.214e+11Hz 0.577109 -0.80063
+ 1.215e+11Hz 0.576482 -0.801074
+ 1.216e+11Hz 0.575854 -0.801519
+ 1.217e+11Hz 0.575226 -0.801962
+ 1.218e+11Hz 0.574598 -0.802406
+ 1.219e+11Hz 0.573969 -0.802848
+ 1.22e+11Hz 0.57334 -0.803291
+ 1.221e+11Hz 0.572711 -0.803733
+ 1.222e+11Hz 0.572081 -0.804174
+ 1.223e+11Hz 0.571451 -0.804615
+ 1.224e+11Hz 0.570821 -0.805055
+ 1.225e+11Hz 0.57019 -0.805495
+ 1.226e+11Hz 0.569559 -0.805935
+ 1.227e+11Hz 0.568928 -0.806374
+ 1.228e+11Hz 0.568296 -0.806813
+ 1.229e+11Hz 0.567664 -0.807251
+ 1.23e+11Hz 0.567032 -0.807689
+ 1.231e+11Hz 0.566399 -0.808126
+ 1.232e+11Hz 0.565765 -0.808563
+ 1.233e+11Hz 0.565132 -0.808999
+ 1.234e+11Hz 0.564498 -0.809435
+ 1.235e+11Hz 0.563864 -0.80987
+ 1.236e+11Hz 0.563229 -0.810305
+ 1.237e+11Hz 0.562594 -0.810739
+ 1.238e+11Hz 0.561959 -0.811173
+ 1.239e+11Hz 0.561323 -0.811607
+ 1.24e+11Hz 0.560687 -0.81204
+ 1.241e+11Hz 0.56005 -0.812472
+ 1.242e+11Hz 0.559413 -0.812904
+ 1.243e+11Hz 0.558776 -0.813336
+ 1.244e+11Hz 0.558139 -0.813767
+ 1.245e+11Hz 0.557501 -0.814198
+ 1.246e+11Hz 0.556862 -0.814628
+ 1.247e+11Hz 0.556224 -0.815057
+ 1.248e+11Hz 0.555585 -0.815487
+ 1.249e+11Hz 0.554945 -0.815915
+ 1.25e+11Hz 0.554305 -0.816343
+ 1.251e+11Hz 0.553665 -0.816771
+ 1.252e+11Hz 0.553025 -0.817198
+ 1.253e+11Hz 0.552384 -0.817625
+ 1.254e+11Hz 0.551743 -0.818051
+ 1.255e+11Hz 0.551101 -0.818477
+ 1.256e+11Hz 0.550459 -0.818902
+ 1.257e+11Hz 0.549817 -0.819327
+ 1.258e+11Hz 0.549174 -0.819752
+ 1.259e+11Hz 0.548531 -0.820175
+ 1.26e+11Hz 0.547887 -0.820599
+ 1.261e+11Hz 0.547243 -0.821021
+ 1.262e+11Hz 0.546599 -0.821444
+ 1.263e+11Hz 0.545954 -0.821866
+ 1.264e+11Hz 0.54531 -0.822287
+ 1.265e+11Hz 0.544664 -0.822708
+ 1.266e+11Hz 0.544018 -0.823128
+ 1.267e+11Hz 0.543372 -0.823548
+ 1.268e+11Hz 0.542726 -0.823967
+ 1.269e+11Hz 0.542079 -0.824386
+ 1.27e+11Hz 0.541432 -0.824804
+ 1.271e+11Hz 0.540784 -0.825222
+ 1.272e+11Hz 0.540136 -0.825639
+ 1.273e+11Hz 0.539488 -0.826056
+ 1.274e+11Hz 0.538839 -0.826472
+ 1.275e+11Hz 0.53819 -0.826888
+ 1.276e+11Hz 0.537541 -0.827303
+ 1.277e+11Hz 0.536891 -0.827718
+ 1.278e+11Hz 0.536241 -0.828132
+ 1.279e+11Hz 0.53559 -0.828546
+ 1.28e+11Hz 0.534939 -0.828959
+ 1.281e+11Hz 0.534288 -0.829372
+ 1.282e+11Hz 0.533636 -0.829784
+ 1.283e+11Hz 0.532984 -0.830195
+ 1.284e+11Hz 0.532332 -0.830606
+ 1.285e+11Hz 0.531679 -0.831017
+ 1.286e+11Hz 0.531026 -0.831427
+ 1.287e+11Hz 0.530373 -0.831836
+ 1.288e+11Hz 0.529719 -0.832245
+ 1.289e+11Hz 0.529065 -0.832654
+ 1.29e+11Hz 0.52841 -0.833062
+ 1.291e+11Hz 0.527755 -0.833469
+ 1.292e+11Hz 0.5271 -0.833876
+ 1.293e+11Hz 0.526444 -0.834282
+ 1.294e+11Hz 0.525788 -0.834688
+ 1.295e+11Hz 0.525132 -0.835093
+ 1.296e+11Hz 0.524475 -0.835498
+ 1.297e+11Hz 0.523818 -0.835902
+ 1.298e+11Hz 0.52316 -0.836305
+ 1.299e+11Hz 0.522503 -0.836708
+ 1.3e+11Hz 0.521844 -0.837111
+ 1.301e+11Hz 0.521186 -0.837513
+ 1.302e+11Hz 0.520527 -0.837914
+ 1.303e+11Hz 0.519868 -0.838315
+ 1.304e+11Hz 0.519208 -0.838715
+ 1.305e+11Hz 0.518548 -0.839115
+ 1.306e+11Hz 0.517888 -0.839514
+ 1.307e+11Hz 0.517228 -0.839912
+ 1.308e+11Hz 0.516567 -0.84031
+ 1.309e+11Hz 0.515905 -0.840708
+ 1.31e+11Hz 0.515244 -0.841105
+ 1.311e+11Hz 0.514582 -0.841501
+ 1.312e+11Hz 0.513919 -0.841897
+ 1.313e+11Hz 0.513257 -0.842292
+ 1.314e+11Hz 0.512594 -0.842687
+ 1.315e+11Hz 0.51193 -0.843081
+ 1.316e+11Hz 0.511267 -0.843475
+ 1.317e+11Hz 0.510603 -0.843868
+ 1.318e+11Hz 0.509938 -0.84426
+ 1.319e+11Hz 0.509274 -0.844652
+ 1.32e+11Hz 0.508609 -0.845043
+ 1.321e+11Hz 0.507943 -0.845434
+ 1.322e+11Hz 0.507278 -0.845824
+ 1.323e+11Hz 0.506612 -0.846214
+ 1.324e+11Hz 0.505945 -0.846603
+ 1.325e+11Hz 0.505279 -0.846992
+ 1.326e+11Hz 0.504612 -0.847379
+ 1.327e+11Hz 0.503944 -0.847767
+ 1.328e+11Hz 0.503277 -0.848154
+ 1.329e+11Hz 0.502609 -0.84854
+ 1.33e+11Hz 0.501941 -0.848925
+ 1.331e+11Hz 0.501272 -0.84931
+ 1.332e+11Hz 0.500603 -0.849695
+ 1.333e+11Hz 0.499934 -0.850079
+ 1.334e+11Hz 0.499265 -0.850462
+ 1.335e+11Hz 0.498595 -0.850845
+ 1.336e+11Hz 0.497925 -0.851227
+ 1.337e+11Hz 0.497254 -0.851609
+ 1.338e+11Hz 0.496584 -0.85199
+ 1.339e+11Hz 0.495913 -0.85237
+ 1.34e+11Hz 0.495241 -0.85275
+ 1.341e+11Hz 0.49457 -0.85313
+ 1.342e+11Hz 0.493898 -0.853509
+ 1.343e+11Hz 0.493225 -0.853887
+ 1.344e+11Hz 0.492553 -0.854264
+ 1.345e+11Hz 0.49188 -0.854641
+ 1.346e+11Hz 0.491207 -0.855018
+ 1.347e+11Hz 0.490534 -0.855394
+ 1.348e+11Hz 0.48986 -0.855769
+ 1.349e+11Hz 0.489186 -0.856144
+ 1.35e+11Hz 0.488512 -0.856518
+ 1.351e+11Hz 0.487837 -0.856892
+ 1.352e+11Hz 0.487162 -0.857265
+ 1.353e+11Hz 0.486487 -0.857637
+ 1.354e+11Hz 0.485812 -0.858009
+ 1.355e+11Hz 0.485136 -0.858381
+ 1.356e+11Hz 0.48446 -0.858751
+ 1.357e+11Hz 0.483784 -0.859122
+ 1.358e+11Hz 0.483107 -0.859491
+ 1.359e+11Hz 0.48243 -0.85986
+ 1.36e+11Hz 0.481753 -0.860229
+ 1.361e+11Hz 0.481076 -0.860597
+ 1.362e+11Hz 0.480398 -0.860964
+ 1.363e+11Hz 0.47972 -0.861331
+ 1.364e+11Hz 0.479042 -0.861697
+ 1.365e+11Hz 0.478363 -0.862063
+ 1.366e+11Hz 0.477684 -0.862428
+ 1.367e+11Hz 0.477005 -0.862792
+ 1.368e+11Hz 0.476326 -0.863156
+ 1.369e+11Hz 0.475646 -0.86352
+ 1.37e+11Hz 0.474967 -0.863882
+ 1.371e+11Hz 0.474286 -0.864245
+ 1.372e+11Hz 0.473606 -0.864606
+ 1.373e+11Hz 0.472925 -0.864967
+ 1.374e+11Hz 0.472244 -0.865328
+ 1.375e+11Hz 0.471563 -0.865688
+ 1.376e+11Hz 0.470882 -0.866047
+ 1.377e+11Hz 0.4702 -0.866406
+ 1.378e+11Hz 0.469518 -0.866765
+ 1.379e+11Hz 0.468836 -0.867122
+ 1.38e+11Hz 0.468153 -0.867479
+ 1.381e+11Hz 0.46747 -0.867836
+ 1.382e+11Hz 0.466787 -0.868192
+ 1.383e+11Hz 0.466104 -0.868548
+ 1.384e+11Hz 0.46542 -0.868903
+ 1.385e+11Hz 0.464737 -0.869257
+ 1.386e+11Hz 0.464053 -0.869611
+ 1.387e+11Hz 0.463368 -0.869964
+ 1.388e+11Hz 0.462684 -0.870317
+ 1.389e+11Hz 0.461999 -0.870669
+ 1.39e+11Hz 0.461314 -0.871021
+ 1.391e+11Hz 0.460628 -0.871372
+ 1.392e+11Hz 0.459942 -0.871722
+ 1.393e+11Hz 0.459257 -0.872072
+ 1.394e+11Hz 0.45857 -0.872422
+ 1.395e+11Hz 0.457884 -0.87277
+ 1.396e+11Hz 0.457197 -0.873119
+ 1.397e+11Hz 0.45651 -0.873466
+ 1.398e+11Hz 0.455823 -0.873814
+ 1.399e+11Hz 0.455136 -0.87416
+ 1.4e+11Hz 0.454448 -0.874506
+ 1.401e+11Hz 0.45376 -0.874852
+ 1.402e+11Hz 0.453072 -0.875197
+ 1.403e+11Hz 0.452383 -0.875541
+ 1.404e+11Hz 0.451694 -0.875885
+ 1.405e+11Hz 0.451005 -0.876229
+ 1.406e+11Hz 0.450316 -0.876571
+ 1.407e+11Hz 0.449627 -0.876914
+ 1.408e+11Hz 0.448937 -0.877255
+ 1.409e+11Hz 0.448247 -0.877597
+ 1.41e+11Hz 0.447556 -0.877937
+ 1.411e+11Hz 0.446866 -0.878277
+ 1.412e+11Hz 0.446175 -0.878617
+ 1.413e+11Hz 0.445484 -0.878956
+ 1.414e+11Hz 0.444793 -0.879294
+ 1.415e+11Hz 0.444101 -0.879632
+ 1.416e+11Hz 0.443409 -0.879969
+ 1.417e+11Hz 0.442717 -0.880306
+ 1.418e+11Hz 0.442025 -0.880642
+ 1.419e+11Hz 0.441332 -0.880978
+ 1.42e+11Hz 0.440639 -0.881313
+ 1.421e+11Hz 0.439946 -0.881648
+ 1.422e+11Hz 0.439252 -0.881982
+ 1.423e+11Hz 0.438559 -0.882316
+ 1.424e+11Hz 0.437865 -0.882649
+ 1.425e+11Hz 0.437171 -0.882981
+ 1.426e+11Hz 0.436476 -0.883313
+ 1.427e+11Hz 0.435781 -0.883644
+ 1.428e+11Hz 0.435086 -0.883975
+ 1.429e+11Hz 0.434391 -0.884305
+ 1.43e+11Hz 0.433695 -0.884635
+ 1.431e+11Hz 0.433 -0.884964
+ 1.432e+11Hz 0.432304 -0.885293
+ 1.433e+11Hz 0.431607 -0.885621
+ 1.434e+11Hz 0.430911 -0.885948
+ 1.435e+11Hz 0.430214 -0.886275
+ 1.436e+11Hz 0.429517 -0.886602
+ 1.437e+11Hz 0.428819 -0.886927
+ 1.438e+11Hz 0.428121 -0.887253
+ 1.439e+11Hz 0.427423 -0.887578
+ 1.44e+11Hz 0.426725 -0.887902
+ 1.441e+11Hz 0.426027 -0.888225
+ 1.442e+11Hz 0.425328 -0.888548
+ 1.443e+11Hz 0.424629 -0.888871
+ 1.444e+11Hz 0.42393 -0.889193
+ 1.445e+11Hz 0.42323 -0.889514
+ 1.446e+11Hz 0.42253 -0.889835
+ 1.447e+11Hz 0.42183 -0.890156
+ 1.448e+11Hz 0.42113 -0.890476
+ 1.449e+11Hz 0.420429 -0.890795
+ 1.45e+11Hz 0.419728 -0.891113
+ 1.451e+11Hz 0.419027 -0.891432
+ 1.452e+11Hz 0.418325 -0.891749
+ 1.453e+11Hz 0.417623 -0.892066
+ 1.454e+11Hz 0.416921 -0.892382
+ 1.455e+11Hz 0.416219 -0.892698
+ 1.456e+11Hz 0.415517 -0.893014
+ 1.457e+11Hz 0.414814 -0.893328
+ 1.458e+11Hz 0.41411 -0.893643
+ 1.459e+11Hz 0.413407 -0.893956
+ 1.46e+11Hz 0.412703 -0.894269
+ 1.461e+11Hz 0.411999 -0.894582
+ 1.462e+11Hz 0.411295 -0.894894
+ 1.463e+11Hz 0.410591 -0.895205
+ 1.464e+11Hz 0.409886 -0.895516
+ 1.465e+11Hz 0.409181 -0.895826
+ 1.466e+11Hz 0.408475 -0.896136
+ 1.467e+11Hz 0.40777 -0.896445
+ 1.468e+11Hz 0.407064 -0.896753
+ 1.469e+11Hz 0.406358 -0.897061
+ 1.47e+11Hz 0.405651 -0.897368
+ 1.471e+11Hz 0.404944 -0.897675
+ 1.472e+11Hz 0.404237 -0.897981
+ 1.473e+11Hz 0.40353 -0.898287
+ 1.474e+11Hz 0.402823 -0.898592
+ 1.475e+11Hz 0.402115 -0.898896
+ 1.476e+11Hz 0.401407 -0.8992
+ 1.477e+11Hz 0.400698 -0.899503
+ 1.478e+11Hz 0.39999 -0.899806
+ 1.479e+11Hz 0.399281 -0.900108
+ 1.48e+11Hz 0.398572 -0.900409
+ 1.481e+11Hz 0.397862 -0.90071
+ 1.482e+11Hz 0.397152 -0.90101
+ 1.483e+11Hz 0.396442 -0.90131
+ 1.484e+11Hz 0.395732 -0.901609
+ 1.485e+11Hz 0.395021 -0.901908
+ 1.486e+11Hz 0.394311 -0.902205
+ 1.487e+11Hz 0.393599 -0.902503
+ 1.488e+11Hz 0.392888 -0.902799
+ 1.489e+11Hz 0.392176 -0.903095
+ 1.49e+11Hz 0.391465 -0.903391
+ 1.491e+11Hz 0.390752 -0.903686
+ 1.492e+11Hz 0.39004 -0.90398
+ 1.493e+11Hz 0.389327 -0.904274
+ 1.494e+11Hz 0.388614 -0.904567
+ 1.495e+11Hz 0.387901 -0.904859
+ 1.496e+11Hz 0.387187 -0.905151
+ 1.497e+11Hz 0.386474 -0.905442
+ 1.498e+11Hz 0.38576 -0.905733
+ 1.499e+11Hz 0.385045 -0.906023
+ 1.5e+11Hz 0.384331 -0.906312
+ 1.501e+11Hz 0.383616 -0.906601
+ 1.502e+11Hz 0.382901 -0.906889
+ 1.503e+11Hz 0.382186 -0.907176
+ 1.504e+11Hz 0.38147 -0.907463
+ 1.505e+11Hz 0.380754 -0.907749
+ 1.506e+11Hz 0.380038 -0.908035
+ 1.507e+11Hz 0.379322 -0.90832
+ 1.508e+11Hz 0.378605 -0.908604
+ 1.509e+11Hz 0.377888 -0.908888
+ 1.51e+11Hz 0.377171 -0.909171
+ 1.511e+11Hz 0.376454 -0.909453
+ 1.512e+11Hz 0.375736 -0.909735
+ 1.513e+11Hz 0.375018 -0.910016
+ 1.514e+11Hz 0.3743 -0.910297
+ 1.515e+11Hz 0.373582 -0.910577
+ 1.516e+11Hz 0.372863 -0.910856
+ 1.517e+11Hz 0.372145 -0.911135
+ 1.518e+11Hz 0.371426 -0.911413
+ 1.519e+11Hz 0.370706 -0.91169
+ 1.52e+11Hz 0.369987 -0.911967
+ 1.521e+11Hz 0.369267 -0.912243
+ 1.522e+11Hz 0.368547 -0.912518
+ 1.523e+11Hz 0.367827 -0.912793
+ 1.524e+11Hz 0.367107 -0.913067
+ 1.525e+11Hz 0.366386 -0.91334
+ 1.526e+11Hz 0.365665 -0.913613
+ 1.527e+11Hz 0.364944 -0.913885
+ 1.528e+11Hz 0.364223 -0.914157
+ 1.529e+11Hz 0.363501 -0.914428
+ 1.53e+11Hz 0.362779 -0.914698
+ 1.531e+11Hz 0.362057 -0.914967
+ 1.532e+11Hz 0.361335 -0.915236
+ 1.533e+11Hz 0.360613 -0.915504
+ 1.534e+11Hz 0.35989 -0.915772
+ 1.535e+11Hz 0.359167 -0.916039
+ 1.536e+11Hz 0.358444 -0.916305
+ 1.537e+11Hz 0.357721 -0.916571
+ 1.538e+11Hz 0.356997 -0.916836
+ 1.539e+11Hz 0.356274 -0.9171
+ 1.54e+11Hz 0.35555 -0.917364
+ 1.541e+11Hz 0.354826 -0.917627
+ 1.542e+11Hz 0.354102 -0.917889
+ 1.543e+11Hz 0.353377 -0.91815
+ 1.544e+11Hz 0.352652 -0.918411
+ 1.545e+11Hz 0.351928 -0.918672
+ 1.546e+11Hz 0.351203 -0.918931
+ 1.547e+11Hz 0.350477 -0.91919
+ 1.548e+11Hz 0.349752 -0.919449
+ 1.549e+11Hz 0.349026 -0.919706
+ 1.55e+11Hz 0.348301 -0.919963
+ 1.551e+11Hz 0.347575 -0.92022
+ 1.552e+11Hz 0.346849 -0.920475
+ 1.553e+11Hz 0.346122 -0.920731
+ 1.554e+11Hz 0.345396 -0.920985
+ 1.555e+11Hz 0.344669 -0.921239
+ 1.556e+11Hz 0.343942 -0.921492
+ 1.557e+11Hz 0.343215 -0.921744
+ 1.558e+11Hz 0.342488 -0.921996
+ 1.559e+11Hz 0.341761 -0.922247
+ 1.56e+11Hz 0.341033 -0.922497
+ 1.561e+11Hz 0.340306 -0.922747
+ 1.562e+11Hz 0.339578 -0.922996
+ 1.563e+11Hz 0.33885 -0.923244
+ 1.564e+11Hz 0.338122 -0.923492
+ 1.565e+11Hz 0.337393 -0.923739
+ 1.566e+11Hz 0.336665 -0.923985
+ 1.567e+11Hz 0.335936 -0.924231
+ 1.568e+11Hz 0.335207 -0.924476
+ 1.569e+11Hz 0.334479 -0.924721
+ 1.57e+11Hz 0.33375 -0.924964
+ 1.571e+11Hz 0.33302 -0.925207
+ 1.572e+11Hz 0.332291 -0.92545
+ 1.573e+11Hz 0.331561 -0.925692
+ 1.574e+11Hz 0.330832 -0.925933
+ 1.575e+11Hz 0.330102 -0.926173
+ 1.576e+11Hz 0.329372 -0.926413
+ 1.577e+11Hz 0.328642 -0.926652
+ 1.578e+11Hz 0.327912 -0.92689
+ 1.579e+11Hz 0.327182 -0.927128
+ 1.58e+11Hz 0.326451 -0.927365
+ 1.581e+11Hz 0.325721 -0.927602
+ 1.582e+11Hz 0.32499 -0.927838
+ 1.583e+11Hz 0.324259 -0.928073
+ 1.584e+11Hz 0.323528 -0.928307
+ 1.585e+11Hz 0.322797 -0.928541
+ 1.586e+11Hz 0.322066 -0.928774
+ 1.587e+11Hz 0.321335 -0.929007
+ 1.588e+11Hz 0.320603 -0.929239
+ 1.589e+11Hz 0.319872 -0.92947
+ 1.59e+11Hz 0.31914 -0.929701
+ 1.591e+11Hz 0.318408 -0.929931
+ 1.592e+11Hz 0.317676 -0.93016
+ 1.593e+11Hz 0.316944 -0.930389
+ 1.594e+11Hz 0.316212 -0.930617
+ 1.595e+11Hz 0.31548 -0.930844
+ 1.596e+11Hz 0.314747 -0.931071
+ 1.597e+11Hz 0.314015 -0.931297
+ 1.598e+11Hz 0.313282 -0.931522
+ 1.599e+11Hz 0.31255 -0.931747
+ 1.6e+11Hz 0.311817 -0.931971
+ 1.601e+11Hz 0.311084 -0.932194
+ 1.602e+11Hz 0.310351 -0.932417
+ 1.603e+11Hz 0.309618 -0.932639
+ 1.604e+11Hz 0.308885 -0.932861
+ 1.605e+11Hz 0.308152 -0.933082
+ 1.606e+11Hz 0.307418 -0.933302
+ 1.607e+11Hz 0.306685 -0.933522
+ 1.608e+11Hz 0.305951 -0.933741
+ 1.609e+11Hz 0.305217 -0.933959
+ 1.61e+11Hz 0.304484 -0.934177
+ 1.611e+11Hz 0.30375 -0.934394
+ 1.612e+11Hz 0.303016 -0.93461
+ 1.613e+11Hz 0.302282 -0.934826
+ 1.614e+11Hz 0.301548 -0.935041
+ 1.615e+11Hz 0.300813 -0.935256
+ 1.616e+11Hz 0.300079 -0.935469
+ 1.617e+11Hz 0.299345 -0.935683
+ 1.618e+11Hz 0.29861 -0.935895
+ 1.619e+11Hz 0.297876 -0.936107
+ 1.62e+11Hz 0.297141 -0.936319
+ 1.621e+11Hz 0.296406 -0.936529
+ 1.622e+11Hz 0.295671 -0.936739
+ 1.623e+11Hz 0.294937 -0.936949
+ 1.624e+11Hz 0.294202 -0.937158
+ 1.625e+11Hz 0.293466 -0.937366
+ 1.626e+11Hz 0.292731 -0.937574
+ 1.627e+11Hz 0.291996 -0.93778
+ 1.628e+11Hz 0.291261 -0.937987
+ 1.629e+11Hz 0.290525 -0.938193
+ 1.63e+11Hz 0.28979 -0.938398
+ 1.631e+11Hz 0.289054 -0.938602
+ 1.632e+11Hz 0.288319 -0.938806
+ 1.633e+11Hz 0.287583 -0.939009
+ 1.634e+11Hz 0.286847 -0.939212
+ 1.635e+11Hz 0.286111 -0.939414
+ 1.636e+11Hz 0.285375 -0.939615
+ 1.637e+11Hz 0.284639 -0.939816
+ 1.638e+11Hz 0.283903 -0.940016
+ 1.639e+11Hz 0.283167 -0.940215
+ 1.64e+11Hz 0.282431 -0.940414
+ 1.641e+11Hz 0.281694 -0.940612
+ 1.642e+11Hz 0.280958 -0.94081
+ 1.643e+11Hz 0.280221 -0.941007
+ 1.644e+11Hz 0.279485 -0.941203
+ 1.645e+11Hz 0.278748 -0.941399
+ 1.646e+11Hz 0.278012 -0.941594
+ 1.647e+11Hz 0.277275 -0.941789
+ 1.648e+11Hz 0.276538 -0.941983
+ 1.649e+11Hz 0.275801 -0.942176
+ 1.65e+11Hz 0.275064 -0.942369
+ 1.651e+11Hz 0.274327 -0.942561
+ 1.652e+11Hz 0.27359 -0.942752
+ 1.653e+11Hz 0.272853 -0.942943
+ 1.654e+11Hz 0.272116 -0.943133
+ 1.655e+11Hz 0.271378 -0.943323
+ 1.656e+11Hz 0.270641 -0.943512
+ 1.657e+11Hz 0.269903 -0.9437
+ 1.658e+11Hz 0.269166 -0.943888
+ 1.659e+11Hz 0.268428 -0.944075
+ 1.66e+11Hz 0.267691 -0.944262
+ 1.661e+11Hz 0.266953 -0.944448
+ 1.662e+11Hz 0.266215 -0.944633
+ 1.663e+11Hz 0.265478 -0.944818
+ 1.664e+11Hz 0.26474 -0.945002
+ 1.665e+11Hz 0.264002 -0.945185
+ 1.666e+11Hz 0.263264 -0.945368
+ 1.667e+11Hz 0.262526 -0.945551
+ 1.668e+11Hz 0.261788 -0.945732
+ 1.669e+11Hz 0.261049 -0.945913
+ 1.67e+11Hz 0.260311 -0.946094
+ 1.671e+11Hz 0.259573 -0.946273
+ 1.672e+11Hz 0.258834 -0.946453
+ 1.673e+11Hz 0.258096 -0.946631
+ 1.674e+11Hz 0.257358 -0.946809
+ 1.675e+11Hz 0.256619 -0.946987
+ 1.676e+11Hz 0.255881 -0.947163
+ 1.677e+11Hz 0.255142 -0.94734
+ 1.678e+11Hz 0.254403 -0.947515
+ 1.679e+11Hz 0.253665 -0.94769
+ 1.68e+11Hz 0.252926 -0.947864
+ 1.681e+11Hz 0.252187 -0.948038
+ 1.682e+11Hz 0.251448 -0.948211
+ 1.683e+11Hz 0.250709 -0.948384
+ 1.684e+11Hz 0.24997 -0.948556
+ 1.685e+11Hz 0.249231 -0.948727
+ 1.686e+11Hz 0.248492 -0.948898
+ 1.687e+11Hz 0.247753 -0.949068
+ 1.688e+11Hz 0.247014 -0.949237
+ 1.689e+11Hz 0.246275 -0.949406
+ 1.69e+11Hz 0.245535 -0.949574
+ 1.691e+11Hz 0.244796 -0.949742
+ 1.692e+11Hz 0.244057 -0.949909
+ 1.693e+11Hz 0.243317 -0.950075
+ 1.694e+11Hz 0.242578 -0.950241
+ 1.695e+11Hz 0.241839 -0.950406
+ 1.696e+11Hz 0.241099 -0.950571
+ 1.697e+11Hz 0.24036 -0.950735
+ 1.698e+11Hz 0.23962 -0.950898
+ 1.699e+11Hz 0.23888 -0.951061
+ 1.7e+11Hz 0.238141 -0.951223
+ 1.701e+11Hz 0.237401 -0.951384
+ 1.702e+11Hz 0.236662 -0.951545
+ 1.703e+11Hz 0.235922 -0.951706
+ 1.704e+11Hz 0.235182 -0.951865
+ 1.705e+11Hz 0.234442 -0.952024
+ 1.706e+11Hz 0.233703 -0.952183
+ 1.707e+11Hz 0.232963 -0.952341
+ 1.708e+11Hz 0.232223 -0.952498
+ 1.709e+11Hz 0.231483 -0.952655
+ 1.71e+11Hz 0.230743 -0.952811
+ 1.711e+11Hz 0.230003 -0.952966
+ 1.712e+11Hz 0.229263 -0.953121
+ 1.713e+11Hz 0.228523 -0.953275
+ 1.714e+11Hz 0.227783 -0.953429
+ 1.715e+11Hz 0.227043 -0.953582
+ 1.716e+11Hz 0.226303 -0.953735
+ 1.717e+11Hz 0.225563 -0.953886
+ 1.718e+11Hz 0.224823 -0.954038
+ 1.719e+11Hz 0.224083 -0.954188
+ 1.72e+11Hz 0.223343 -0.954338
+ 1.721e+11Hz 0.222603 -0.954488
+ 1.722e+11Hz 0.221863 -0.954637
+ 1.723e+11Hz 0.221123 -0.954785
+ 1.724e+11Hz 0.220383 -0.954933
+ 1.725e+11Hz 0.219643 -0.95508
+ 1.726e+11Hz 0.218903 -0.955226
+ 1.727e+11Hz 0.218163 -0.955372
+ 1.728e+11Hz 0.217423 -0.955517
+ 1.729e+11Hz 0.216683 -0.955662
+ 1.73e+11Hz 0.215943 -0.955806
+ 1.731e+11Hz 0.215203 -0.955949
+ 1.732e+11Hz 0.214463 -0.956092
+ 1.733e+11Hz 0.213723 -0.956234
+ 1.734e+11Hz 0.212983 -0.956376
+ 1.735e+11Hz 0.212243 -0.956517
+ 1.736e+11Hz 0.211503 -0.956658
+ 1.737e+11Hz 0.210763 -0.956798
+ 1.738e+11Hz 0.210023 -0.956937
+ 1.739e+11Hz 0.209283 -0.957076
+ 1.74e+11Hz 0.208543 -0.957214
+ 1.741e+11Hz 0.207803 -0.957352
+ 1.742e+11Hz 0.207063 -0.957489
+ 1.743e+11Hz 0.206323 -0.957625
+ 1.744e+11Hz 0.205583 -0.957761
+ 1.745e+11Hz 0.204844 -0.957896
+ 1.746e+11Hz 0.204104 -0.958031
+ 1.747e+11Hz 0.203364 -0.958165
+ 1.748e+11Hz 0.202624 -0.958298
+ 1.749e+11Hz 0.201884 -0.958431
+ 1.75e+11Hz 0.201145 -0.958564
+ 1.751e+11Hz 0.200405 -0.958696
+ 1.752e+11Hz 0.199665 -0.958827
+ 1.753e+11Hz 0.198926 -0.958957
+ 1.754e+11Hz 0.198186 -0.959088
+ 1.755e+11Hz 0.197447 -0.959217
+ 1.756e+11Hz 0.196707 -0.959346
+ 1.757e+11Hz 0.195968 -0.959474
+ 1.758e+11Hz 0.195228 -0.959602
+ 1.759e+11Hz 0.194489 -0.95973
+ 1.76e+11Hz 0.19375 -0.959856
+ 1.761e+11Hz 0.19301 -0.959983
+ 1.762e+11Hz 0.192271 -0.960108
+ 1.763e+11Hz 0.191532 -0.960233
+ 1.764e+11Hz 0.190792 -0.960358
+ 1.765e+11Hz 0.190053 -0.960482
+ 1.766e+11Hz 0.189314 -0.960605
+ 1.767e+11Hz 0.188575 -0.960728
+ 1.768e+11Hz 0.187836 -0.96085
+ 1.769e+11Hz 0.187097 -0.960972
+ 1.77e+11Hz 0.186358 -0.961093
+ 1.771e+11Hz 0.185619 -0.961214
+ 1.772e+11Hz 0.18488 -0.961334
+ 1.773e+11Hz 0.184142 -0.961454
+ 1.774e+11Hz 0.183403 -0.961573
+ 1.775e+11Hz 0.182664 -0.961692
+ 1.776e+11Hz 0.181926 -0.96181
+ 1.777e+11Hz 0.181187 -0.961927
+ 1.778e+11Hz 0.180448 -0.962044
+ 1.779e+11Hz 0.17971 -0.962161
+ 1.78e+11Hz 0.178971 -0.962277
+ 1.781e+11Hz 0.178233 -0.962392
+ 1.782e+11Hz 0.177495 -0.962507
+ 1.783e+11Hz 0.176756 -0.962622
+ 1.784e+11Hz 0.176018 -0.962735
+ 1.785e+11Hz 0.17528 -0.962849
+ 1.786e+11Hz 0.174542 -0.962962
+ 1.787e+11Hz 0.173804 -0.963074
+ 1.788e+11Hz 0.173066 -0.963186
+ 1.789e+11Hz 0.172328 -0.963297
+ 1.79e+11Hz 0.17159 -0.963408
+ 1.791e+11Hz 0.170852 -0.963518
+ 1.792e+11Hz 0.170114 -0.963628
+ 1.793e+11Hz 0.169376 -0.963738
+ 1.794e+11Hz 0.168638 -0.963847
+ 1.795e+11Hz 0.167901 -0.963955
+ 1.796e+11Hz 0.167163 -0.964063
+ 1.797e+11Hz 0.166425 -0.96417
+ 1.798e+11Hz 0.165688 -0.964277
+ 1.799e+11Hz 0.16495 -0.964384
+ 1.8e+11Hz 0.164213 -0.96449
+ 1.801e+11Hz 0.163475 -0.964595
+ 1.802e+11Hz 0.162738 -0.9647
+ 1.803e+11Hz 0.162001 -0.964805
+ 1.804e+11Hz 0.161263 -0.964909
+ 1.805e+11Hz 0.160526 -0.965012
+ 1.806e+11Hz 0.159789 -0.965115
+ 1.807e+11Hz 0.159052 -0.965218
+ 1.808e+11Hz 0.158314 -0.96532
+ 1.809e+11Hz 0.157577 -0.965422
+ 1.81e+11Hz 0.15684 -0.965523
+ 1.811e+11Hz 0.156103 -0.965624
+ 1.812e+11Hz 0.155366 -0.965724
+ 1.813e+11Hz 0.154629 -0.965824
+ 1.814e+11Hz 0.153892 -0.965923
+ 1.815e+11Hz 0.153155 -0.966022
+ 1.816e+11Hz 0.152418 -0.966121
+ 1.817e+11Hz 0.151682 -0.966219
+ 1.818e+11Hz 0.150945 -0.966317
+ 1.819e+11Hz 0.150208 -0.966414
+ 1.82e+11Hz 0.149471 -0.96651
+ 1.821e+11Hz 0.148734 -0.966607
+ 1.822e+11Hz 0.147998 -0.966703
+ 1.823e+11Hz 0.147261 -0.966798
+ 1.824e+11Hz 0.146524 -0.966893
+ 1.825e+11Hz 0.145787 -0.966987
+ 1.826e+11Hz 0.145051 -0.967081
+ 1.827e+11Hz 0.144314 -0.967175
+ 1.828e+11Hz 0.143577 -0.967268
+ 1.829e+11Hz 0.142841 -0.967361
+ 1.83e+11Hz 0.142104 -0.967453
+ 1.831e+11Hz 0.141367 -0.967545
+ 1.832e+11Hz 0.140631 -0.967637
+ 1.833e+11Hz 0.139894 -0.967728
+ 1.834e+11Hz 0.139158 -0.967818
+ 1.835e+11Hz 0.138421 -0.967908
+ 1.836e+11Hz 0.137684 -0.967998
+ 1.837e+11Hz 0.136948 -0.968088
+ 1.838e+11Hz 0.136211 -0.968176
+ 1.839e+11Hz 0.135474 -0.968265
+ 1.84e+11Hz 0.134738 -0.968353
+ 1.841e+11Hz 0.134001 -0.968441
+ 1.842e+11Hz 0.133264 -0.968528
+ 1.843e+11Hz 0.132527 -0.968615
+ 1.844e+11Hz 0.131791 -0.968701
+ 1.845e+11Hz 0.131054 -0.968787
+ 1.846e+11Hz 0.130317 -0.968872
+ 1.847e+11Hz 0.12958 -0.968957
+ 1.848e+11Hz 0.128843 -0.969042
+ 1.849e+11Hz 0.128106 -0.969126
+ 1.85e+11Hz 0.127369 -0.96921
+ 1.851e+11Hz 0.126632 -0.969293
+ 1.852e+11Hz 0.125895 -0.969376
+ 1.853e+11Hz 0.125158 -0.969459
+ 1.854e+11Hz 0.124421 -0.969541
+ 1.855e+11Hz 0.123684 -0.969623
+ 1.856e+11Hz 0.122947 -0.969704
+ 1.857e+11Hz 0.12221 -0.969785
+ 1.858e+11Hz 0.121472 -0.969866
+ 1.859e+11Hz 0.120735 -0.969946
+ 1.86e+11Hz 0.119998 -0.970025
+ 1.861e+11Hz 0.11926 -0.970104
+ 1.862e+11Hz 0.118523 -0.970183
+ 1.863e+11Hz 0.117785 -0.970261
+ 1.864e+11Hz 0.117047 -0.970339
+ 1.865e+11Hz 0.11631 -0.970417
+ 1.866e+11Hz 0.115572 -0.970494
+ 1.867e+11Hz 0.114834 -0.970571
+ 1.868e+11Hz 0.114096 -0.970647
+ 1.869e+11Hz 0.113358 -0.970723
+ 1.87e+11Hz 0.11262 -0.970798
+ 1.871e+11Hz 0.111882 -0.970873
+ 1.872e+11Hz 0.111144 -0.970947
+ 1.873e+11Hz 0.110405 -0.971021
+ 1.874e+11Hz 0.109667 -0.971095
+ 1.875e+11Hz 0.108928 -0.971168
+ 1.876e+11Hz 0.10819 -0.971241
+ 1.877e+11Hz 0.107451 -0.971313
+ 1.878e+11Hz 0.106712 -0.971385
+ 1.879e+11Hz 0.105973 -0.971457
+ 1.88e+11Hz 0.105234 -0.971528
+ 1.881e+11Hz 0.104495 -0.971598
+ 1.882e+11Hz 0.103756 -0.971668
+ 1.883e+11Hz 0.103017 -0.971738
+ 1.884e+11Hz 0.102277 -0.971807
+ 1.885e+11Hz 0.101538 -0.971876
+ 1.886e+11Hz 0.100798 -0.971944
+ 1.887e+11Hz 0.100059 -0.972012
+ 1.888e+11Hz 0.0993189 -0.972079
+ 1.889e+11Hz 0.098579 -0.972146
+ 1.89e+11Hz 0.097839 -0.972213
+ 1.891e+11Hz 0.0970988 -0.972279
+ 1.892e+11Hz 0.0963586 -0.972344
+ 1.893e+11Hz 0.0956182 -0.97241
+ 1.894e+11Hz 0.0948777 -0.972474
+ 1.895e+11Hz 0.0941371 -0.972538
+ 1.896e+11Hz 0.0933963 -0.972602
+ 1.897e+11Hz 0.0926555 -0.972665
+ 1.898e+11Hz 0.0919145 -0.972728
+ 1.899e+11Hz 0.0911734 -0.97279
+ 1.9e+11Hz 0.0904321 -0.972852
+ 1.901e+11Hz 0.0896908 -0.972914
+ 1.902e+11Hz 0.0889493 -0.972974
+ 1.903e+11Hz 0.0882077 -0.973035
+ 1.904e+11Hz 0.0874659 -0.973095
+ 1.905e+11Hz 0.0867241 -0.973154
+ 1.906e+11Hz 0.0859821 -0.973213
+ 1.907e+11Hz 0.0852399 -0.973271
+ 1.908e+11Hz 0.0844977 -0.973329
+ 1.909e+11Hz 0.0837553 -0.973387
+ 1.91e+11Hz 0.0830128 -0.973444
+ 1.911e+11Hz 0.0822701 -0.9735
+ 1.912e+11Hz 0.0815273 -0.973556
+ 1.913e+11Hz 0.0807844 -0.973611
+ 1.914e+11Hz 0.0800413 -0.973666
+ 1.915e+11Hz 0.0792981 -0.97372
+ 1.916e+11Hz 0.0785548 -0.973774
+ 1.917e+11Hz 0.0778114 -0.973828
+ 1.918e+11Hz 0.0770678 -0.97388
+ 1.919e+11Hz 0.076324 -0.973933
+ 1.92e+11Hz 0.0755802 -0.973985
+ 1.921e+11Hz 0.0748362 -0.974036
+ 1.922e+11Hz 0.074092 -0.974086
+ 1.923e+11Hz 0.0733478 -0.974137
+ 1.924e+11Hz 0.0726034 -0.974186
+ 1.925e+11Hz 0.0718589 -0.974235
+ 1.926e+11Hz 0.0711142 -0.974284
+ 1.927e+11Hz 0.0703694 -0.974332
+ 1.928e+11Hz 0.0696245 -0.974379
+ 1.929e+11Hz 0.0688794 -0.974426
+ 1.93e+11Hz 0.0681342 -0.974473
+ 1.931e+11Hz 0.0673889 -0.974519
+ 1.932e+11Hz 0.0666435 -0.974564
+ 1.933e+11Hz 0.0658979 -0.974609
+ 1.934e+11Hz 0.0651522 -0.974653
+ 1.935e+11Hz 0.0644063 -0.974696
+ 1.936e+11Hz 0.0636604 -0.974739
+ 1.937e+11Hz 0.0629143 -0.974782
+ 1.938e+11Hz 0.0621681 -0.974824
+ 1.939e+11Hz 0.0614217 -0.974865
+ 1.94e+11Hz 0.0606753 -0.974906
+ 1.941e+11Hz 0.0599287 -0.974946
+ 1.942e+11Hz 0.059182 -0.974985
+ 1.943e+11Hz 0.0584352 -0.975025
+ 1.944e+11Hz 0.0576883 -0.975063
+ 1.945e+11Hz 0.0569412 -0.975101
+ 1.946e+11Hz 0.056194 -0.975138
+ 1.947e+11Hz 0.0554468 -0.975175
+ 1.948e+11Hz 0.0546994 -0.975211
+ 1.949e+11Hz 0.0539519 -0.975246
+ 1.95e+11Hz 0.0532043 -0.975281
+ 1.951e+11Hz 0.0524565 -0.975316
+ 1.952e+11Hz 0.0517087 -0.975349
+ 1.953e+11Hz 0.0509608 -0.975382
+ 1.954e+11Hz 0.0502128 -0.975415
+ 1.955e+11Hz 0.0494646 -0.975447
+ 1.956e+11Hz 0.0487164 -0.975478
+ 1.957e+11Hz 0.0479681 -0.975509
+ 1.958e+11Hz 0.0472196 -0.975539
+ 1.959e+11Hz 0.0464711 -0.975568
+ 1.96e+11Hz 0.0457225 -0.975597
+ 1.961e+11Hz 0.0449738 -0.975625
+ 1.962e+11Hz 0.044225 -0.975653
+ 1.963e+11Hz 0.0434761 -0.97568
+ 1.964e+11Hz 0.0427272 -0.975706
+ 1.965e+11Hz 0.0419781 -0.975732
+ 1.966e+11Hz 0.041229 -0.975757
+ 1.967e+11Hz 0.0404798 -0.975782
+ 1.968e+11Hz 0.0397305 -0.975806
+ 1.969e+11Hz 0.0389812 -0.975829
+ 1.97e+11Hz 0.0382317 -0.975852
+ 1.971e+11Hz 0.0374822 -0.975874
+ 1.972e+11Hz 0.0367327 -0.975895
+ 1.973e+11Hz 0.035983 -0.975916
+ 1.974e+11Hz 0.0352333 -0.975936
+ 1.975e+11Hz 0.0344836 -0.975955
+ 1.976e+11Hz 0.0337338 -0.975974
+ 1.977e+11Hz 0.0329839 -0.975992
+ 1.978e+11Hz 0.032234 -0.97601
+ 1.979e+11Hz 0.031484 -0.976027
+ 1.98e+11Hz 0.0307339 -0.976043
+ 1.981e+11Hz 0.0299839 -0.976059
+ 1.982e+11Hz 0.0292337 -0.976074
+ 1.983e+11Hz 0.0284836 -0.976088
+ 1.984e+11Hz 0.0277334 -0.976102
+ 1.985e+11Hz 0.0269831 -0.976115
+ 1.986e+11Hz 0.0262328 -0.976128
+ 1.987e+11Hz 0.0254825 -0.97614
+ 1.988e+11Hz 0.0247321 -0.976151
+ 1.989e+11Hz 0.0239817 -0.976161
+ 1.99e+11Hz 0.0232313 -0.976171
+ 1.991e+11Hz 0.0224809 -0.976181
+ 1.992e+11Hz 0.0217304 -0.976189
+ 1.993e+11Hz 0.0209799 -0.976197
+ 1.994e+11Hz 0.0202294 -0.976205
+ 1.995e+11Hz 0.0194789 -0.976211
+ 1.996e+11Hz 0.0187284 -0.976217
+ 1.997e+11Hz 0.0179778 -0.976223
+ 1.998e+11Hz 0.0172273 -0.976227
+ 1.999e+11Hz 0.0164767 -0.976232
+ 2e+11Hz 0.0157261 -0.976235
+ 2.001e+11Hz 0.0149755 -0.976238
+ 2.002e+11Hz 0.014225 -0.97624
+ 2.003e+11Hz 0.0134744 -0.976242
+ 2.004e+11Hz 0.0127238 -0.976242
+ 2.005e+11Hz 0.0119732 -0.976243
+ 2.006e+11Hz 0.0112227 -0.976242
+ 2.007e+11Hz 0.0104721 -0.976241
+ 2.008e+11Hz 0.00972156 -0.97624
+ 2.009e+11Hz 0.00897103 -0.976237
+ 2.01e+11Hz 0.00822051 -0.976234
+ 2.011e+11Hz 0.00747001 -0.976231
+ 2.012e+11Hz 0.00671953 -0.976226
+ 2.013e+11Hz 0.00596907 -0.976222
+ 2.014e+11Hz 0.00521864 -0.976216
+ 2.015e+11Hz 0.00446823 -0.97621
+ 2.016e+11Hz 0.00371784 -0.976203
+ 2.017e+11Hz 0.00296749 -0.976196
+ 2.018e+11Hz 0.00221717 -0.976187
+ 2.019e+11Hz 0.00146688 -0.976179
+ 2.02e+11Hz 0.00071662 -0.976169
+ 2.021e+11Hz -3.35995e-05 -0.976159
+ 2.022e+11Hz -0.00078378 -0.976149
+ 2.023e+11Hz -0.00153392 -0.976137
+ 2.024e+11Hz -0.00228402 -0.976125
+ 2.025e+11Hz -0.00303408 -0.976113
+ 2.026e+11Hz -0.00378409 -0.9761
+ 2.027e+11Hz -0.00453405 -0.976086
+ 2.028e+11Hz -0.00528396 -0.976071
+ 2.029e+11Hz -0.00603383 -0.976056
+ 2.03e+11Hz -0.00678364 -0.97604
+ 2.031e+11Hz -0.0075334 -0.976024
+ 2.032e+11Hz -0.0082831 -0.976007
+ 2.033e+11Hz -0.00903275 -0.975989
+ 2.034e+11Hz -0.00978234 -0.975971
+ 2.035e+11Hz -0.0105319 -0.975952
+ 2.036e+11Hz -0.0112813 -0.975933
+ 2.037e+11Hz -0.0120307 -0.975913
+ 2.038e+11Hz -0.0127801 -0.975892
+ 2.039e+11Hz -0.0135294 -0.97587
+ 2.04e+11Hz -0.0142786 -0.975848
+ 2.041e+11Hz -0.0150277 -0.975826
+ 2.042e+11Hz -0.0157768 -0.975802
+ 2.043e+11Hz -0.0165258 -0.975779
+ 2.044e+11Hz -0.0172747 -0.975754
+ 2.045e+11Hz -0.0180236 -0.975729
+ 2.046e+11Hz -0.0187723 -0.975703
+ 2.047e+11Hz -0.019521 -0.975677
+ 2.048e+11Hz -0.0202697 -0.97565
+ 2.049e+11Hz -0.0210182 -0.975622
+ 2.05e+11Hz -0.0217667 -0.975594
+ 2.051e+11Hz -0.0225151 -0.975565
+ 2.052e+11Hz -0.0232634 -0.975536
+ 2.053e+11Hz -0.0240116 -0.975506
+ 2.054e+11Hz -0.0247597 -0.975475
+ 2.055e+11Hz -0.0255078 -0.975444
+ 2.056e+11Hz -0.0262557 -0.975412
+ 2.057e+11Hz -0.0270036 -0.975379
+ 2.058e+11Hz -0.0277514 -0.975346
+ 2.059e+11Hz -0.0284991 -0.975312
+ 2.06e+11Hz -0.0292467 -0.975278
+ 2.061e+11Hz -0.0299942 -0.975243
+ 2.062e+11Hz -0.0307416 -0.975208
+ 2.063e+11Hz -0.0314889 -0.975171
+ 2.064e+11Hz -0.0322361 -0.975135
+ 2.065e+11Hz -0.0329833 -0.975097
+ 2.066e+11Hz -0.0337303 -0.975059
+ 2.067e+11Hz -0.0344772 -0.975021
+ 2.068e+11Hz -0.0352241 -0.974982
+ 2.069e+11Hz -0.0359708 -0.974942
+ 2.07e+11Hz -0.0367175 -0.974901
+ 2.071e+11Hz -0.037464 -0.97486
+ 2.072e+11Hz -0.0382104 -0.974819
+ 2.073e+11Hz -0.0389567 -0.974777
+ 2.074e+11Hz -0.039703 -0.974734
+ 2.075e+11Hz -0.0404491 -0.974691
+ 2.076e+11Hz -0.0411951 -0.974647
+ 2.077e+11Hz -0.041941 -0.974602
+ 2.078e+11Hz -0.0426868 -0.974557
+ 2.079e+11Hz -0.0434324 -0.974511
+ 2.08e+11Hz -0.044178 -0.974465
+ 2.081e+11Hz -0.0449235 -0.974418
+ 2.082e+11Hz -0.0456688 -0.97437
+ 2.083e+11Hz -0.046414 -0.974322
+ 2.084e+11Hz -0.0471591 -0.974274
+ 2.085e+11Hz -0.0479041 -0.974224
+ 2.086e+11Hz -0.048649 -0.974174
+ 2.087e+11Hz -0.0493938 -0.974124
+ 2.088e+11Hz -0.0501384 -0.974073
+ 2.089e+11Hz -0.050883 -0.974021
+ 2.09e+11Hz -0.0516274 -0.973969
+ 2.091e+11Hz -0.0523716 -0.973916
+ 2.092e+11Hz -0.0531158 -0.973863
+ 2.093e+11Hz -0.0538598 -0.973809
+ 2.094e+11Hz -0.0546038 -0.973754
+ 2.095e+11Hz -0.0553475 -0.973699
+ 2.096e+11Hz -0.0560912 -0.973644
+ 2.097e+11Hz -0.0568347 -0.973587
+ 2.098e+11Hz -0.0575781 -0.97353
+ 2.099e+11Hz -0.0583214 -0.973473
+ 2.1e+11Hz -0.0590646 -0.973415
+ 2.101e+11Hz -0.0598076 -0.973356
+ 2.102e+11Hz -0.0605504 -0.973297
+ 2.103e+11Hz -0.0612932 -0.973237
+ 2.104e+11Hz -0.0620358 -0.973177
+ 2.105e+11Hz -0.0627783 -0.973116
+ 2.106e+11Hz -0.0635206 -0.973055
+ 2.107e+11Hz -0.0642628 -0.972992
+ 2.108e+11Hz -0.0650049 -0.97293
+ 2.109e+11Hz -0.0657468 -0.972867
+ 2.11e+11Hz -0.0664885 -0.972803
+ 2.111e+11Hz -0.0672302 -0.972739
+ 2.112e+11Hz -0.0679717 -0.972674
+ 2.113e+11Hz -0.068713 -0.972608
+ 2.114e+11Hz -0.0694542 -0.972542
+ 2.115e+11Hz -0.0701952 -0.972475
+ 2.116e+11Hz -0.0709361 -0.972408
+ 2.117e+11Hz -0.0716769 -0.97234
+ 2.118e+11Hz -0.0724175 -0.972272
+ 2.119e+11Hz -0.0731579 -0.972203
+ 2.12e+11Hz -0.0738982 -0.972134
+ 2.121e+11Hz -0.0746383 -0.972064
+ 2.122e+11Hz -0.0753783 -0.971993
+ 2.123e+11Hz -0.0761181 -0.971922
+ 2.124e+11Hz -0.0768577 -0.97185
+ 2.125e+11Hz -0.0775972 -0.971778
+ 2.126e+11Hz -0.0783366 -0.971705
+ 2.127e+11Hz -0.0790757 -0.971632
+ 2.128e+11Hz -0.0798147 -0.971558
+ 2.129e+11Hz -0.0805536 -0.971484
+ 2.13e+11Hz -0.0812922 -0.971409
+ 2.131e+11Hz -0.0820307 -0.971333
+ 2.132e+11Hz -0.0827691 -0.971257
+ 2.133e+11Hz -0.0835072 -0.97118
+ 2.134e+11Hz -0.0842452 -0.971103
+ 2.135e+11Hz -0.084983 -0.971026
+ 2.136e+11Hz -0.0857206 -0.970947
+ 2.137e+11Hz -0.0864581 -0.970868
+ 2.138e+11Hz -0.0871954 -0.970789
+ 2.139e+11Hz -0.0879325 -0.970709
+ 2.14e+11Hz -0.0886694 -0.970629
+ 2.141e+11Hz -0.0894061 -0.970548
+ 2.142e+11Hz -0.0901427 -0.970466
+ 2.143e+11Hz -0.090879 -0.970384
+ 2.144e+11Hz -0.0916152 -0.970302
+ 2.145e+11Hz -0.0923512 -0.970219
+ 2.146e+11Hz -0.093087 -0.970135
+ 2.147e+11Hz -0.0938226 -0.970051
+ 2.148e+11Hz -0.0945581 -0.969966
+ 2.149e+11Hz -0.0952933 -0.969881
+ 2.15e+11Hz -0.0960283 -0.969795
+ 2.151e+11Hz -0.0967632 -0.969709
+ 2.152e+11Hz -0.0974978 -0.969622
+ 2.153e+11Hz -0.0982323 -0.969535
+ 2.154e+11Hz -0.0989665 -0.969447
+ 2.155e+11Hz -0.0997006 -0.969359
+ 2.156e+11Hz -0.100434 -0.96927
+ 2.157e+11Hz -0.101168 -0.969181
+ 2.158e+11Hz -0.101902 -0.969091
+ 2.159e+11Hz -0.102635 -0.969001
+ 2.16e+11Hz -0.103368 -0.96891
+ 2.161e+11Hz -0.104101 -0.968819
+ 2.162e+11Hz -0.104833 -0.968727
+ 2.163e+11Hz -0.105566 -0.968635
+ 2.164e+11Hz -0.106298 -0.968542
+ 2.165e+11Hz -0.10703 -0.968449
+ 2.166e+11Hz -0.107762 -0.968355
+ 2.167e+11Hz -0.108493 -0.968261
+ 2.168e+11Hz -0.109225 -0.968166
+ 2.169e+11Hz -0.109956 -0.968071
+ 2.17e+11Hz -0.110687 -0.967976
+ 2.171e+11Hz -0.111418 -0.96788
+ 2.172e+11Hz -0.112148 -0.967783
+ 2.173e+11Hz -0.112878 -0.967686
+ 2.174e+11Hz -0.113608 -0.967589
+ 2.175e+11Hz -0.114338 -0.967491
+ 2.176e+11Hz -0.115068 -0.967392
+ 2.177e+11Hz -0.115797 -0.967294
+ 2.178e+11Hz -0.116527 -0.967194
+ 2.179e+11Hz -0.117256 -0.967095
+ 2.18e+11Hz -0.117984 -0.966995
+ 2.181e+11Hz -0.118713 -0.966894
+ 2.182e+11Hz -0.119441 -0.966793
+ 2.183e+11Hz -0.12017 -0.966691
+ 2.184e+11Hz -0.120898 -0.96659
+ 2.185e+11Hz -0.121625 -0.966487
+ 2.186e+11Hz -0.122353 -0.966385
+ 2.187e+11Hz -0.12308 -0.966281
+ 2.188e+11Hz -0.123807 -0.966178
+ 2.189e+11Hz -0.124534 -0.966074
+ 2.19e+11Hz -0.125261 -0.96597
+ 2.191e+11Hz -0.125987 -0.965865
+ 2.192e+11Hz -0.126713 -0.96576
+ 2.193e+11Hz -0.127439 -0.965654
+ 2.194e+11Hz -0.128165 -0.965548
+ 2.195e+11Hz -0.128891 -0.965442
+ 2.196e+11Hz -0.129616 -0.965335
+ 2.197e+11Hz -0.130341 -0.965228
+ 2.198e+11Hz -0.131066 -0.96512
+ 2.199e+11Hz -0.131791 -0.965012
+ 2.2e+11Hz -0.132516 -0.964904
+ 2.201e+11Hz -0.13324 -0.964795
+ 2.202e+11Hz -0.133964 -0.964686
+ 2.203e+11Hz -0.134688 -0.964577
+ 2.204e+11Hz -0.135412 -0.964467
+ 2.205e+11Hz -0.136136 -0.964357
+ 2.206e+11Hz -0.136859 -0.964247
+ 2.207e+11Hz -0.137582 -0.964136
+ 2.208e+11Hz -0.138305 -0.964025
+ 2.209e+11Hz -0.139028 -0.963913
+ 2.21e+11Hz -0.139751 -0.963801
+ 2.211e+11Hz -0.140473 -0.963689
+ 2.212e+11Hz -0.141195 -0.963576
+ 2.213e+11Hz -0.141917 -0.963464
+ 2.214e+11Hz -0.142639 -0.96335
+ 2.215e+11Hz -0.143361 -0.963237
+ 2.216e+11Hz -0.144083 -0.963123
+ 2.217e+11Hz -0.144804 -0.963009
+ 2.218e+11Hz -0.145525 -0.962894
+ 2.219e+11Hz -0.146246 -0.96278
+ 2.22e+11Hz -0.146967 -0.962665
+ 2.221e+11Hz -0.147688 -0.962549
+ 2.222e+11Hz -0.148409 -0.962433
+ 2.223e+11Hz -0.149129 -0.962317
+ 2.224e+11Hz -0.149849 -0.962201
+ 2.225e+11Hz -0.15057 -0.962085
+ 2.226e+11Hz -0.15129 -0.961968
+ 2.227e+11Hz -0.152009 -0.96185
+ 2.228e+11Hz -0.152729 -0.961733
+ 2.229e+11Hz -0.153449 -0.961615
+ 2.23e+11Hz -0.154168 -0.961497
+ 2.231e+11Hz -0.154888 -0.961379
+ 2.232e+11Hz -0.155607 -0.96126
+ 2.233e+11Hz -0.156326 -0.961141
+ 2.234e+11Hz -0.157045 -0.961022
+ 2.235e+11Hz -0.157764 -0.960903
+ 2.236e+11Hz -0.158483 -0.960783
+ 2.237e+11Hz -0.159202 -0.960663
+ 2.238e+11Hz -0.15992 -0.960543
+ 2.239e+11Hz -0.160639 -0.960422
+ 2.24e+11Hz -0.161357 -0.960302
+ 2.241e+11Hz -0.162076 -0.960181
+ 2.242e+11Hz -0.162794 -0.960059
+ 2.243e+11Hz -0.163512 -0.959938
+ 2.244e+11Hz -0.16423 -0.959816
+ 2.245e+11Hz -0.164948 -0.959694
+ 2.246e+11Hz -0.165667 -0.959572
+ 2.247e+11Hz -0.166385 -0.959449
+ 2.248e+11Hz -0.167102 -0.959326
+ 2.249e+11Hz -0.16782 -0.959203
+ 2.25e+11Hz -0.168538 -0.95908
+ 2.251e+11Hz -0.169256 -0.958956
+ 2.252e+11Hz -0.169974 -0.958832
+ 2.253e+11Hz -0.170692 -0.958708
+ 2.254e+11Hz -0.17141 -0.958584
+ 2.255e+11Hz -0.172127 -0.958459
+ 2.256e+11Hz -0.172845 -0.958335
+ 2.257e+11Hz -0.173563 -0.95821
+ 2.258e+11Hz -0.174281 -0.958084
+ 2.259e+11Hz -0.174999 -0.957959
+ 2.26e+11Hz -0.175716 -0.957833
+ 2.261e+11Hz -0.176434 -0.957707
+ 2.262e+11Hz -0.177152 -0.95758
+ 2.263e+11Hz -0.17787 -0.957454
+ 2.264e+11Hz -0.178588 -0.957327
+ 2.265e+11Hz -0.179306 -0.9572
+ 2.266e+11Hz -0.180024 -0.957073
+ 2.267e+11Hz -0.180742 -0.956945
+ 2.268e+11Hz -0.18146 -0.956817
+ 2.269e+11Hz -0.182178 -0.956689
+ 2.27e+11Hz -0.182897 -0.956561
+ 2.271e+11Hz -0.183615 -0.956432
+ 2.272e+11Hz -0.184333 -0.956303
+ 2.273e+11Hz -0.185052 -0.956174
+ 2.274e+11Hz -0.18577 -0.956044
+ 2.275e+11Hz -0.186489 -0.955915
+ 2.276e+11Hz -0.187208 -0.955785
+ 2.277e+11Hz -0.187927 -0.955655
+ 2.278e+11Hz -0.188646 -0.955524
+ 2.279e+11Hz -0.189365 -0.955393
+ 2.28e+11Hz -0.190084 -0.955262
+ 2.281e+11Hz -0.190804 -0.955131
+ 2.282e+11Hz -0.191523 -0.954999
+ 2.283e+11Hz -0.192243 -0.954867
+ 2.284e+11Hz -0.192963 -0.954735
+ 2.285e+11Hz -0.193683 -0.954602
+ 2.286e+11Hz -0.194403 -0.954469
+ 2.287e+11Hz -0.195123 -0.954336
+ 2.288e+11Hz -0.195844 -0.954203
+ 2.289e+11Hz -0.196564 -0.954069
+ 2.29e+11Hz -0.197285 -0.953935
+ 2.291e+11Hz -0.198006 -0.9538
+ 2.292e+11Hz -0.198727 -0.953665
+ 2.293e+11Hz -0.199449 -0.95353
+ 2.294e+11Hz -0.20017 -0.953395
+ 2.295e+11Hz -0.200892 -0.953259
+ 2.296e+11Hz -0.201614 -0.953123
+ 2.297e+11Hz -0.202336 -0.952986
+ 2.298e+11Hz -0.203058 -0.952849
+ 2.299e+11Hz -0.203781 -0.952712
+ 2.3e+11Hz -0.204504 -0.952575
+ 2.301e+11Hz -0.205227 -0.952437
+ 2.302e+11Hz -0.20595 -0.952298
+ 2.303e+11Hz -0.206673 -0.952159
+ 2.304e+11Hz -0.207397 -0.95202
+ 2.305e+11Hz -0.208121 -0.951881
+ 2.306e+11Hz -0.208845 -0.951741
+ 2.307e+11Hz -0.209569 -0.951601
+ 2.308e+11Hz -0.210294 -0.95146
+ 2.309e+11Hz -0.211019 -0.951319
+ 2.31e+11Hz -0.211744 -0.951177
+ 2.311e+11Hz -0.212469 -0.951035
+ 2.312e+11Hz -0.213195 -0.950893
+ 2.313e+11Hz -0.213921 -0.95075
+ 2.314e+11Hz -0.214647 -0.950606
+ 2.315e+11Hz -0.215374 -0.950462
+ 2.316e+11Hz -0.2161 -0.950318
+ 2.317e+11Hz -0.216827 -0.950173
+ 2.318e+11Hz -0.217554 -0.950028
+ 2.319e+11Hz -0.218282 -0.949883
+ 2.32e+11Hz -0.21901 -0.949736
+ 2.321e+11Hz -0.219738 -0.94959
+ 2.322e+11Hz -0.220466 -0.949442
+ 2.323e+11Hz -0.221195 -0.949295
+ 2.324e+11Hz -0.221923 -0.949146
+ 2.325e+11Hz -0.222653 -0.948998
+ 2.326e+11Hz -0.223382 -0.948848
+ 2.327e+11Hz -0.224112 -0.948699
+ 2.328e+11Hz -0.224842 -0.948548
+ 2.329e+11Hz -0.225572 -0.948397
+ 2.33e+11Hz -0.226302 -0.948246
+ 2.331e+11Hz -0.227033 -0.948094
+ 2.332e+11Hz -0.227764 -0.947941
+ 2.333e+11Hz -0.228495 -0.947788
+ 2.334e+11Hz -0.229227 -0.947634
+ 2.335e+11Hz -0.229959 -0.947479
+ 2.336e+11Hz -0.230691 -0.947324
+ 2.337e+11Hz -0.231424 -0.947169
+ 2.338e+11Hz -0.232156 -0.947012
+ 2.339e+11Hz -0.232889 -0.946855
+ 2.34e+11Hz -0.233623 -0.946698
+ 2.341e+11Hz -0.234356 -0.94654
+ 2.342e+11Hz -0.23509 -0.946381
+ 2.343e+11Hz -0.235824 -0.946221
+ 2.344e+11Hz -0.236558 -0.946061
+ 2.345e+11Hz -0.237293 -0.9459
+ 2.346e+11Hz -0.238028 -0.945739
+ 2.347e+11Hz -0.238763 -0.945577
+ 2.348e+11Hz -0.239498 -0.945414
+ 2.349e+11Hz -0.240234 -0.94525
+ 2.35e+11Hz -0.240969 -0.945086
+ 2.351e+11Hz -0.241706 -0.944921
+ 2.352e+11Hz -0.242442 -0.944755
+ 2.353e+11Hz -0.243178 -0.944589
+ 2.354e+11Hz -0.243915 -0.944421
+ 2.355e+11Hz -0.244652 -0.944253
+ 2.356e+11Hz -0.245389 -0.944085
+ 2.357e+11Hz -0.246127 -0.943915
+ 2.358e+11Hz -0.246865 -0.943745
+ 2.359e+11Hz -0.247602 -0.943574
+ 2.36e+11Hz -0.248341 -0.943402
+ 2.361e+11Hz -0.249079 -0.94323
+ 2.362e+11Hz -0.249817 -0.943057
+ 2.363e+11Hz -0.250556 -0.942882
+ 2.364e+11Hz -0.251295 -0.942708
+ 2.365e+11Hz -0.252034 -0.942532
+ 2.366e+11Hz -0.252773 -0.942355
+ 2.367e+11Hz -0.253513 -0.942178
+ 2.368e+11Hz -0.254252 -0.942
+ 2.369e+11Hz -0.254992 -0.941821
+ 2.37e+11Hz -0.255732 -0.941641
+ 2.371e+11Hz -0.256472 -0.94146
+ 2.372e+11Hz -0.257212 -0.941279
+ 2.373e+11Hz -0.257952 -0.941096
+ 2.374e+11Hz -0.258693 -0.940913
+ 2.375e+11Hz -0.259433 -0.940729
+ 2.376e+11Hz -0.260174 -0.940544
+ 2.377e+11Hz -0.260915 -0.940359
+ 2.378e+11Hz -0.261656 -0.940172
+ 2.379e+11Hz -0.262397 -0.939984
+ 2.38e+11Hz -0.263138 -0.939796
+ 2.381e+11Hz -0.263879 -0.939607
+ 2.382e+11Hz -0.26462 -0.939417
+ 2.383e+11Hz -0.265362 -0.939225
+ 2.384e+11Hz -0.266103 -0.939034
+ 2.385e+11Hz -0.266845 -0.938841
+ 2.386e+11Hz -0.267586 -0.938647
+ 2.387e+11Hz -0.268328 -0.938452
+ 2.388e+11Hz -0.269069 -0.938257
+ 2.389e+11Hz -0.269811 -0.93806
+ 2.39e+11Hz -0.270553 -0.937863
+ 2.391e+11Hz -0.271294 -0.937665
+ 2.392e+11Hz -0.272036 -0.937465
+ 2.393e+11Hz -0.272778 -0.937265
+ 2.394e+11Hz -0.273519 -0.937064
+ 2.395e+11Hz -0.274261 -0.936862
+ 2.396e+11Hz -0.275003 -0.936659
+ 2.397e+11Hz -0.275744 -0.936456
+ 2.398e+11Hz -0.276486 -0.936251
+ 2.399e+11Hz -0.277227 -0.936045
+ 2.4e+11Hz -0.277969 -0.935839
+ 2.401e+11Hz -0.27871 -0.935631
+ 2.402e+11Hz -0.279451 -0.935423
+ 2.403e+11Hz -0.280193 -0.935213
+ 2.404e+11Hz -0.280934 -0.935003
+ 2.405e+11Hz -0.281675 -0.934792
+ 2.406e+11Hz -0.282416 -0.93458
+ 2.407e+11Hz -0.283157 -0.934367
+ 2.408e+11Hz -0.283898 -0.934153
+ 2.409e+11Hz -0.284638 -0.933938
+ 2.41e+11Hz -0.285379 -0.933722
+ 2.411e+11Hz -0.286119 -0.933505
+ 2.412e+11Hz -0.286859 -0.933287
+ 2.413e+11Hz -0.287599 -0.933069
+ 2.414e+11Hz -0.288339 -0.932849
+ 2.415e+11Hz -0.289079 -0.932629
+ 2.416e+11Hz -0.289819 -0.932407
+ 2.417e+11Hz -0.290558 -0.932185
+ 2.418e+11Hz -0.291297 -0.931962
+ 2.419e+11Hz -0.292036 -0.931737
+ 2.42e+11Hz -0.292775 -0.931512
+ 2.421e+11Hz -0.293514 -0.931286
+ 2.422e+11Hz -0.294252 -0.931059
+ 2.423e+11Hz -0.29499 -0.930832
+ 2.424e+11Hz -0.295728 -0.930603
+ 2.425e+11Hz -0.296466 -0.930373
+ 2.426e+11Hz -0.297203 -0.930143
+ 2.427e+11Hz -0.29794 -0.929911
+ 2.428e+11Hz -0.298677 -0.929679
+ 2.429e+11Hz -0.299414 -0.929446
+ 2.43e+11Hz -0.30015 -0.929212
+ 2.431e+11Hz -0.300887 -0.928977
+ 2.432e+11Hz -0.301622 -0.928741
+ 2.433e+11Hz -0.302358 -0.928504
+ 2.434e+11Hz -0.303093 -0.928267
+ 2.435e+11Hz -0.303828 -0.928028
+ 2.436e+11Hz -0.304563 -0.927789
+ 2.437e+11Hz -0.305297 -0.927549
+ 2.438e+11Hz -0.306031 -0.927308
+ 2.439e+11Hz -0.306765 -0.927066
+ 2.44e+11Hz -0.307498 -0.926823
+ 2.441e+11Hz -0.308231 -0.926579
+ 2.442e+11Hz -0.308964 -0.926335
+ 2.443e+11Hz -0.309697 -0.92609
+ 2.444e+11Hz -0.310429 -0.925844
+ 2.445e+11Hz -0.31116 -0.925597
+ 2.446e+11Hz -0.311892 -0.925349
+ 2.447e+11Hz -0.312623 -0.925101
+ 2.448e+11Hz -0.313353 -0.924851
+ 2.449e+11Hz -0.314083 -0.924601
+ 2.45e+11Hz -0.314813 -0.92435
+ 2.451e+11Hz -0.315543 -0.924099
+ 2.452e+11Hz -0.316272 -0.923846
+ 2.453e+11Hz -0.317001 -0.923593
+ 2.454e+11Hz -0.317729 -0.923339
+ 2.455e+11Hz -0.318457 -0.923084
+ 2.456e+11Hz -0.319185 -0.922828
+ 2.457e+11Hz -0.319912 -0.922572
+ 2.458e+11Hz -0.320639 -0.922315
+ 2.459e+11Hz -0.321365 -0.922057
+ 2.46e+11Hz -0.322091 -0.921798
+ 2.461e+11Hz -0.322817 -0.921539
+ 2.462e+11Hz -0.323542 -0.921279
+ 2.463e+11Hz -0.324267 -0.921018
+ 2.464e+11Hz -0.324991 -0.920756
+ 2.465e+11Hz -0.325715 -0.920494
+ 2.466e+11Hz -0.326439 -0.920231
+ 2.467e+11Hz -0.327162 -0.919968
+ 2.468e+11Hz -0.327884 -0.919703
+ 2.469e+11Hz -0.328607 -0.919438
+ 2.47e+11Hz -0.329329 -0.919172
+ 2.471e+11Hz -0.33005 -0.918906
+ 2.472e+11Hz -0.330771 -0.918639
+ 2.473e+11Hz -0.331492 -0.918371
+ 2.474e+11Hz -0.332212 -0.918103
+ 2.475e+11Hz -0.332932 -0.917833
+ 2.476e+11Hz -0.333651 -0.917564
+ 2.477e+11Hz -0.33437 -0.917293
+ 2.478e+11Hz -0.335089 -0.917022
+ 2.479e+11Hz -0.335807 -0.91675
+ 2.48e+11Hz -0.336524 -0.916478
+ 2.481e+11Hz -0.337242 -0.916205
+ 2.482e+11Hz -0.337958 -0.915931
+ 2.483e+11Hz -0.338675 -0.915657
+ 2.484e+11Hz -0.339391 -0.915382
+ 2.485e+11Hz -0.340106 -0.915107
+ 2.486e+11Hz -0.340821 -0.914831
+ 2.487e+11Hz -0.341536 -0.914554
+ 2.488e+11Hz -0.342251 -0.914277
+ 2.489e+11Hz -0.342964 -0.913999
+ 2.49e+11Hz -0.343678 -0.91372
+ 2.491e+11Hz -0.344391 -0.913441
+ 2.492e+11Hz -0.345104 -0.913162
+ 2.493e+11Hz -0.345816 -0.912881
+ 2.494e+11Hz -0.346528 -0.912601
+ 2.495e+11Hz -0.347239 -0.912319
+ 2.496e+11Hz -0.34795 -0.912037
+ 2.497e+11Hz -0.348661 -0.911755
+ 2.498e+11Hz -0.349371 -0.911472
+ 2.499e+11Hz -0.350081 -0.911188
+ 2.5e+11Hz -0.35079 -0.910904
+ 2.501e+11Hz -0.351499 -0.910619
+ 2.502e+11Hz -0.352208 -0.910334
+ 2.503e+11Hz -0.352916 -0.910048
+ 2.504e+11Hz -0.353624 -0.909762
+ 2.505e+11Hz -0.354332 -0.909475
+ 2.506e+11Hz -0.355039 -0.909187
+ 2.507e+11Hz -0.355745 -0.908899
+ 2.508e+11Hz -0.356452 -0.908611
+ 2.509e+11Hz -0.357158 -0.908322
+ 2.51e+11Hz -0.357863 -0.908032
+ 2.511e+11Hz -0.358568 -0.907742
+ 2.512e+11Hz -0.359273 -0.907452
+ 2.513e+11Hz -0.359978 -0.907161
+ 2.514e+11Hz -0.360682 -0.906869
+ 2.515e+11Hz -0.361386 -0.906577
+ 2.516e+11Hz -0.362089 -0.906284
+ 2.517e+11Hz -0.362792 -0.905991
+ 2.518e+11Hz -0.363495 -0.905697
+ 2.519e+11Hz -0.364197 -0.905403
+ 2.52e+11Hz -0.364899 -0.905108
+ 2.521e+11Hz -0.3656 -0.904813
+ 2.522e+11Hz -0.366302 -0.904517
+ 2.523e+11Hz -0.367003 -0.904221
+ 2.524e+11Hz -0.367703 -0.903924
+ 2.525e+11Hz -0.368404 -0.903627
+ 2.526e+11Hz -0.369103 -0.903329
+ 2.527e+11Hz -0.369803 -0.903031
+ 2.528e+11Hz -0.370502 -0.902732
+ 2.529e+11Hz -0.371201 -0.902433
+ 2.53e+11Hz -0.3719 -0.902133
+ 2.531e+11Hz -0.372598 -0.901833
+ 2.532e+11Hz -0.373296 -0.901532
+ 2.533e+11Hz -0.373994 -0.901231
+ 2.534e+11Hz -0.374691 -0.900929
+ 2.535e+11Hz -0.375388 -0.900627
+ 2.536e+11Hz -0.376085 -0.900324
+ 2.537e+11Hz -0.376781 -0.90002
+ 2.538e+11Hz -0.377477 -0.899717
+ 2.539e+11Hz -0.378173 -0.899412
+ 2.54e+11Hz -0.378868 -0.899107
+ 2.541e+11Hz -0.379564 -0.898802
+ 2.542e+11Hz -0.380258 -0.898496
+ 2.543e+11Hz -0.380953 -0.89819
+ 2.544e+11Hz -0.381647 -0.897883
+ 2.545e+11Hz -0.382341 -0.897575
+ 2.546e+11Hz -0.383035 -0.897267
+ 2.547e+11Hz -0.383728 -0.896959
+ 2.548e+11Hz -0.384421 -0.89665
+ 2.549e+11Hz -0.385114 -0.89634
+ 2.55e+11Hz -0.385806 -0.89603
+ 2.551e+11Hz -0.386498 -0.89572
+ 2.552e+11Hz -0.38719 -0.895409
+ 2.553e+11Hz -0.387882 -0.895097
+ 2.554e+11Hz -0.388573 -0.894785
+ 2.555e+11Hz -0.389264 -0.894472
+ 2.556e+11Hz -0.389955 -0.894159
+ 2.557e+11Hz -0.390645 -0.893845
+ 2.558e+11Hz -0.391335 -0.893531
+ 2.559e+11Hz -0.392025 -0.893216
+ 2.56e+11Hz -0.392715 -0.892901
+ 2.561e+11Hz -0.393404 -0.892585
+ 2.562e+11Hz -0.394093 -0.892269
+ 2.563e+11Hz -0.394782 -0.891952
+ 2.564e+11Hz -0.39547 -0.891634
+ 2.565e+11Hz -0.396158 -0.891316
+ 2.566e+11Hz -0.396846 -0.890997
+ 2.567e+11Hz -0.397533 -0.890678
+ 2.568e+11Hz -0.39822 -0.890359
+ 2.569e+11Hz -0.398907 -0.890038
+ 2.57e+11Hz -0.399594 -0.889717
+ 2.571e+11Hz -0.40028 -0.889396
+ 2.572e+11Hz -0.400966 -0.889074
+ 2.573e+11Hz -0.401652 -0.888751
+ 2.574e+11Hz -0.402337 -0.888428
+ 2.575e+11Hz -0.403022 -0.888105
+ 2.576e+11Hz -0.403707 -0.88778
+ 2.577e+11Hz -0.404391 -0.887456
+ 2.578e+11Hz -0.405075 -0.88713
+ 2.579e+11Hz -0.405759 -0.886804
+ 2.58e+11Hz -0.406442 -0.886478
+ 2.581e+11Hz -0.407125 -0.886151
+ 2.582e+11Hz -0.407808 -0.885823
+ 2.583e+11Hz -0.408491 -0.885495
+ 2.584e+11Hz -0.409173 -0.885166
+ 2.585e+11Hz -0.409855 -0.884837
+ 2.586e+11Hz -0.410536 -0.884507
+ 2.587e+11Hz -0.411217 -0.884176
+ 2.588e+11Hz -0.411898 -0.883845
+ 2.589e+11Hz -0.412578 -0.883513
+ 2.59e+11Hz -0.413258 -0.883181
+ 2.591e+11Hz -0.413938 -0.882848
+ 2.592e+11Hz -0.414617 -0.882515
+ 2.593e+11Hz -0.415296 -0.882181
+ 2.594e+11Hz -0.415975 -0.881846
+ 2.595e+11Hz -0.416653 -0.881511
+ 2.596e+11Hz -0.417331 -0.881175
+ 2.597e+11Hz -0.418009 -0.880839
+ 2.598e+11Hz -0.418686 -0.880502
+ 2.599e+11Hz -0.419363 -0.880164
+ 2.6e+11Hz -0.420039 -0.879826
+ 2.601e+11Hz -0.420715 -0.879487
+ 2.602e+11Hz -0.42139 -0.879148
+ 2.603e+11Hz -0.422066 -0.878808
+ 2.604e+11Hz -0.42274 -0.878468
+ 2.605e+11Hz -0.423415 -0.878127
+ 2.606e+11Hz -0.424089 -0.877785
+ 2.607e+11Hz -0.424762 -0.877443
+ 2.608e+11Hz -0.425435 -0.8771
+ 2.609e+11Hz -0.426108 -0.876757
+ 2.61e+11Hz -0.42678 -0.876413
+ 2.611e+11Hz -0.427452 -0.876069
+ 2.612e+11Hz -0.428124 -0.875724
+ 2.613e+11Hz -0.428794 -0.875378
+ 2.614e+11Hz -0.429465 -0.875032
+ 2.615e+11Hz -0.430135 -0.874686
+ 2.616e+11Hz -0.430805 -0.874338
+ 2.617e+11Hz -0.431474 -0.873991
+ 2.618e+11Hz -0.432143 -0.873642
+ 2.619e+11Hz -0.432811 -0.873293
+ 2.62e+11Hz -0.433479 -0.872944
+ 2.621e+11Hz -0.434146 -0.872594
+ 2.622e+11Hz -0.434813 -0.872244
+ 2.623e+11Hz -0.435479 -0.871893
+ 2.624e+11Hz -0.436145 -0.871541
+ 2.625e+11Hz -0.43681 -0.871189
+ 2.626e+11Hz -0.437475 -0.870837
+ 2.627e+11Hz -0.43814 -0.870484
+ 2.628e+11Hz -0.438803 -0.87013
+ 2.629e+11Hz -0.439467 -0.869776
+ 2.63e+11Hz -0.44013 -0.869422
+ 2.631e+11Hz -0.440792 -0.869067
+ 2.632e+11Hz -0.441454 -0.868711
+ 2.633e+11Hz -0.442115 -0.868355
+ 2.634e+11Hz -0.442776 -0.867999
+ 2.635e+11Hz -0.443437 -0.867642
+ 2.636e+11Hz -0.444096 -0.867284
+ 2.637e+11Hz -0.444756 -0.866926
+ 2.638e+11Hz -0.445415 -0.866568
+ 2.639e+11Hz -0.446073 -0.866209
+ 2.64e+11Hz -0.44673 -0.86585
+ 2.641e+11Hz -0.447388 -0.86549
+ 2.642e+11Hz -0.448044 -0.86513
+ 2.643e+11Hz -0.4487 -0.86477
+ 2.644e+11Hz -0.449356 -0.864409
+ 2.645e+11Hz -0.450011 -0.864048
+ 2.646e+11Hz -0.450666 -0.863686
+ 2.647e+11Hz -0.45132 -0.863324
+ 2.648e+11Hz -0.451973 -0.862961
+ 2.649e+11Hz -0.452626 -0.862598
+ 2.65e+11Hz -0.453278 -0.862235
+ 2.651e+11Hz -0.45393 -0.861871
+ 2.652e+11Hz -0.454581 -0.861507
+ 2.653e+11Hz -0.455232 -0.861143
+ 2.654e+11Hz -0.455882 -0.860778
+ 2.655e+11Hz -0.456532 -0.860413
+ 2.656e+11Hz -0.457181 -0.860048
+ 2.657e+11Hz -0.45783 -0.859682
+ 2.658e+11Hz -0.458478 -0.859316
+ 2.659e+11Hz -0.459125 -0.858949
+ 2.66e+11Hz -0.459772 -0.858583
+ 2.661e+11Hz -0.460419 -0.858216
+ 2.662e+11Hz -0.461065 -0.857848
+ 2.663e+11Hz -0.46171 -0.857481
+ 2.664e+11Hz -0.462355 -0.857113
+ 2.665e+11Hz -0.462999 -0.856745
+ 2.666e+11Hz -0.463643 -0.856377
+ 2.667e+11Hz -0.464286 -0.856008
+ 2.668e+11Hz -0.464929 -0.855639
+ 2.669e+11Hz -0.465571 -0.85527
+ 2.67e+11Hz -0.466213 -0.854901
+ 2.671e+11Hz -0.466854 -0.854531
+ 2.672e+11Hz -0.467495 -0.854161
+ 2.673e+11Hz -0.468135 -0.853791
+ 2.674e+11Hz -0.468775 -0.853421
+ 2.675e+11Hz -0.469414 -0.85305
+ 2.676e+11Hz -0.470053 -0.85268
+ 2.677e+11Hz -0.470691 -0.852309
+ 2.678e+11Hz -0.471329 -0.851938
+ 2.679e+11Hz -0.471966 -0.851567
+ 2.68e+11Hz -0.472603 -0.851196
+ 2.681e+11Hz -0.473239 -0.850824
+ 2.682e+11Hz -0.473875 -0.850452
+ 2.683e+11Hz -0.47451 -0.850081
+ 2.684e+11Hz -0.475145 -0.849709
+ 2.685e+11Hz -0.47578 -0.849337
+ 2.686e+11Hz -0.476414 -0.848964
+ 2.687e+11Hz -0.477048 -0.848592
+ 2.688e+11Hz -0.477681 -0.84822
+ 2.689e+11Hz -0.478314 -0.847847
+ 2.69e+11Hz -0.478946 -0.847475
+ 2.691e+11Hz -0.479578 -0.847102
+ 2.692e+11Hz -0.48021 -0.846729
+ 2.693e+11Hz -0.480841 -0.846356
+ 2.694e+11Hz -0.481472 -0.845983
+ 2.695e+11Hz -0.482102 -0.84561
+ 2.696e+11Hz -0.482732 -0.845237
+ 2.697e+11Hz -0.483362 -0.844864
+ 2.698e+11Hz -0.483992 -0.84449
+ 2.699e+11Hz -0.484621 -0.844117
+ 2.7e+11Hz -0.48525 -0.843743
+ 2.701e+11Hz -0.485878 -0.84337
+ 2.702e+11Hz -0.486506 -0.842996
+ 2.703e+11Hz -0.487134 -0.842623
+ 2.704e+11Hz -0.487761 -0.842249
+ 2.705e+11Hz -0.488389 -0.841875
+ 2.706e+11Hz -0.489016 -0.841502
+ 2.707e+11Hz -0.489642 -0.841128
+ 2.708e+11Hz -0.490269 -0.840754
+ 2.709e+11Hz -0.490895 -0.84038
+ 2.71e+11Hz -0.491521 -0.840006
+ 2.711e+11Hz -0.492147 -0.839633
+ 2.712e+11Hz -0.492772 -0.839259
+ 2.713e+11Hz -0.493398 -0.838885
+ 2.714e+11Hz -0.494023 -0.838511
+ 2.715e+11Hz -0.494648 -0.838137
+ 2.716e+11Hz -0.495272 -0.837763
+ 2.717e+11Hz -0.495897 -0.837388
+ 2.718e+11Hz -0.496522 -0.837014
+ 2.719e+11Hz -0.497146 -0.83664
+ 2.72e+11Hz -0.49777 -0.836266
+ 2.721e+11Hz -0.498394 -0.835892
+ 2.722e+11Hz -0.499018 -0.835517
+ 2.723e+11Hz -0.499642 -0.835143
+ 2.724e+11Hz -0.500265 -0.834769
+ 2.725e+11Hz -0.500889 -0.834394
+ 2.726e+11Hz -0.501513 -0.83402
+ 2.727e+11Hz -0.502136 -0.833646
+ 2.728e+11Hz -0.502759 -0.833271
+ 2.729e+11Hz -0.503383 -0.832897
+ 2.73e+11Hz -0.504006 -0.832522
+ 2.731e+11Hz -0.50463 -0.832147
+ 2.732e+11Hz -0.505253 -0.831772
+ 2.733e+11Hz -0.505876 -0.831398
+ 2.734e+11Hz -0.506499 -0.831023
+ 2.735e+11Hz -0.507123 -0.830648
+ 2.736e+11Hz -0.507746 -0.830273
+ 2.737e+11Hz -0.50837 -0.829898
+ 2.738e+11Hz -0.508993 -0.829522
+ 2.739e+11Hz -0.509616 -0.829147
+ 2.74e+11Hz -0.51024 -0.828772
+ 2.741e+11Hz -0.510864 -0.828396
+ 2.742e+11Hz -0.511487 -0.828021
+ 2.743e+11Hz -0.512111 -0.827645
+ 2.744e+11Hz -0.512735 -0.827269
+ 2.745e+11Hz -0.513359 -0.826893
+ 2.746e+11Hz -0.513983 -0.826517
+ 2.747e+11Hz -0.514607 -0.82614
+ 2.748e+11Hz -0.515232 -0.825764
+ 2.749e+11Hz -0.515856 -0.825387
+ 2.75e+11Hz -0.516481 -0.82501
+ 2.751e+11Hz -0.517106 -0.824633
+ 2.752e+11Hz -0.517731 -0.824256
+ 2.753e+11Hz -0.518356 -0.823879
+ 2.754e+11Hz -0.518981 -0.823501
+ 2.755e+11Hz -0.519607 -0.823123
+ 2.756e+11Hz -0.520232 -0.822745
+ 2.757e+11Hz -0.520858 -0.822367
+ 2.758e+11Hz -0.521484 -0.821988
+ 2.759e+11Hz -0.522111 -0.821609
+ 2.76e+11Hz -0.522737 -0.82123
+ 2.761e+11Hz -0.523364 -0.820851
+ 2.762e+11Hz -0.523991 -0.820471
+ 2.763e+11Hz -0.524618 -0.820091
+ 2.764e+11Hz -0.525246 -0.819711
+ 2.765e+11Hz -0.525873 -0.81933
+ 2.766e+11Hz -0.526501 -0.818949
+ 2.767e+11Hz -0.527129 -0.818568
+ 2.768e+11Hz -0.527758 -0.818186
+ 2.769e+11Hz -0.528386 -0.817804
+ 2.77e+11Hz -0.529015 -0.817422
+ 2.771e+11Hz -0.529645 -0.817039
+ 2.772e+11Hz -0.530274 -0.816655
+ 2.773e+11Hz -0.530904 -0.816272
+ 2.774e+11Hz -0.531534 -0.815888
+ 2.775e+11Hz -0.532164 -0.815503
+ 2.776e+11Hz -0.532795 -0.815118
+ 2.777e+11Hz -0.533426 -0.814733
+ 2.778e+11Hz -0.534057 -0.814347
+ 2.779e+11Hz -0.534688 -0.81396
+ 2.78e+11Hz -0.53532 -0.813573
+ 2.781e+11Hz -0.535952 -0.813186
+ 2.782e+11Hz -0.536584 -0.812798
+ 2.783e+11Hz -0.537217 -0.812409
+ 2.784e+11Hz -0.537849 -0.81202
+ 2.785e+11Hz -0.538482 -0.81163
+ 2.786e+11Hz -0.539116 -0.81124
+ 2.787e+11Hz -0.539749 -0.810849
+ 2.788e+11Hz -0.540383 -0.810457
+ 2.789e+11Hz -0.541017 -0.810065
+ 2.79e+11Hz -0.541652 -0.809673
+ 2.791e+11Hz -0.542287 -0.809279
+ 2.792e+11Hz -0.542921 -0.808885
+ 2.793e+11Hz -0.543557 -0.80849
+ 2.794e+11Hz -0.544192 -0.808095
+ 2.795e+11Hz -0.544828 -0.807699
+ 2.796e+11Hz -0.545464 -0.807302
+ 2.797e+11Hz -0.5461 -0.806904
+ 2.798e+11Hz -0.546736 -0.806506
+ 2.799e+11Hz -0.547373 -0.806107
+ 2.8e+11Hz -0.54801 -0.805707
+ 2.801e+11Hz -0.548647 -0.805307
+ 2.802e+11Hz -0.549284 -0.804905
+ 2.803e+11Hz -0.549921 -0.804503
+ 2.804e+11Hz -0.550559 -0.8041
+ 2.805e+11Hz -0.551197 -0.803697
+ 2.806e+11Hz -0.551835 -0.803292
+ 2.807e+11Hz -0.552473 -0.802887
+ 2.808e+11Hz -0.553111 -0.80248
+ 2.809e+11Hz -0.55375 -0.802073
+ 2.81e+11Hz -0.554389 -0.801665
+ 2.811e+11Hz -0.555027 -0.801256
+ 2.812e+11Hz -0.555666 -0.800847
+ 2.813e+11Hz -0.556305 -0.800436
+ 2.814e+11Hz -0.556945 -0.800024
+ 2.815e+11Hz -0.557584 -0.799612
+ 2.816e+11Hz -0.558223 -0.799198
+ 2.817e+11Hz -0.558863 -0.798784
+ 2.818e+11Hz -0.559502 -0.798369
+ 2.819e+11Hz -0.560142 -0.797953
+ 2.82e+11Hz -0.560781 -0.797535
+ 2.821e+11Hz -0.561421 -0.797117
+ 2.822e+11Hz -0.562061 -0.796698
+ 2.823e+11Hz -0.5627 -0.796278
+ 2.824e+11Hz -0.56334 -0.795857
+ 2.825e+11Hz -0.56398 -0.795435
+ 2.826e+11Hz -0.564619 -0.795012
+ 2.827e+11Hz -0.565259 -0.794588
+ 2.828e+11Hz -0.565899 -0.794162
+ 2.829e+11Hz -0.566538 -0.793736
+ 2.83e+11Hz -0.567178 -0.793309
+ 2.831e+11Hz -0.567817 -0.792881
+ 2.832e+11Hz -0.568456 -0.792452
+ 2.833e+11Hz -0.569096 -0.792021
+ 2.834e+11Hz -0.569735 -0.79159
+ 2.835e+11Hz -0.570374 -0.791158
+ 2.836e+11Hz -0.571012 -0.790724
+ 2.837e+11Hz -0.571651 -0.79029
+ 2.838e+11Hz -0.572289 -0.789854
+ 2.839e+11Hz -0.572928 -0.789418
+ 2.84e+11Hz -0.573566 -0.78898
+ 2.841e+11Hz -0.574204 -0.788541
+ 2.842e+11Hz -0.574841 -0.788102
+ 2.843e+11Hz -0.575479 -0.787661
+ 2.844e+11Hz -0.576116 -0.787219
+ 2.845e+11Hz -0.576753 -0.786776
+ 2.846e+11Hz -0.577389 -0.786332
+ 2.847e+11Hz -0.578026 -0.785887
+ 2.848e+11Hz -0.578662 -0.78544
+ 2.849e+11Hz -0.579297 -0.784993
+ 2.85e+11Hz -0.579933 -0.784545
+ 2.851e+11Hz -0.580568 -0.784095
+ 2.852e+11Hz -0.581202 -0.783645
+ 2.853e+11Hz -0.581836 -0.783193
+ 2.854e+11Hz -0.58247 -0.782741
+ 2.855e+11Hz -0.583104 -0.782287
+ 2.856e+11Hz -0.583737 -0.781833
+ 2.857e+11Hz -0.58437 -0.781377
+ 2.858e+11Hz -0.585002 -0.78092
+ 2.859e+11Hz -0.585633 -0.780462
+ 2.86e+11Hz -0.586265 -0.780003
+ 2.861e+11Hz -0.586896 -0.779544
+ 2.862e+11Hz -0.587526 -0.779083
+ 2.863e+11Hz -0.588156 -0.778621
+ 2.864e+11Hz -0.588785 -0.778158
+ 2.865e+11Hz -0.589414 -0.777694
+ 2.866e+11Hz -0.590042 -0.777229
+ 2.867e+11Hz -0.59067 -0.776763
+ 2.868e+11Hz -0.591297 -0.776296
+ 2.869e+11Hz -0.591923 -0.775828
+ 2.87e+11Hz -0.592549 -0.775359
+ 2.871e+11Hz -0.593175 -0.774889
+ 2.872e+11Hz -0.593799 -0.774418
+ 2.873e+11Hz -0.594423 -0.773946
+ 2.874e+11Hz -0.595047 -0.773473
+ 2.875e+11Hz -0.59567 -0.773
+ 2.876e+11Hz -0.596292 -0.772525
+ 2.877e+11Hz -0.596914 -0.772049
+ 2.878e+11Hz -0.597535 -0.771573
+ 2.879e+11Hz -0.598155 -0.771095
+ 2.88e+11Hz -0.598774 -0.770617
+ 2.881e+11Hz -0.599393 -0.770138
+ 2.882e+11Hz -0.600011 -0.769658
+ 2.883e+11Hz -0.600629 -0.769177
+ 2.884e+11Hz -0.601246 -0.768695
+ 2.885e+11Hz -0.601862 -0.768212
+ 2.886e+11Hz -0.602477 -0.767729
+ 2.887e+11Hz -0.603091 -0.767245
+ 2.888e+11Hz -0.603705 -0.766759
+ 2.889e+11Hz -0.604318 -0.766273
+ 2.89e+11Hz -0.604931 -0.765787
+ 2.891e+11Hz -0.605542 -0.765299
+ 2.892e+11Hz -0.606153 -0.764811
+ 2.893e+11Hz -0.606763 -0.764322
+ 2.894e+11Hz -0.607372 -0.763832
+ 2.895e+11Hz -0.607981 -0.763341
+ 2.896e+11Hz -0.608588 -0.76285
+ 2.897e+11Hz -0.609195 -0.762358
+ 2.898e+11Hz -0.609801 -0.761865
+ 2.899e+11Hz -0.610407 -0.761372
+ 2.9e+11Hz -0.611011 -0.760878
+ 2.901e+11Hz -0.611615 -0.760383
+ 2.902e+11Hz -0.612218 -0.759888
+ 2.903e+11Hz -0.61282 -0.759392
+ 2.904e+11Hz -0.613421 -0.758895
+ 2.905e+11Hz -0.614021 -0.758398
+ 2.906e+11Hz -0.614621 -0.7579
+ 2.907e+11Hz -0.61522 -0.757401
+ 2.908e+11Hz -0.615818 -0.756902
+ 2.909e+11Hz -0.616415 -0.756402
+ 2.91e+11Hz -0.617011 -0.755902
+ 2.911e+11Hz -0.617607 -0.755401
+ 2.912e+11Hz -0.618202 -0.7549
+ 2.913e+11Hz -0.618796 -0.754398
+ 2.914e+11Hz -0.619389 -0.753896
+ 2.915e+11Hz -0.619981 -0.753393
+ 2.916e+11Hz -0.620573 -0.752889
+ 2.917e+11Hz -0.621163 -0.752385
+ 2.918e+11Hz -0.621753 -0.751881
+ 2.919e+11Hz -0.622342 -0.751376
+ 2.92e+11Hz -0.622931 -0.750871
+ 2.921e+11Hz -0.623518 -0.750365
+ 2.922e+11Hz -0.624105 -0.749859
+ 2.923e+11Hz -0.624691 -0.749352
+ 2.924e+11Hz -0.625276 -0.748845
+ 2.925e+11Hz -0.625861 -0.748338
+ 2.926e+11Hz -0.626444 -0.74783
+ 2.927e+11Hz -0.627027 -0.747322
+ 2.928e+11Hz -0.627609 -0.746813
+ 2.929e+11Hz -0.628191 -0.746304
+ 2.93e+11Hz -0.628771 -0.745795
+ 2.931e+11Hz -0.629351 -0.745285
+ 2.932e+11Hz -0.62993 -0.744775
+ 2.933e+11Hz -0.630509 -0.744264
+ 2.934e+11Hz -0.631086 -0.743754
+ 2.935e+11Hz -0.631663 -0.743243
+ 2.936e+11Hz -0.63224 -0.742731
+ 2.937e+11Hz -0.632815 -0.74222
+ 2.938e+11Hz -0.63339 -0.741708
+ 2.939e+11Hz -0.633964 -0.741195
+ 2.94e+11Hz -0.634538 -0.740683
+ 2.941e+11Hz -0.63511 -0.74017
+ 2.942e+11Hz -0.635683 -0.739657
+ 2.943e+11Hz -0.636254 -0.739143
+ 2.944e+11Hz -0.636825 -0.73863
+ 2.945e+11Hz -0.637395 -0.738116
+ 2.946e+11Hz -0.637965 -0.737602
+ 2.947e+11Hz -0.638533 -0.737087
+ 2.948e+11Hz -0.639102 -0.736573
+ 2.949e+11Hz -0.639669 -0.736058
+ 2.95e+11Hz -0.640237 -0.735543
+ 2.951e+11Hz -0.640803 -0.735027
+ 2.952e+11Hz -0.641369 -0.734512
+ 2.953e+11Hz -0.641934 -0.733996
+ 2.954e+11Hz -0.642499 -0.73348
+ 2.955e+11Hz -0.643063 -0.732963
+ 2.956e+11Hz -0.643627 -0.732447
+ 2.957e+11Hz -0.64419 -0.73193
+ 2.958e+11Hz -0.644752 -0.731413
+ 2.959e+11Hz -0.645314 -0.730896
+ 2.96e+11Hz -0.645876 -0.730378
+ 2.961e+11Hz -0.646437 -0.729861
+ 2.962e+11Hz -0.646997 -0.729343
+ 2.963e+11Hz -0.647557 -0.728825
+ 2.964e+11Hz -0.648117 -0.728307
+ 2.965e+11Hz -0.648676 -0.727788
+ 2.966e+11Hz -0.649235 -0.727269
+ 2.967e+11Hz -0.649793 -0.72675
+ 2.968e+11Hz -0.65035 -0.726231
+ 2.969e+11Hz -0.650908 -0.725712
+ 2.97e+11Hz -0.651464 -0.725192
+ 2.971e+11Hz -0.652021 -0.724672
+ 2.972e+11Hz -0.652577 -0.724152
+ 2.973e+11Hz -0.653132 -0.723631
+ 2.974e+11Hz -0.653687 -0.723111
+ 2.975e+11Hz -0.654242 -0.72259
+ 2.976e+11Hz -0.654797 -0.722069
+ 2.977e+11Hz -0.655351 -0.721547
+ 2.978e+11Hz -0.655904 -0.721026
+ 2.979e+11Hz -0.656457 -0.720504
+ 2.98e+11Hz -0.65701 -0.719981
+ 2.981e+11Hz -0.657563 -0.719459
+ 2.982e+11Hz -0.658115 -0.718936
+ 2.983e+11Hz -0.658667 -0.718413
+ 2.984e+11Hz -0.659218 -0.71789
+ 2.985e+11Hz -0.659769 -0.717366
+ 2.986e+11Hz -0.66032 -0.716842
+ 2.987e+11Hz -0.66087 -0.716318
+ 2.988e+11Hz -0.66142 -0.715793
+ 2.989e+11Hz -0.66197 -0.715268
+ 2.99e+11Hz -0.66252 -0.714743
+ 2.991e+11Hz -0.663069 -0.714218
+ 2.992e+11Hz -0.663618 -0.713692
+ 2.993e+11Hz -0.664166 -0.713165
+ 2.994e+11Hz -0.664715 -0.712639
+ 2.995e+11Hz -0.665262 -0.712112
+ 2.996e+11Hz -0.66581 -0.711584
+ 2.997e+11Hz -0.666357 -0.711057
+ 2.998e+11Hz -0.666905 -0.710528
+ 2.999e+11Hz -0.667451 -0.71
+ 3e+11Hz -0.667998 -0.709471
+ ]

A21 %vd(10 3) %vd(21, 22) xfer3
.model xfer3 xfer R_I=true table=[
+ 0Hz 0.995382 0
+ 1e+08Hz 0.995382 -0.000812217
+ 2e+08Hz 0.99538 -0.00162442
+ 3e+08Hz 0.995377 -0.0024366
+ 4e+08Hz 0.995372 -0.00324873
+ 5e+08Hz 0.995367 -0.00406082
+ 6e+08Hz 0.99536 -0.00487284
+ 7e+08Hz 0.995352 -0.00568478
+ 8e+08Hz 0.995343 -0.00649662
+ 9e+08Hz 0.995333 -0.00730836
+ 1e+09Hz 0.995321 -0.00811999
+ 1.1e+09Hz 0.995308 -0.00893148
+ 1.2e+09Hz 0.995294 -0.00974282
+ 1.3e+09Hz 0.995279 -0.010554
+ 1.4e+09Hz 0.995263 -0.011365
+ 1.5e+09Hz 0.995245 -0.0121759
+ 1.6e+09Hz 0.995226 -0.0129865
+ 1.7e+09Hz 0.995206 -0.013797
+ 1.8e+09Hz 0.995185 -0.0146072
+ 1.9e+09Hz 0.995163 -0.0154172
+ 2e+09Hz 0.995139 -0.0162269
+ 2.1e+09Hz 0.995115 -0.0170364
+ 2.2e+09Hz 0.995089 -0.0178456
+ 2.3e+09Hz 0.995062 -0.0186546
+ 2.4e+09Hz 0.995034 -0.0194632
+ 2.5e+09Hz 0.995005 -0.0202716
+ 2.6e+09Hz 0.994974 -0.0210796
+ 2.7e+09Hz 0.994943 -0.0218873
+ 2.8e+09Hz 0.99491 -0.0226947
+ 2.9e+09Hz 0.994876 -0.0235018
+ 3e+09Hz 0.994841 -0.0243085
+ 3.1e+09Hz 0.994806 -0.0251148
+ 3.2e+09Hz 0.994768 -0.0259208
+ 3.3e+09Hz 0.99473 -0.0267263
+ 3.4e+09Hz 0.994691 -0.0275315
+ 3.5e+09Hz 0.994651 -0.0283363
+ 3.6e+09Hz 0.99461 -0.0291407
+ 3.7e+09Hz 0.994567 -0.0299446
+ 3.8e+09Hz 0.994524 -0.0307482
+ 3.9e+09Hz 0.99448 -0.0315512
+ 4e+09Hz 0.994434 -0.0323539
+ 4.1e+09Hz 0.994388 -0.0331561
+ 4.2e+09Hz 0.99434 -0.0339578
+ 4.3e+09Hz 0.994292 -0.0347591
+ 4.4e+09Hz 0.994243 -0.0355599
+ 4.5e+09Hz 0.994192 -0.0363602
+ 4.6e+09Hz 0.994141 -0.0371601
+ 4.7e+09Hz 0.994089 -0.0379594
+ 4.8e+09Hz 0.994036 -0.0387583
+ 4.9e+09Hz 0.993982 -0.0395566
+ 5e+09Hz 0.993927 -0.0403545
+ 5.1e+09Hz 0.993871 -0.0411518
+ 5.2e+09Hz 0.993814 -0.0419486
+ 5.3e+09Hz 0.993757 -0.0427449
+ 5.4e+09Hz 0.993698 -0.0435407
+ 5.5e+09Hz 0.993639 -0.0443359
+ 5.6e+09Hz 0.993579 -0.0451306
+ 5.7e+09Hz 0.993518 -0.0459248
+ 5.8e+09Hz 0.993456 -0.0467184
+ 5.9e+09Hz 0.993394 -0.0475115
+ 6e+09Hz 0.99333 -0.048304
+ 6.1e+09Hz 0.993266 -0.049096
+ 6.2e+09Hz 0.993201 -0.0498875
+ 6.3e+09Hz 0.993135 -0.0506783
+ 6.4e+09Hz 0.993069 -0.0514687
+ 6.5e+09Hz 0.993002 -0.0522585
+ 6.6e+09Hz 0.992934 -0.0530477
+ 6.7e+09Hz 0.992865 -0.0538364
+ 6.8e+09Hz 0.992796 -0.0546245
+ 6.9e+09Hz 0.992726 -0.0554121
+ 7e+09Hz 0.992655 -0.0561991
+ 7.1e+09Hz 0.992584 -0.0569855
+ 7.2e+09Hz 0.992512 -0.0577714
+ 7.3e+09Hz 0.992439 -0.0585568
+ 7.4e+09Hz 0.992366 -0.0593416
+ 7.5e+09Hz 0.992292 -0.0601258
+ 7.6e+09Hz 0.992217 -0.0609095
+ 7.7e+09Hz 0.992142 -0.0616927
+ 7.8e+09Hz 0.992066 -0.0624753
+ 7.9e+09Hz 0.99199 -0.0632574
+ 8e+09Hz 0.991913 -0.0640389
+ 8.1e+09Hz 0.991836 -0.0648199
+ 8.2e+09Hz 0.991758 -0.0656004
+ 8.3e+09Hz 0.991679 -0.0663804
+ 8.4e+09Hz 0.9916 -0.0671598
+ 8.5e+09Hz 0.991521 -0.0679387
+ 8.6e+09Hz 0.99144 -0.0687171
+ 8.7e+09Hz 0.99136 -0.0694949
+ 8.8e+09Hz 0.991279 -0.0702723
+ 8.9e+09Hz 0.991197 -0.0710492
+ 9e+09Hz 0.991115 -0.0718255
+ 9.1e+09Hz 0.991033 -0.0726014
+ 9.2e+09Hz 0.99095 -0.0733768
+ 9.3e+09Hz 0.990866 -0.0741517
+ 9.4e+09Hz 0.990782 -0.0749261
+ 9.5e+09Hz 0.990698 -0.0757001
+ 9.6e+09Hz 0.990613 -0.0764736
+ 9.7e+09Hz 0.990528 -0.0772466
+ 9.8e+09Hz 0.990443 -0.0780192
+ 9.9e+09Hz 0.990357 -0.0787913
+ 1e+10Hz 0.99027 -0.079563
+ 1.01e+10Hz 0.990184 -0.0803343
+ 1.02e+10Hz 0.990097 -0.0811051
+ 1.03e+10Hz 0.990009 -0.0818755
+ 1.04e+10Hz 0.989921 -0.0826455
+ 1.05e+10Hz 0.989833 -0.0834151
+ 1.06e+10Hz 0.989744 -0.0841844
+ 1.07e+10Hz 0.989655 -0.0849532
+ 1.08e+10Hz 0.989566 -0.0857216
+ 1.09e+10Hz 0.989477 -0.0864897
+ 1.1e+10Hz 0.989387 -0.0872574
+ 1.11e+10Hz 0.989296 -0.0880247
+ 1.12e+10Hz 0.989206 -0.0887917
+ 1.13e+10Hz 0.989115 -0.0895584
+ 1.14e+10Hz 0.989023 -0.0903247
+ 1.15e+10Hz 0.988932 -0.0910906
+ 1.16e+10Hz 0.98884 -0.0918563
+ 1.17e+10Hz 0.988748 -0.0926217
+ 1.18e+10Hz 0.988655 -0.0933867
+ 1.19e+10Hz 0.988563 -0.0941515
+ 1.2e+10Hz 0.988469 -0.0949159
+ 1.21e+10Hz 0.988376 -0.0956801
+ 1.22e+10Hz 0.988282 -0.096444
+ 1.23e+10Hz 0.988188 -0.0972077
+ 1.24e+10Hz 0.988094 -0.0979711
+ 1.25e+10Hz 0.988 -0.0987343
+ 1.26e+10Hz 0.987905 -0.0994972
+ 1.27e+10Hz 0.98781 -0.10026
+ 1.28e+10Hz 0.987714 -0.101022
+ 1.29e+10Hz 0.987618 -0.101785
+ 1.3e+10Hz 0.987523 -0.102547
+ 1.31e+10Hz 0.987426 -0.103309
+ 1.32e+10Hz 0.98733 -0.10407
+ 1.33e+10Hz 0.987233 -0.104832
+ 1.34e+10Hz 0.987136 -0.105593
+ 1.35e+10Hz 0.987038 -0.106354
+ 1.36e+10Hz 0.986941 -0.107115
+ 1.37e+10Hz 0.986843 -0.107876
+ 1.38e+10Hz 0.986744 -0.108637
+ 1.39e+10Hz 0.986646 -0.109397
+ 1.4e+10Hz 0.986547 -0.110158
+ 1.41e+10Hz 0.986448 -0.110918
+ 1.42e+10Hz 0.986348 -0.111678
+ 1.43e+10Hz 0.986249 -0.112438
+ 1.44e+10Hz 0.986149 -0.113198
+ 1.45e+10Hz 0.986048 -0.113958
+ 1.46e+10Hz 0.985948 -0.114718
+ 1.47e+10Hz 0.985847 -0.115478
+ 1.48e+10Hz 0.985745 -0.116237
+ 1.49e+10Hz 0.985644 -0.116997
+ 1.5e+10Hz 0.985542 -0.117756
+ 1.51e+10Hz 0.98544 -0.118516
+ 1.52e+10Hz 0.985337 -0.119275
+ 1.53e+10Hz 0.985234 -0.120035
+ 1.54e+10Hz 0.985131 -0.120794
+ 1.55e+10Hz 0.985028 -0.121554
+ 1.56e+10Hz 0.984924 -0.122313
+ 1.57e+10Hz 0.98482 -0.123072
+ 1.58e+10Hz 0.984715 -0.123831
+ 1.59e+10Hz 0.98461 -0.124591
+ 1.6e+10Hz 0.984505 -0.12535
+ 1.61e+10Hz 0.984399 -0.126109
+ 1.62e+10Hz 0.984293 -0.126869
+ 1.63e+10Hz 0.984187 -0.127628
+ 1.64e+10Hz 0.98408 -0.128387
+ 1.65e+10Hz 0.983973 -0.129147
+ 1.66e+10Hz 0.983865 -0.129906
+ 1.67e+10Hz 0.983758 -0.130665
+ 1.68e+10Hz 0.983649 -0.131425
+ 1.69e+10Hz 0.983541 -0.132184
+ 1.7e+10Hz 0.983431 -0.132944
+ 1.71e+10Hz 0.983322 -0.133703
+ 1.72e+10Hz 0.983212 -0.134463
+ 1.73e+10Hz 0.983102 -0.135222
+ 1.74e+10Hz 0.982991 -0.135982
+ 1.75e+10Hz 0.98288 -0.136742
+ 1.76e+10Hz 0.982768 -0.137502
+ 1.77e+10Hz 0.982656 -0.138262
+ 1.78e+10Hz 0.982543 -0.139021
+ 1.79e+10Hz 0.98243 -0.139781
+ 1.8e+10Hz 0.982317 -0.140541
+ 1.81e+10Hz 0.982203 -0.141302
+ 1.82e+10Hz 0.982088 -0.142062
+ 1.83e+10Hz 0.981973 -0.142822
+ 1.84e+10Hz 0.981858 -0.143582
+ 1.85e+10Hz 0.981742 -0.144343
+ 1.86e+10Hz 0.981625 -0.145103
+ 1.87e+10Hz 0.981508 -0.145863
+ 1.88e+10Hz 0.981391 -0.146624
+ 1.89e+10Hz 0.981273 -0.147385
+ 1.9e+10Hz 0.981154 -0.148145
+ 1.91e+10Hz 0.981035 -0.148906
+ 1.92e+10Hz 0.980916 -0.149667
+ 1.93e+10Hz 0.980796 -0.150428
+ 1.94e+10Hz 0.980675 -0.151189
+ 1.95e+10Hz 0.980554 -0.15195
+ 1.96e+10Hz 0.980432 -0.152711
+ 1.97e+10Hz 0.980309 -0.153472
+ 1.98e+10Hz 0.980186 -0.154233
+ 1.99e+10Hz 0.980063 -0.154995
+ 2e+10Hz 0.979939 -0.155756
+ 2.01e+10Hz 0.979814 -0.156517
+ 2.02e+10Hz 0.979689 -0.157279
+ 2.03e+10Hz 0.979563 -0.15804
+ 2.04e+10Hz 0.979436 -0.158802
+ 2.05e+10Hz 0.979309 -0.159563
+ 2.06e+10Hz 0.979182 -0.160325
+ 2.07e+10Hz 0.979053 -0.161087
+ 2.08e+10Hz 0.978924 -0.161848
+ 2.09e+10Hz 0.978795 -0.16261
+ 2.1e+10Hz 0.978665 -0.163372
+ 2.11e+10Hz 0.978534 -0.164134
+ 2.12e+10Hz 0.978402 -0.164896
+ 2.13e+10Hz 0.97827 -0.165657
+ 2.14e+10Hz 0.978137 -0.166419
+ 2.15e+10Hz 0.978004 -0.167181
+ 2.16e+10Hz 0.97787 -0.167943
+ 2.17e+10Hz 0.977735 -0.168705
+ 2.18e+10Hz 0.977599 -0.169467
+ 2.19e+10Hz 0.977463 -0.170229
+ 2.2e+10Hz 0.977327 -0.170991
+ 2.21e+10Hz 0.977189 -0.171753
+ 2.22e+10Hz 0.977051 -0.172515
+ 2.23e+10Hz 0.976912 -0.173276
+ 2.24e+10Hz 0.976773 -0.174038
+ 2.25e+10Hz 0.976633 -0.1748
+ 2.26e+10Hz 0.976492 -0.175562
+ 2.27e+10Hz 0.97635 -0.176324
+ 2.28e+10Hz 0.976208 -0.177085
+ 2.29e+10Hz 0.976065 -0.177847
+ 2.3e+10Hz 0.975921 -0.178609
+ 2.31e+10Hz 0.975777 -0.17937
+ 2.32e+10Hz 0.975632 -0.180132
+ 2.33e+10Hz 0.975486 -0.180893
+ 2.34e+10Hz 0.97534 -0.181655
+ 2.35e+10Hz 0.975192 -0.182416
+ 2.36e+10Hz 0.975045 -0.183177
+ 2.37e+10Hz 0.974896 -0.183938
+ 2.38e+10Hz 0.974747 -0.184699
+ 2.39e+10Hz 0.974597 -0.18546
+ 2.4e+10Hz 0.974446 -0.186221
+ 2.41e+10Hz 0.974294 -0.186982
+ 2.42e+10Hz 0.974142 -0.187743
+ 2.43e+10Hz 0.973989 -0.188503
+ 2.44e+10Hz 0.973836 -0.189263
+ 2.45e+10Hz 0.973682 -0.190024
+ 2.46e+10Hz 0.973527 -0.190784
+ 2.47e+10Hz 0.973371 -0.191544
+ 2.48e+10Hz 0.973214 -0.192304
+ 2.49e+10Hz 0.973057 -0.193064
+ 2.5e+10Hz 0.9729 -0.193823
+ 2.51e+10Hz 0.972741 -0.194583
+ 2.52e+10Hz 0.972582 -0.195342
+ 2.53e+10Hz 0.972422 -0.196101
+ 2.54e+10Hz 0.972261 -0.19686
+ 2.55e+10Hz 0.9721 -0.197619
+ 2.56e+10Hz 0.971938 -0.198378
+ 2.57e+10Hz 0.971775 -0.199136
+ 2.58e+10Hz 0.971611 -0.199894
+ 2.59e+10Hz 0.971447 -0.200652
+ 2.6e+10Hz 0.971282 -0.20141
+ 2.61e+10Hz 0.971117 -0.202168
+ 2.62e+10Hz 0.970951 -0.202925
+ 2.63e+10Hz 0.970784 -0.203683
+ 2.64e+10Hz 0.970616 -0.20444
+ 2.65e+10Hz 0.970448 -0.205197
+ 2.66e+10Hz 0.970279 -0.205953
+ 2.67e+10Hz 0.970109 -0.20671
+ 2.68e+10Hz 0.969939 -0.207466
+ 2.69e+10Hz 0.969768 -0.208222
+ 2.7e+10Hz 0.969596 -0.208978
+ 2.71e+10Hz 0.969424 -0.209733
+ 2.72e+10Hz 0.969251 -0.210489
+ 2.73e+10Hz 0.969077 -0.211244
+ 2.74e+10Hz 0.968903 -0.211998
+ 2.75e+10Hz 0.968728 -0.212753
+ 2.76e+10Hz 0.968552 -0.213507
+ 2.77e+10Hz 0.968376 -0.214261
+ 2.78e+10Hz 0.968199 -0.215015
+ 2.79e+10Hz 0.968021 -0.215769
+ 2.8e+10Hz 0.967843 -0.216522
+ 2.81e+10Hz 0.967664 -0.217275
+ 2.82e+10Hz 0.967485 -0.218028
+ 2.83e+10Hz 0.967304 -0.21878
+ 2.84e+10Hz 0.967124 -0.219533
+ 2.85e+10Hz 0.966942 -0.220285
+ 2.86e+10Hz 0.96676 -0.221036
+ 2.87e+10Hz 0.966578 -0.221788
+ 2.88e+10Hz 0.966395 -0.222539
+ 2.89e+10Hz 0.966211 -0.22329
+ 2.9e+10Hz 0.966026 -0.22404
+ 2.91e+10Hz 0.965842 -0.224791
+ 2.92e+10Hz 0.965656 -0.225541
+ 2.93e+10Hz 0.96547 -0.226291
+ 2.94e+10Hz 0.965283 -0.22704
+ 2.95e+10Hz 0.965096 -0.227789
+ 2.96e+10Hz 0.964908 -0.228538
+ 2.97e+10Hz 0.964719 -0.229287
+ 2.98e+10Hz 0.96453 -0.230035
+ 2.99e+10Hz 0.964341 -0.230784
+ 3e+10Hz 0.96415 -0.231531
+ 3.01e+10Hz 0.96396 -0.232279
+ 3.02e+10Hz 0.963768 -0.233026
+ 3.03e+10Hz 0.963577 -0.233773
+ 3.04e+10Hz 0.963384 -0.23452
+ 3.05e+10Hz 0.963191 -0.235266
+ 3.06e+10Hz 0.962998 -0.236013
+ 3.07e+10Hz 0.962804 -0.236758
+ 3.08e+10Hz 0.962609 -0.237504
+ 3.09e+10Hz 0.962414 -0.238249
+ 3.1e+10Hz 0.962219 -0.238994
+ 3.11e+10Hz 0.962023 -0.239739
+ 3.12e+10Hz 0.961826 -0.240484
+ 3.13e+10Hz 0.961629 -0.241228
+ 3.14e+10Hz 0.961431 -0.241972
+ 3.15e+10Hz 0.961233 -0.242716
+ 3.16e+10Hz 0.961034 -0.243459
+ 3.17e+10Hz 0.960835 -0.244202
+ 3.18e+10Hz 0.960636 -0.244945
+ 3.19e+10Hz 0.960435 -0.245688
+ 3.2e+10Hz 0.960235 -0.24643
+ 3.21e+10Hz 0.960034 -0.247172
+ 3.22e+10Hz 0.959832 -0.247914
+ 3.23e+10Hz 0.95963 -0.248656
+ 3.24e+10Hz 0.959427 -0.249397
+ 3.25e+10Hz 0.959224 -0.250138
+ 3.26e+10Hz 0.959021 -0.250879
+ 3.27e+10Hz 0.958817 -0.25162
+ 3.28e+10Hz 0.958612 -0.25236
+ 3.29e+10Hz 0.958407 -0.2531
+ 3.3e+10Hz 0.958202 -0.25384
+ 3.31e+10Hz 0.957996 -0.25458
+ 3.32e+10Hz 0.957789 -0.255319
+ 3.33e+10Hz 0.957583 -0.256058
+ 3.34e+10Hz 0.957375 -0.256797
+ 3.35e+10Hz 0.957168 -0.257536
+ 3.36e+10Hz 0.956959 -0.258275
+ 3.37e+10Hz 0.956751 -0.259013
+ 3.38e+10Hz 0.956542 -0.259751
+ 3.39e+10Hz 0.956332 -0.260489
+ 3.4e+10Hz 0.956122 -0.261227
+ 3.41e+10Hz 0.955911 -0.261964
+ 3.42e+10Hz 0.955701 -0.262701
+ 3.43e+10Hz 0.955489 -0.263438
+ 3.44e+10Hz 0.955277 -0.264175
+ 3.45e+10Hz 0.955065 -0.264912
+ 3.46e+10Hz 0.954852 -0.265649
+ 3.47e+10Hz 0.954639 -0.266385
+ 3.48e+10Hz 0.954426 -0.267121
+ 3.49e+10Hz 0.954212 -0.267857
+ 3.5e+10Hz 0.953997 -0.268593
+ 3.51e+10Hz 0.953782 -0.269328
+ 3.52e+10Hz 0.953567 -0.270064
+ 3.53e+10Hz 0.953351 -0.270799
+ 3.54e+10Hz 0.953134 -0.271534
+ 3.55e+10Hz 0.952918 -0.272269
+ 3.56e+10Hz 0.952701 -0.273003
+ 3.57e+10Hz 0.952483 -0.273738
+ 3.58e+10Hz 0.952265 -0.274472
+ 3.59e+10Hz 0.952046 -0.275207
+ 3.6e+10Hz 0.951827 -0.275941
+ 3.61e+10Hz 0.951608 -0.276675
+ 3.62e+10Hz 0.951388 -0.277409
+ 3.63e+10Hz 0.951168 -0.278142
+ 3.64e+10Hz 0.950947 -0.278876
+ 3.65e+10Hz 0.950725 -0.279609
+ 3.66e+10Hz 0.950504 -0.280342
+ 3.67e+10Hz 0.950282 -0.281075
+ 3.68e+10Hz 0.950059 -0.281808
+ 3.69e+10Hz 0.949836 -0.282541
+ 3.7e+10Hz 0.949612 -0.283274
+ 3.71e+10Hz 0.949388 -0.284007
+ 3.72e+10Hz 0.949164 -0.284739
+ 3.73e+10Hz 0.948939 -0.285471
+ 3.74e+10Hz 0.948713 -0.286204
+ 3.75e+10Hz 0.948487 -0.286936
+ 3.76e+10Hz 0.948261 -0.287668
+ 3.77e+10Hz 0.948034 -0.2884
+ 3.78e+10Hz 0.947807 -0.289132
+ 3.79e+10Hz 0.947579 -0.289863
+ 3.8e+10Hz 0.947351 -0.290595
+ 3.81e+10Hz 0.947122 -0.291326
+ 3.82e+10Hz 0.946893 -0.292058
+ 3.83e+10Hz 0.946663 -0.292789
+ 3.84e+10Hz 0.946433 -0.29352
+ 3.85e+10Hz 0.946202 -0.294251
+ 3.86e+10Hz 0.945971 -0.294982
+ 3.87e+10Hz 0.945739 -0.295713
+ 3.88e+10Hz 0.945507 -0.296444
+ 3.89e+10Hz 0.945274 -0.297175
+ 3.9e+10Hz 0.945041 -0.297905
+ 3.91e+10Hz 0.944807 -0.298636
+ 3.92e+10Hz 0.944573 -0.299366
+ 3.93e+10Hz 0.944338 -0.300097
+ 3.94e+10Hz 0.944103 -0.300827
+ 3.95e+10Hz 0.943867 -0.301557
+ 3.96e+10Hz 0.94363 -0.302287
+ 3.97e+10Hz 0.943394 -0.303017
+ 3.98e+10Hz 0.943156 -0.303747
+ 3.99e+10Hz 0.942918 -0.304477
+ 4e+10Hz 0.94268 -0.305206
+ 4.01e+10Hz 0.942441 -0.305936
+ 4.02e+10Hz 0.942201 -0.306666
+ 4.03e+10Hz 0.941961 -0.307395
+ 4.04e+10Hz 0.94172 -0.308124
+ 4.05e+10Hz 0.941479 -0.308854
+ 4.06e+10Hz 0.941237 -0.309583
+ 4.07e+10Hz 0.940995 -0.310312
+ 4.08e+10Hz 0.940752 -0.311041
+ 4.09e+10Hz 0.940509 -0.31177
+ 4.1e+10Hz 0.940265 -0.312499
+ 4.11e+10Hz 0.94002 -0.313227
+ 4.12e+10Hz 0.939775 -0.313956
+ 4.13e+10Hz 0.939529 -0.314685
+ 4.14e+10Hz 0.939283 -0.315413
+ 4.15e+10Hz 0.939036 -0.316141
+ 4.16e+10Hz 0.938789 -0.31687
+ 4.17e+10Hz 0.938541 -0.317598
+ 4.18e+10Hz 0.938292 -0.318326
+ 4.19e+10Hz 0.938043 -0.319054
+ 4.2e+10Hz 0.937793 -0.319782
+ 4.21e+10Hz 0.937543 -0.320509
+ 4.22e+10Hz 0.937292 -0.321237
+ 4.23e+10Hz 0.93704 -0.321965
+ 4.24e+10Hz 0.936788 -0.322692
+ 4.25e+10Hz 0.936535 -0.323419
+ 4.26e+10Hz 0.936282 -0.324146
+ 4.27e+10Hz 0.936028 -0.324874
+ 4.28e+10Hz 0.935773 -0.3256
+ 4.29e+10Hz 0.935518 -0.326327
+ 4.3e+10Hz 0.935262 -0.327054
+ 4.31e+10Hz 0.935006 -0.327781
+ 4.32e+10Hz 0.934749 -0.328507
+ 4.33e+10Hz 0.934491 -0.329233
+ 4.34e+10Hz 0.934233 -0.32996
+ 4.35e+10Hz 0.933974 -0.330686
+ 4.36e+10Hz 0.933714 -0.331412
+ 4.37e+10Hz 0.933454 -0.332137
+ 4.38e+10Hz 0.933193 -0.332863
+ 4.39e+10Hz 0.932932 -0.333589
+ 4.4e+10Hz 0.932669 -0.334314
+ 4.41e+10Hz 0.932407 -0.335039
+ 4.42e+10Hz 0.932143 -0.335764
+ 4.43e+10Hz 0.931879 -0.336489
+ 4.44e+10Hz 0.931615 -0.337214
+ 4.45e+10Hz 0.93135 -0.337938
+ 4.46e+10Hz 0.931084 -0.338663
+ 4.47e+10Hz 0.930817 -0.339387
+ 4.48e+10Hz 0.93055 -0.340111
+ 4.49e+10Hz 0.930282 -0.340835
+ 4.5e+10Hz 0.930014 -0.341559
+ 4.51e+10Hz 0.929744 -0.342282
+ 4.52e+10Hz 0.929475 -0.343006
+ 4.53e+10Hz 0.929204 -0.343729
+ 4.54e+10Hz 0.928933 -0.344452
+ 4.55e+10Hz 0.928662 -0.345175
+ 4.56e+10Hz 0.928389 -0.345897
+ 4.57e+10Hz 0.928116 -0.34662
+ 4.58e+10Hz 0.927843 -0.347342
+ 4.59e+10Hz 0.927568 -0.348064
+ 4.6e+10Hz 0.927293 -0.348786
+ 4.61e+10Hz 0.927018 -0.349507
+ 4.62e+10Hz 0.926742 -0.350229
+ 4.63e+10Hz 0.926465 -0.35095
+ 4.64e+10Hz 0.926187 -0.351671
+ 4.65e+10Hz 0.925909 -0.352391
+ 4.66e+10Hz 0.92563 -0.353112
+ 4.67e+10Hz 0.925351 -0.353832
+ 4.68e+10Hz 0.925071 -0.354552
+ 4.69e+10Hz 0.92479 -0.355272
+ 4.7e+10Hz 0.924509 -0.355992
+ 4.71e+10Hz 0.924227 -0.356711
+ 4.72e+10Hz 0.923944 -0.35743
+ 4.73e+10Hz 0.923661 -0.358149
+ 4.74e+10Hz 0.923377 -0.358867
+ 4.75e+10Hz 0.923092 -0.359586
+ 4.76e+10Hz 0.922807 -0.360304
+ 4.77e+10Hz 0.922521 -0.361022
+ 4.78e+10Hz 0.922235 -0.361739
+ 4.79e+10Hz 0.921948 -0.362457
+ 4.8e+10Hz 0.92166 -0.363174
+ 4.81e+10Hz 0.921371 -0.36389
+ 4.82e+10Hz 0.921082 -0.364607
+ 4.83e+10Hz 0.920793 -0.365323
+ 4.84e+10Hz 0.920503 -0.366039
+ 4.85e+10Hz 0.920212 -0.366755
+ 4.86e+10Hz 0.91992 -0.36747
+ 4.87e+10Hz 0.919628 -0.368185
+ 4.88e+10Hz 0.919335 -0.3689
+ 4.89e+10Hz 0.919042 -0.369615
+ 4.9e+10Hz 0.918748 -0.370329
+ 4.91e+10Hz 0.918454 -0.371043
+ 4.92e+10Hz 0.918158 -0.371756
+ 4.93e+10Hz 0.917863 -0.37247
+ 4.94e+10Hz 0.917566 -0.373183
+ 4.95e+10Hz 0.917269 -0.373896
+ 4.96e+10Hz 0.916972 -0.374608
+ 4.97e+10Hz 0.916673 -0.37532
+ 4.98e+10Hz 0.916375 -0.376032
+ 4.99e+10Hz 0.916075 -0.376744
+ 5e+10Hz 0.915775 -0.377455
+ 5.01e+10Hz 0.915475 -0.378166
+ 5.02e+10Hz 0.915174 -0.378877
+ 5.03e+10Hz 0.914872 -0.379587
+ 5.04e+10Hz 0.914569 -0.380297
+ 5.05e+10Hz 0.914267 -0.381007
+ 5.06e+10Hz 0.913963 -0.381716
+ 5.07e+10Hz 0.913659 -0.382425
+ 5.08e+10Hz 0.913354 -0.383134
+ 5.09e+10Hz 0.913049 -0.383842
+ 5.1e+10Hz 0.912743 -0.38455
+ 5.11e+10Hz 0.912437 -0.385258
+ 5.12e+10Hz 0.91213 -0.385966
+ 5.13e+10Hz 0.911823 -0.386673
+ 5.14e+10Hz 0.911515 -0.38738
+ 5.15e+10Hz 0.911206 -0.388086
+ 5.16e+10Hz 0.910897 -0.388792
+ 5.17e+10Hz 0.910587 -0.389498
+ 5.18e+10Hz 0.910277 -0.390204
+ 5.19e+10Hz 0.909967 -0.390909
+ 5.2e+10Hz 0.909655 -0.391614
+ 5.21e+10Hz 0.909343 -0.392318
+ 5.22e+10Hz 0.909031 -0.393023
+ 5.23e+10Hz 0.908718 -0.393726
+ 5.24e+10Hz 0.908405 -0.39443
+ 5.25e+10Hz 0.908091 -0.395133
+ 5.26e+10Hz 0.907776 -0.395836
+ 5.27e+10Hz 0.907461 -0.396539
+ 5.28e+10Hz 0.907146 -0.397241
+ 5.29e+10Hz 0.90683 -0.397943
+ 5.3e+10Hz 0.906513 -0.398645
+ 5.31e+10Hz 0.906196 -0.399346
+ 5.32e+10Hz 0.905878 -0.400047
+ 5.33e+10Hz 0.90556 -0.400748
+ 5.34e+10Hz 0.905242 -0.401448
+ 5.35e+10Hz 0.904922 -0.402148
+ 5.36e+10Hz 0.904603 -0.402848
+ 5.37e+10Hz 0.904283 -0.403547
+ 5.38e+10Hz 0.903962 -0.404246
+ 5.39e+10Hz 0.903641 -0.404945
+ 5.4e+10Hz 0.903319 -0.405643
+ 5.41e+10Hz 0.902997 -0.406341
+ 5.42e+10Hz 0.902675 -0.407039
+ 5.43e+10Hz 0.902351 -0.407737
+ 5.44e+10Hz 0.902028 -0.408434
+ 5.45e+10Hz 0.901704 -0.409131
+ 5.46e+10Hz 0.901379 -0.409827
+ 5.47e+10Hz 0.901054 -0.410523
+ 5.48e+10Hz 0.900729 -0.411219
+ 5.49e+10Hz 0.900403 -0.411915
+ 5.5e+10Hz 0.900076 -0.41261
+ 5.51e+10Hz 0.899749 -0.413305
+ 5.52e+10Hz 0.899422 -0.414
+ 5.53e+10Hz 0.899094 -0.414694
+ 5.54e+10Hz 0.898765 -0.415388
+ 5.55e+10Hz 0.898437 -0.416082
+ 5.56e+10Hz 0.898107 -0.416776
+ 5.57e+10Hz 0.897778 -0.417469
+ 5.58e+10Hz 0.897447 -0.418162
+ 5.59e+10Hz 0.897117 -0.418854
+ 5.6e+10Hz 0.896785 -0.419547
+ 5.61e+10Hz 0.896454 -0.420239
+ 5.62e+10Hz 0.896122 -0.420931
+ 5.63e+10Hz 0.895789 -0.421622
+ 5.64e+10Hz 0.895456 -0.422313
+ 5.65e+10Hz 0.895122 -0.423004
+ 5.66e+10Hz 0.894788 -0.423695
+ 5.67e+10Hz 0.894454 -0.424385
+ 5.68e+10Hz 0.894119 -0.425075
+ 5.69e+10Hz 0.893784 -0.425765
+ 5.7e+10Hz 0.893448 -0.426455
+ 5.71e+10Hz 0.893112 -0.427144
+ 5.72e+10Hz 0.892775 -0.427833
+ 5.73e+10Hz 0.892438 -0.428522
+ 5.74e+10Hz 0.8921 -0.42921
+ 5.75e+10Hz 0.891762 -0.429898
+ 5.76e+10Hz 0.891424 -0.430586
+ 5.77e+10Hz 0.891085 -0.431274
+ 5.78e+10Hz 0.890745 -0.431961
+ 5.79e+10Hz 0.890405 -0.432648
+ 5.8e+10Hz 0.890065 -0.433335
+ 5.81e+10Hz 0.889724 -0.434022
+ 5.82e+10Hz 0.889383 -0.434708
+ 5.83e+10Hz 0.889041 -0.435394
+ 5.84e+10Hz 0.888699 -0.43608
+ 5.85e+10Hz 0.888356 -0.436766
+ 5.86e+10Hz 0.888013 -0.437451
+ 5.87e+10Hz 0.887669 -0.438137
+ 5.88e+10Hz 0.887325 -0.438821
+ 5.89e+10Hz 0.886981 -0.439506
+ 5.9e+10Hz 0.886636 -0.440191
+ 5.91e+10Hz 0.88629 -0.440875
+ 5.92e+10Hz 0.885944 -0.441559
+ 5.93e+10Hz 0.885598 -0.442242
+ 5.94e+10Hz 0.885251 -0.442926
+ 5.95e+10Hz 0.884904 -0.443609
+ 5.96e+10Hz 0.884556 -0.444292
+ 5.97e+10Hz 0.884208 -0.444975
+ 5.98e+10Hz 0.883859 -0.445658
+ 5.99e+10Hz 0.88351 -0.44634
+ 6e+10Hz 0.88316 -0.447022
+ 6.01e+10Hz 0.88281 -0.447704
+ 6.02e+10Hz 0.88246 -0.448385
+ 6.03e+10Hz 0.882108 -0.449067
+ 6.04e+10Hz 0.881757 -0.449748
+ 6.05e+10Hz 0.881405 -0.450429
+ 6.06e+10Hz 0.881052 -0.45111
+ 6.07e+10Hz 0.880699 -0.45179
+ 6.08e+10Hz 0.880346 -0.452471
+ 6.09e+10Hz 0.879992 -0.453151
+ 6.1e+10Hz 0.879637 -0.453831
+ 6.11e+10Hz 0.879282 -0.45451
+ 6.12e+10Hz 0.878927 -0.45519
+ 6.13e+10Hz 0.878571 -0.455869
+ 6.14e+10Hz 0.878215 -0.456548
+ 6.15e+10Hz 0.877858 -0.457227
+ 6.16e+10Hz 0.8775 -0.457905
+ 6.17e+10Hz 0.877142 -0.458584
+ 6.18e+10Hz 0.876784 -0.459262
+ 6.19e+10Hz 0.876425 -0.45994
+ 6.2e+10Hz 0.876066 -0.460618
+ 6.21e+10Hz 0.875706 -0.461295
+ 6.22e+10Hz 0.875345 -0.461972
+ 6.23e+10Hz 0.874984 -0.462649
+ 6.24e+10Hz 0.874623 -0.463326
+ 6.25e+10Hz 0.874261 -0.464003
+ 6.26e+10Hz 0.873899 -0.464679
+ 6.27e+10Hz 0.873536 -0.465356
+ 6.28e+10Hz 0.873172 -0.466032
+ 6.29e+10Hz 0.872808 -0.466707
+ 6.3e+10Hz 0.872444 -0.467383
+ 6.31e+10Hz 0.872079 -0.468058
+ 6.32e+10Hz 0.871713 -0.468734
+ 6.33e+10Hz 0.871347 -0.469408
+ 6.34e+10Hz 0.87098 -0.470083
+ 6.35e+10Hz 0.870613 -0.470758
+ 6.36e+10Hz 0.870245 -0.471432
+ 6.37e+10Hz 0.869877 -0.472106
+ 6.38e+10Hz 0.869508 -0.47278
+ 6.39e+10Hz 0.869139 -0.473453
+ 6.4e+10Hz 0.868769 -0.474127
+ 6.41e+10Hz 0.868399 -0.4748
+ 6.42e+10Hz 0.868028 -0.475473
+ 6.43e+10Hz 0.867657 -0.476145
+ 6.44e+10Hz 0.867285 -0.476818
+ 6.45e+10Hz 0.866912 -0.47749
+ 6.46e+10Hz 0.866539 -0.478162
+ 6.47e+10Hz 0.866165 -0.478834
+ 6.48e+10Hz 0.865791 -0.479506
+ 6.49e+10Hz 0.865416 -0.480177
+ 6.5e+10Hz 0.865041 -0.480848
+ 6.51e+10Hz 0.864665 -0.481519
+ 6.52e+10Hz 0.864289 -0.482189
+ 6.53e+10Hz 0.863912 -0.48286
+ 6.54e+10Hz 0.863534 -0.48353
+ 6.55e+10Hz 0.863156 -0.4842
+ 6.56e+10Hz 0.862778 -0.484869
+ 6.57e+10Hz 0.862399 -0.485539
+ 6.58e+10Hz 0.862019 -0.486208
+ 6.59e+10Hz 0.861639 -0.486877
+ 6.6e+10Hz 0.861258 -0.487546
+ 6.61e+10Hz 0.860876 -0.488214
+ 6.62e+10Hz 0.860494 -0.488882
+ 6.63e+10Hz 0.860112 -0.48955
+ 6.64e+10Hz 0.859729 -0.490218
+ 6.65e+10Hz 0.859345 -0.490885
+ 6.66e+10Hz 0.858961 -0.491552
+ 6.67e+10Hz 0.858576 -0.492219
+ 6.68e+10Hz 0.85819 -0.492886
+ 6.69e+10Hz 0.857804 -0.493552
+ 6.7e+10Hz 0.857418 -0.494218
+ 6.71e+10Hz 0.857031 -0.494884
+ 6.72e+10Hz 0.856643 -0.495549
+ 6.73e+10Hz 0.856255 -0.496214
+ 6.74e+10Hz 0.855866 -0.496879
+ 6.75e+10Hz 0.855476 -0.497544
+ 6.76e+10Hz 0.855086 -0.498208
+ 6.77e+10Hz 0.854696 -0.498872
+ 6.78e+10Hz 0.854305 -0.499536
+ 6.79e+10Hz 0.853913 -0.5002
+ 6.8e+10Hz 0.853521 -0.500863
+ 6.81e+10Hz 0.853128 -0.501526
+ 6.82e+10Hz 0.852734 -0.502189
+ 6.83e+10Hz 0.85234 -0.502851
+ 6.84e+10Hz 0.851946 -0.503513
+ 6.85e+10Hz 0.851551 -0.504175
+ 6.86e+10Hz 0.851155 -0.504836
+ 6.87e+10Hz 0.850759 -0.505497
+ 6.88e+10Hz 0.850362 -0.506158
+ 6.89e+10Hz 0.849964 -0.506819
+ 6.9e+10Hz 0.849566 -0.507479
+ 6.91e+10Hz 0.849168 -0.508139
+ 6.92e+10Hz 0.848768 -0.508798
+ 6.93e+10Hz 0.848369 -0.509457
+ 6.94e+10Hz 0.847968 -0.510116
+ 6.95e+10Hz 0.847567 -0.510775
+ 6.96e+10Hz 0.847166 -0.511433
+ 6.97e+10Hz 0.846764 -0.512091
+ 6.98e+10Hz 0.846361 -0.512749
+ 6.99e+10Hz 0.845958 -0.513406
+ 7e+10Hz 0.845554 -0.514063
+ 7.01e+10Hz 0.84515 -0.51472
+ 7.02e+10Hz 0.844745 -0.515376
+ 7.03e+10Hz 0.84434 -0.516032
+ 7.04e+10Hz 0.843934 -0.516687
+ 7.05e+10Hz 0.843527 -0.517343
+ 7.06e+10Hz 0.84312 -0.517998
+ 7.07e+10Hz 0.842712 -0.518652
+ 7.08e+10Hz 0.842304 -0.519306
+ 7.09e+10Hz 0.841895 -0.51996
+ 7.1e+10Hz 0.841486 -0.520614
+ 7.11e+10Hz 0.841076 -0.521267
+ 7.12e+10Hz 0.840665 -0.52192
+ 7.13e+10Hz 0.840254 -0.522572
+ 7.14e+10Hz 0.839843 -0.523224
+ 7.15e+10Hz 0.83943 -0.523876
+ 7.16e+10Hz 0.839018 -0.524527
+ 7.17e+10Hz 0.838605 -0.525178
+ 7.18e+10Hz 0.838191 -0.525829
+ 7.19e+10Hz 0.837776 -0.526479
+ 7.2e+10Hz 0.837362 -0.527129
+ 7.21e+10Hz 0.836946 -0.527779
+ 7.22e+10Hz 0.83653 -0.528428
+ 7.23e+10Hz 0.836114 -0.529077
+ 7.24e+10Hz 0.835697 -0.529725
+ 7.25e+10Hz 0.835279 -0.530373
+ 7.26e+10Hz 0.834861 -0.531021
+ 7.27e+10Hz 0.834442 -0.531668
+ 7.28e+10Hz 0.834023 -0.532315
+ 7.29e+10Hz 0.833604 -0.532961
+ 7.3e+10Hz 0.833183 -0.533608
+ 7.31e+10Hz 0.832763 -0.534253
+ 7.32e+10Hz 0.832341 -0.534899
+ 7.33e+10Hz 0.83192 -0.535544
+ 7.34e+10Hz 0.831497 -0.536188
+ 7.35e+10Hz 0.831075 -0.536833
+ 7.36e+10Hz 0.830651 -0.537476
+ 7.37e+10Hz 0.830227 -0.53812
+ 7.38e+10Hz 0.829803 -0.538763
+ 7.39e+10Hz 0.829378 -0.539406
+ 7.4e+10Hz 0.828953 -0.540048
+ 7.41e+10Hz 0.828527 -0.54069
+ 7.42e+10Hz 0.828101 -0.541331
+ 7.43e+10Hz 0.827674 -0.541972
+ 7.44e+10Hz 0.827246 -0.542613
+ 7.45e+10Hz 0.826818 -0.543254
+ 7.46e+10Hz 0.82639 -0.543894
+ 7.47e+10Hz 0.825961 -0.544533
+ 7.48e+10Hz 0.825532 -0.545172
+ 7.49e+10Hz 0.825102 -0.545811
+ 7.5e+10Hz 0.824672 -0.546449
+ 7.51e+10Hz 0.824241 -0.547087
+ 7.52e+10Hz 0.82381 -0.547725
+ 7.53e+10Hz 0.823378 -0.548362
+ 7.54e+10Hz 0.822946 -0.548999
+ 7.55e+10Hz 0.822513 -0.549636
+ 7.56e+10Hz 0.82208 -0.550272
+ 7.57e+10Hz 0.821646 -0.550907
+ 7.58e+10Hz 0.821212 -0.551542
+ 7.59e+10Hz 0.820777 -0.552177
+ 7.6e+10Hz 0.820342 -0.552812
+ 7.61e+10Hz 0.819906 -0.553446
+ 7.62e+10Hz 0.81947 -0.55408
+ 7.63e+10Hz 0.819034 -0.554713
+ 7.64e+10Hz 0.818597 -0.555346
+ 7.65e+10Hz 0.818159 -0.555978
+ 7.66e+10Hz 0.817721 -0.556611
+ 7.67e+10Hz 0.817283 -0.557242
+ 7.68e+10Hz 0.816844 -0.557874
+ 7.69e+10Hz 0.816405 -0.558505
+ 7.7e+10Hz 0.815965 -0.559135
+ 7.71e+10Hz 0.815525 -0.559765
+ 7.72e+10Hz 0.815084 -0.560395
+ 7.73e+10Hz 0.814643 -0.561025
+ 7.74e+10Hz 0.814202 -0.561654
+ 7.75e+10Hz 0.81376 -0.562282
+ 7.76e+10Hz 0.813317 -0.562911
+ 7.77e+10Hz 0.812874 -0.563539
+ 7.78e+10Hz 0.812431 -0.564166
+ 7.79e+10Hz 0.811987 -0.564793
+ 7.8e+10Hz 0.811543 -0.56542
+ 7.81e+10Hz 0.811098 -0.566047
+ 7.82e+10Hz 0.810653 -0.566673
+ 7.83e+10Hz 0.810208 -0.567298
+ 7.84e+10Hz 0.809762 -0.567924
+ 7.85e+10Hz 0.809315 -0.568549
+ 7.86e+10Hz 0.808868 -0.569173
+ 7.87e+10Hz 0.808421 -0.569797
+ 7.88e+10Hz 0.807973 -0.570421
+ 7.89e+10Hz 0.807525 -0.571044
+ 7.9e+10Hz 0.807076 -0.571668
+ 7.91e+10Hz 0.806627 -0.57229
+ 7.92e+10Hz 0.806178 -0.572913
+ 7.93e+10Hz 0.805728 -0.573535
+ 7.94e+10Hz 0.805278 -0.574156
+ 7.95e+10Hz 0.804827 -0.574777
+ 7.96e+10Hz 0.804376 -0.575398
+ 7.97e+10Hz 0.803924 -0.576019
+ 7.98e+10Hz 0.803472 -0.576639
+ 7.99e+10Hz 0.80302 -0.577259
+ 8e+10Hz 0.802567 -0.577878
+ 8.01e+10Hz 0.802113 -0.578497
+ 8.02e+10Hz 0.80166 -0.579116
+ 8.03e+10Hz 0.801205 -0.579734
+ 8.04e+10Hz 0.800751 -0.580352
+ 8.05e+10Hz 0.800296 -0.58097
+ 8.06e+10Hz 0.79984 -0.581587
+ 8.07e+10Hz 0.799384 -0.582204
+ 8.08e+10Hz 0.798928 -0.582821
+ 8.09e+10Hz 0.798471 -0.583437
+ 8.1e+10Hz 0.798014 -0.584053
+ 8.11e+10Hz 0.797556 -0.584669
+ 8.12e+10Hz 0.797098 -0.585284
+ 8.13e+10Hz 0.79664 -0.585899
+ 8.14e+10Hz 0.796181 -0.586514
+ 8.15e+10Hz 0.795721 -0.587128
+ 8.16e+10Hz 0.795262 -0.587742
+ 8.17e+10Hz 0.794801 -0.588355
+ 8.18e+10Hz 0.794341 -0.588969
+ 8.19e+10Hz 0.79388 -0.589581
+ 8.2e+10Hz 0.793418 -0.590194
+ 8.21e+10Hz 0.792956 -0.590806
+ 8.22e+10Hz 0.792494 -0.591418
+ 8.23e+10Hz 0.792031 -0.59203
+ 8.24e+10Hz 0.791568 -0.592641
+ 8.25e+10Hz 0.791104 -0.593252
+ 8.26e+10Hz 0.79064 -0.593862
+ 8.27e+10Hz 0.790176 -0.594472
+ 8.28e+10Hz 0.789711 -0.595082
+ 8.29e+10Hz 0.789245 -0.595692
+ 8.3e+10Hz 0.788779 -0.596301
+ 8.31e+10Hz 0.788313 -0.59691
+ 8.32e+10Hz 0.787846 -0.597518
+ 8.33e+10Hz 0.787379 -0.598127
+ 8.34e+10Hz 0.786912 -0.598735
+ 8.35e+10Hz 0.786444 -0.599342
+ 8.36e+10Hz 0.785975 -0.599949
+ 8.37e+10Hz 0.785506 -0.600556
+ 8.38e+10Hz 0.785037 -0.601163
+ 8.39e+10Hz 0.784567 -0.601769
+ 8.4e+10Hz 0.784097 -0.602375
+ 8.41e+10Hz 0.783626 -0.602981
+ 8.42e+10Hz 0.783155 -0.603586
+ 8.43e+10Hz 0.782683 -0.604191
+ 8.44e+10Hz 0.782211 -0.604796
+ 8.45e+10Hz 0.781739 -0.6054
+ 8.46e+10Hz 0.781266 -0.606004
+ 8.47e+10Hz 0.780792 -0.606608
+ 8.48e+10Hz 0.780319 -0.607211
+ 8.49e+10Hz 0.779844 -0.607814
+ 8.5e+10Hz 0.779369 -0.608417
+ 8.51e+10Hz 0.778894 -0.609019
+ 8.52e+10Hz 0.778419 -0.609621
+ 8.53e+10Hz 0.777942 -0.610223
+ 8.54e+10Hz 0.777466 -0.610825
+ 8.55e+10Hz 0.776989 -0.611426
+ 8.56e+10Hz 0.776511 -0.612026
+ 8.57e+10Hz 0.776033 -0.612627
+ 8.58e+10Hz 0.775555 -0.613227
+ 8.59e+10Hz 0.775076 -0.613827
+ 8.6e+10Hz 0.774596 -0.614426
+ 8.61e+10Hz 0.774117 -0.615025
+ 8.62e+10Hz 0.773636 -0.615624
+ 8.63e+10Hz 0.773155 -0.616223
+ 8.64e+10Hz 0.772674 -0.616821
+ 8.65e+10Hz 0.772192 -0.617419
+ 8.66e+10Hz 0.77171 -0.618016
+ 8.67e+10Hz 0.771228 -0.618614
+ 8.68e+10Hz 0.770744 -0.61921
+ 8.69e+10Hz 0.770261 -0.619807
+ 8.7e+10Hz 0.769777 -0.620403
+ 8.71e+10Hz 0.769292 -0.620999
+ 8.72e+10Hz 0.768807 -0.621594
+ 8.73e+10Hz 0.768321 -0.62219
+ 8.74e+10Hz 0.767835 -0.622784
+ 8.75e+10Hz 0.767349 -0.623379
+ 8.76e+10Hz 0.766862 -0.623973
+ 8.77e+10Hz 0.766374 -0.624567
+ 8.78e+10Hz 0.765886 -0.625161
+ 8.79e+10Hz 0.765398 -0.625754
+ 8.8e+10Hz 0.764909 -0.626346
+ 8.81e+10Hz 0.76442 -0.626939
+ 8.82e+10Hz 0.76393 -0.627531
+ 8.83e+10Hz 0.763439 -0.628123
+ 8.84e+10Hz 0.762948 -0.628714
+ 8.85e+10Hz 0.762457 -0.629305
+ 8.86e+10Hz 0.761965 -0.629896
+ 8.87e+10Hz 0.761473 -0.630487
+ 8.88e+10Hz 0.76098 -0.631077
+ 8.89e+10Hz 0.760487 -0.631666
+ 8.9e+10Hz 0.759993 -0.632256
+ 8.91e+10Hz 0.759499 -0.632845
+ 8.92e+10Hz 0.759004 -0.633433
+ 8.93e+10Hz 0.758508 -0.634021
+ 8.94e+10Hz 0.758013 -0.634609
+ 8.95e+10Hz 0.757516 -0.635197
+ 8.96e+10Hz 0.757019 -0.635784
+ 8.97e+10Hz 0.756522 -0.636371
+ 8.98e+10Hz 0.756024 -0.636957
+ 8.99e+10Hz 0.755526 -0.637543
+ 9e+10Hz 0.755027 -0.638129
+ 9.01e+10Hz 0.754528 -0.638715
+ 9.02e+10Hz 0.754028 -0.639299
+ 9.03e+10Hz 0.753528 -0.639884
+ 9.04e+10Hz 0.753027 -0.640468
+ 9.05e+10Hz 0.752526 -0.641052
+ 9.06e+10Hz 0.752024 -0.641636
+ 9.07e+10Hz 0.751522 -0.642219
+ 9.08e+10Hz 0.751019 -0.642801
+ 9.09e+10Hz 0.750516 -0.643384
+ 9.1e+10Hz 0.750012 -0.643966
+ 9.11e+10Hz 0.749508 -0.644547
+ 9.12e+10Hz 0.749003 -0.645128
+ 9.13e+10Hz 0.748498 -0.645709
+ 9.14e+10Hz 0.747992 -0.64629
+ 9.15e+10Hz 0.747486 -0.64687
+ 9.16e+10Hz 0.74698 -0.647449
+ 9.17e+10Hz 0.746472 -0.648028
+ 9.18e+10Hz 0.745965 -0.648607
+ 9.19e+10Hz 0.745456 -0.649186
+ 9.2e+10Hz 0.744948 -0.649764
+ 9.21e+10Hz 0.744439 -0.650341
+ 9.22e+10Hz 0.743929 -0.650919
+ 9.23e+10Hz 0.743419 -0.651495
+ 9.24e+10Hz 0.742908 -0.652072
+ 9.25e+10Hz 0.742397 -0.652648
+ 9.26e+10Hz 0.741885 -0.653223
+ 9.27e+10Hz 0.741373 -0.653799
+ 9.28e+10Hz 0.740861 -0.654373
+ 9.29e+10Hz 0.740347 -0.654948
+ 9.3e+10Hz 0.739834 -0.655522
+ 9.31e+10Hz 0.73932 -0.656095
+ 9.32e+10Hz 0.738805 -0.656668
+ 9.33e+10Hz 0.73829 -0.657241
+ 9.34e+10Hz 0.737775 -0.657813
+ 9.35e+10Hz 0.737259 -0.658385
+ 9.36e+10Hz 0.736742 -0.658956
+ 9.37e+10Hz 0.736225 -0.659527
+ 9.38e+10Hz 0.735708 -0.660098
+ 9.39e+10Hz 0.73519 -0.660668
+ 9.4e+10Hz 0.734671 -0.661238
+ 9.41e+10Hz 0.734153 -0.661807
+ 9.42e+10Hz 0.733633 -0.662376
+ 9.43e+10Hz 0.733113 -0.662944
+ 9.44e+10Hz 0.732593 -0.663512
+ 9.45e+10Hz 0.732072 -0.66408
+ 9.46e+10Hz 0.731551 -0.664647
+ 9.47e+10Hz 0.731029 -0.665214
+ 9.48e+10Hz 0.730507 -0.66578
+ 9.49e+10Hz 0.729984 -0.666346
+ 9.5e+10Hz 0.729461 -0.666911
+ 9.51e+10Hz 0.728938 -0.667476
+ 9.52e+10Hz 0.728414 -0.66804
+ 9.53e+10Hz 0.727889 -0.668605
+ 9.54e+10Hz 0.727364 -0.669168
+ 9.55e+10Hz 0.726839 -0.669731
+ 9.56e+10Hz 0.726313 -0.670294
+ 9.57e+10Hz 0.725787 -0.670856
+ 9.58e+10Hz 0.72526 -0.671418
+ 9.59e+10Hz 0.724733 -0.671979
+ 9.6e+10Hz 0.724205 -0.67254
+ 9.61e+10Hz 0.723677 -0.673101
+ 9.62e+10Hz 0.723148 -0.673661
+ 9.63e+10Hz 0.722619 -0.67422
+ 9.64e+10Hz 0.72209 -0.674779
+ 9.65e+10Hz 0.72156 -0.675338
+ 9.66e+10Hz 0.721029 -0.675896
+ 9.67e+10Hz 0.720498 -0.676454
+ 9.68e+10Hz 0.719967 -0.677011
+ 9.69e+10Hz 0.719436 -0.677568
+ 9.7e+10Hz 0.718903 -0.678125
+ 9.71e+10Hz 0.718371 -0.678681
+ 9.72e+10Hz 0.717838 -0.679236
+ 9.73e+10Hz 0.717304 -0.679791
+ 9.74e+10Hz 0.71677 -0.680346
+ 9.75e+10Hz 0.716236 -0.6809
+ 9.76e+10Hz 0.715701 -0.681453
+ 9.77e+10Hz 0.715166 -0.682007
+ 9.78e+10Hz 0.714631 -0.682559
+ 9.79e+10Hz 0.714095 -0.683112
+ 9.8e+10Hz 0.713558 -0.683664
+ 9.81e+10Hz 0.713021 -0.684215
+ 9.82e+10Hz 0.712484 -0.684766
+ 9.83e+10Hz 0.711946 -0.685316
+ 9.84e+10Hz 0.711408 -0.685866
+ 9.85e+10Hz 0.71087 -0.686416
+ 9.86e+10Hz 0.710331 -0.686965
+ 9.87e+10Hz 0.709791 -0.687514
+ 9.88e+10Hz 0.709252 -0.688062
+ 9.89e+10Hz 0.708712 -0.68861
+ 9.9e+10Hz 0.708171 -0.689157
+ 9.91e+10Hz 0.70763 -0.689704
+ 9.92e+10Hz 0.707089 -0.69025
+ 9.93e+10Hz 0.706547 -0.690796
+ 9.94e+10Hz 0.706004 -0.691342
+ 9.95e+10Hz 0.705462 -0.691887
+ 9.96e+10Hz 0.704919 -0.692431
+ 9.97e+10Hz 0.704375 -0.692975
+ 9.98e+10Hz 0.703832 -0.693519
+ 9.99e+10Hz 0.703287 -0.694062
+ 1e+11Hz 0.702743 -0.694605
+ 1.001e+11Hz 0.702198 -0.695147
+ 1.002e+11Hz 0.701652 -0.695689
+ 1.003e+11Hz 0.701106 -0.696231
+ 1.004e+11Hz 0.70056 -0.696772
+ 1.005e+11Hz 0.700014 -0.697312
+ 1.006e+11Hz 0.699467 -0.697852
+ 1.007e+11Hz 0.698919 -0.698392
+ 1.008e+11Hz 0.698372 -0.698931
+ 1.009e+11Hz 0.697823 -0.69947
+ 1.01e+11Hz 0.697275 -0.700008
+ 1.011e+11Hz 0.696726 -0.700546
+ 1.012e+11Hz 0.696177 -0.701083
+ 1.013e+11Hz 0.695627 -0.70162
+ 1.014e+11Hz 0.695077 -0.702157
+ 1.015e+11Hz 0.694526 -0.702693
+ 1.016e+11Hz 0.693975 -0.703229
+ 1.017e+11Hz 0.693424 -0.703764
+ 1.018e+11Hz 0.692873 -0.704299
+ 1.019e+11Hz 0.692321 -0.704833
+ 1.02e+11Hz 0.691768 -0.705367
+ 1.021e+11Hz 0.691215 -0.7059
+ 1.022e+11Hz 0.690662 -0.706433
+ 1.023e+11Hz 0.690109 -0.706966
+ 1.024e+11Hz 0.689555 -0.707498
+ 1.025e+11Hz 0.689 -0.70803
+ 1.026e+11Hz 0.688446 -0.708561
+ 1.027e+11Hz 0.687891 -0.709092
+ 1.028e+11Hz 0.687335 -0.709622
+ 1.029e+11Hz 0.686779 -0.710152
+ 1.03e+11Hz 0.686223 -0.710682
+ 1.031e+11Hz 0.685667 -0.711211
+ 1.032e+11Hz 0.68511 -0.71174
+ 1.033e+11Hz 0.684552 -0.712268
+ 1.034e+11Hz 0.683995 -0.712796
+ 1.035e+11Hz 0.683437 -0.713323
+ 1.036e+11Hz 0.682878 -0.71385
+ 1.037e+11Hz 0.682319 -0.714377
+ 1.038e+11Hz 0.68176 -0.714903
+ 1.039e+11Hz 0.681201 -0.715428
+ 1.04e+11Hz 0.680641 -0.715954
+ 1.041e+11Hz 0.68008 -0.716479
+ 1.042e+11Hz 0.67952 -0.717003
+ 1.043e+11Hz 0.678958 -0.717527
+ 1.044e+11Hz 0.678397 -0.718051
+ 1.045e+11Hz 0.677835 -0.718574
+ 1.046e+11Hz 0.677273 -0.719097
+ 1.047e+11Hz 0.67671 -0.719619
+ 1.048e+11Hz 0.676147 -0.720141
+ 1.049e+11Hz 0.675584 -0.720662
+ 1.05e+11Hz 0.67502 -0.721183
+ 1.051e+11Hz 0.674456 -0.721704
+ 1.052e+11Hz 0.673891 -0.722224
+ 1.053e+11Hz 0.673327 -0.722744
+ 1.054e+11Hz 0.672761 -0.723264
+ 1.055e+11Hz 0.672196 -0.723783
+ 1.056e+11Hz 0.67163 -0.724301
+ 1.057e+11Hz 0.671063 -0.72482
+ 1.058e+11Hz 0.670496 -0.725337
+ 1.059e+11Hz 0.669929 -0.725855
+ 1.06e+11Hz 0.669362 -0.726372
+ 1.061e+11Hz 0.668794 -0.726888
+ 1.062e+11Hz 0.668225 -0.727404
+ 1.063e+11Hz 0.667657 -0.72792
+ 1.064e+11Hz 0.667087 -0.728435
+ 1.065e+11Hz 0.666518 -0.72895
+ 1.066e+11Hz 0.665948 -0.729465
+ 1.067e+11Hz 0.665378 -0.729979
+ 1.068e+11Hz 0.664807 -0.730493
+ 1.069e+11Hz 0.664236 -0.731006
+ 1.07e+11Hz 0.663665 -0.731519
+ 1.071e+11Hz 0.663093 -0.732031
+ 1.072e+11Hz 0.662521 -0.732543
+ 1.073e+11Hz 0.661948 -0.733055
+ 1.074e+11Hz 0.661375 -0.733566
+ 1.075e+11Hz 0.660801 -0.734077
+ 1.076e+11Hz 0.660228 -0.734587
+ 1.077e+11Hz 0.659653 -0.735097
+ 1.078e+11Hz 0.659079 -0.735607
+ 1.079e+11Hz 0.658504 -0.736116
+ 1.08e+11Hz 0.657928 -0.736625
+ 1.081e+11Hz 0.657353 -0.737133
+ 1.082e+11Hz 0.656776 -0.737641
+ 1.083e+11Hz 0.6562 -0.738148
+ 1.084e+11Hz 0.655623 -0.738655
+ 1.085e+11Hz 0.655045 -0.739162
+ 1.086e+11Hz 0.654468 -0.739668
+ 1.087e+11Hz 0.653889 -0.740174
+ 1.088e+11Hz 0.653311 -0.74068
+ 1.089e+11Hz 0.652732 -0.741185
+ 1.09e+11Hz 0.652152 -0.741689
+ 1.091e+11Hz 0.651573 -0.742194
+ 1.092e+11Hz 0.650992 -0.742697
+ 1.093e+11Hz 0.650412 -0.743201
+ 1.094e+11Hz 0.649831 -0.743704
+ 1.095e+11Hz 0.649249 -0.744206
+ 1.096e+11Hz 0.648667 -0.744708
+ 1.097e+11Hz 0.648085 -0.74521
+ 1.098e+11Hz 0.647502 -0.745711
+ 1.099e+11Hz 0.646919 -0.746212
+ 1.1e+11Hz 0.646336 -0.746713
+ 1.101e+11Hz 0.645752 -0.747213
+ 1.102e+11Hz 0.645167 -0.747712
+ 1.103e+11Hz 0.644583 -0.748212
+ 1.104e+11Hz 0.643998 -0.74871
+ 1.105e+11Hz 0.643412 -0.749209
+ 1.106e+11Hz 0.642826 -0.749706
+ 1.107e+11Hz 0.64224 -0.750204
+ 1.108e+11Hz 0.641653 -0.750701
+ 1.109e+11Hz 0.641065 -0.751198
+ 1.11e+11Hz 0.640478 -0.751694
+ 1.111e+11Hz 0.63989 -0.75219
+ 1.112e+11Hz 0.639301 -0.752685
+ 1.113e+11Hz 0.638712 -0.75318
+ 1.114e+11Hz 0.638123 -0.753674
+ 1.115e+11Hz 0.637533 -0.754168
+ 1.116e+11Hz 0.636943 -0.754662
+ 1.117e+11Hz 0.636352 -0.755155
+ 1.118e+11Hz 0.635761 -0.755648
+ 1.119e+11Hz 0.63517 -0.75614
+ 1.12e+11Hz 0.634578 -0.756632
+ 1.121e+11Hz 0.633986 -0.757123
+ 1.122e+11Hz 0.633393 -0.757614
+ 1.123e+11Hz 0.6328 -0.758105
+ 1.124e+11Hz 0.632206 -0.758595
+ 1.125e+11Hz 0.631612 -0.759084
+ 1.126e+11Hz 0.631018 -0.759573
+ 1.127e+11Hz 0.630423 -0.760062
+ 1.128e+11Hz 0.629828 -0.76055
+ 1.129e+11Hz 0.629232 -0.761038
+ 1.13e+11Hz 0.628636 -0.761526
+ 1.131e+11Hz 0.628039 -0.762012
+ 1.132e+11Hz 0.627442 -0.762499
+ 1.133e+11Hz 0.626845 -0.762985
+ 1.134e+11Hz 0.626247 -0.76347
+ 1.135e+11Hz 0.625649 -0.763955
+ 1.136e+11Hz 0.62505 -0.76444
+ 1.137e+11Hz 0.624451 -0.764924
+ 1.138e+11Hz 0.623852 -0.765408
+ 1.139e+11Hz 0.623252 -0.765891
+ 1.14e+11Hz 0.622651 -0.766374
+ 1.141e+11Hz 0.622051 -0.766856
+ 1.142e+11Hz 0.621449 -0.767338
+ 1.143e+11Hz 0.620848 -0.767819
+ 1.144e+11Hz 0.620246 -0.7683
+ 1.145e+11Hz 0.619643 -0.76878
+ 1.146e+11Hz 0.61904 -0.76926
+ 1.147e+11Hz 0.618437 -0.76974
+ 1.148e+11Hz 0.617833 -0.770218
+ 1.149e+11Hz 0.617229 -0.770697
+ 1.15e+11Hz 0.616625 -0.771175
+ 1.151e+11Hz 0.61602 -0.771652
+ 1.152e+11Hz 0.615414 -0.772129
+ 1.153e+11Hz 0.614808 -0.772606
+ 1.154e+11Hz 0.614202 -0.773082
+ 1.155e+11Hz 0.613596 -0.773557
+ 1.156e+11Hz 0.612989 -0.774032
+ 1.157e+11Hz 0.612381 -0.774507
+ 1.158e+11Hz 0.611773 -0.774981
+ 1.159e+11Hz 0.611165 -0.775455
+ 1.16e+11Hz 0.610556 -0.775928
+ 1.161e+11Hz 0.609947 -0.7764
+ 1.162e+11Hz 0.609338 -0.776872
+ 1.163e+11Hz 0.608728 -0.777344
+ 1.164e+11Hz 0.608117 -0.777815
+ 1.165e+11Hz 0.607507 -0.778286
+ 1.166e+11Hz 0.606895 -0.778756
+ 1.167e+11Hz 0.606284 -0.779225
+ 1.168e+11Hz 0.605672 -0.779694
+ 1.169e+11Hz 0.60506 -0.780163
+ 1.17e+11Hz 0.604447 -0.780631
+ 1.171e+11Hz 0.603834 -0.781099
+ 1.172e+11Hz 0.60322 -0.781566
+ 1.173e+11Hz 0.602606 -0.782032
+ 1.174e+11Hz 0.601992 -0.782498
+ 1.175e+11Hz 0.601377 -0.782964
+ 1.176e+11Hz 0.600762 -0.783429
+ 1.177e+11Hz 0.600146 -0.783893
+ 1.178e+11Hz 0.59953 -0.784357
+ 1.179e+11Hz 0.598914 -0.784821
+ 1.18e+11Hz 0.598297 -0.785284
+ 1.181e+11Hz 0.59768 -0.785746
+ 1.182e+11Hz 0.597063 -0.786208
+ 1.183e+11Hz 0.596445 -0.786669
+ 1.184e+11Hz 0.595827 -0.78713
+ 1.185e+11Hz 0.595208 -0.78759
+ 1.186e+11Hz 0.594589 -0.78805
+ 1.187e+11Hz 0.593969 -0.78851
+ 1.188e+11Hz 0.59335 -0.788968
+ 1.189e+11Hz 0.592729 -0.789427
+ 1.19e+11Hz 0.592109 -0.789884
+ 1.191e+11Hz 0.591488 -0.790342
+ 1.192e+11Hz 0.590867 -0.790798
+ 1.193e+11Hz 0.590245 -0.791254
+ 1.194e+11Hz 0.589623 -0.79171
+ 1.195e+11Hz 0.589001 -0.792165
+ 1.196e+11Hz 0.588378 -0.79262
+ 1.197e+11Hz 0.587755 -0.793074
+ 1.198e+11Hz 0.587131 -0.793527
+ 1.199e+11Hz 0.586507 -0.79398
+ 1.2e+11Hz 0.585883 -0.794433
+ 1.201e+11Hz 0.585258 -0.794885
+ 1.202e+11Hz 0.584633 -0.795336
+ 1.203e+11Hz 0.584008 -0.795787
+ 1.204e+11Hz 0.583382 -0.796237
+ 1.205e+11Hz 0.582756 -0.796687
+ 1.206e+11Hz 0.58213 -0.797137
+ 1.207e+11Hz 0.581503 -0.797585
+ 1.208e+11Hz 0.580876 -0.798033
+ 1.209e+11Hz 0.580248 -0.798481
+ 1.21e+11Hz 0.579621 -0.798928
+ 1.211e+11Hz 0.578993 -0.799375
+ 1.212e+11Hz 0.578364 -0.799821
+ 1.213e+11Hz 0.577735 -0.800267
+ 1.214e+11Hz 0.577106 -0.800712
+ 1.215e+11Hz 0.576476 -0.801156
+ 1.216e+11Hz 0.575846 -0.8016
+ 1.217e+11Hz 0.575216 -0.802044
+ 1.218e+11Hz 0.574586 -0.802487
+ 1.219e+11Hz 0.573955 -0.802929
+ 1.22e+11Hz 0.573324 -0.803371
+ 1.221e+11Hz 0.572692 -0.803812
+ 1.222e+11Hz 0.57206 -0.804253
+ 1.223e+11Hz 0.571428 -0.804693
+ 1.224e+11Hz 0.570795 -0.805133
+ 1.225e+11Hz 0.570162 -0.805572
+ 1.226e+11Hz 0.569529 -0.806011
+ 1.227e+11Hz 0.568895 -0.806449
+ 1.228e+11Hz 0.568261 -0.806887
+ 1.229e+11Hz 0.567627 -0.807324
+ 1.23e+11Hz 0.566993 -0.807761
+ 1.231e+11Hz 0.566358 -0.808197
+ 1.232e+11Hz 0.565723 -0.808632
+ 1.233e+11Hz 0.565087 -0.809067
+ 1.234e+11Hz 0.564451 -0.809502
+ 1.235e+11Hz 0.563815 -0.809936
+ 1.236e+11Hz 0.563178 -0.810369
+ 1.237e+11Hz 0.562542 -0.810802
+ 1.238e+11Hz 0.561904 -0.811234
+ 1.239e+11Hz 0.561267 -0.811666
+ 1.24e+11Hz 0.560629 -0.812098
+ 1.241e+11Hz 0.559991 -0.812528
+ 1.242e+11Hz 0.559353 -0.812959
+ 1.243e+11Hz 0.558714 -0.813389
+ 1.244e+11Hz 0.558075 -0.813818
+ 1.245e+11Hz 0.557436 -0.814247
+ 1.246e+11Hz 0.556796 -0.814675
+ 1.247e+11Hz 0.556156 -0.815103
+ 1.248e+11Hz 0.555516 -0.81553
+ 1.249e+11Hz 0.554875 -0.815956
+ 1.25e+11Hz 0.554234 -0.816383
+ 1.251e+11Hz 0.553593 -0.816808
+ 1.252e+11Hz 0.552951 -0.817233
+ 1.253e+11Hz 0.552309 -0.817658
+ 1.254e+11Hz 0.551667 -0.818082
+ 1.255e+11Hz 0.551025 -0.818506
+ 1.256e+11Hz 0.550382 -0.818929
+ 1.257e+11Hz 0.549739 -0.819351
+ 1.258e+11Hz 0.549096 -0.819773
+ 1.259e+11Hz 0.548452 -0.820195
+ 1.26e+11Hz 0.547808 -0.820616
+ 1.261e+11Hz 0.547164 -0.821037
+ 1.262e+11Hz 0.546519 -0.821457
+ 1.263e+11Hz 0.545874 -0.821876
+ 1.264e+11Hz 0.545229 -0.822295
+ 1.265e+11Hz 0.544583 -0.822714
+ 1.266e+11Hz 0.543937 -0.823132
+ 1.267e+11Hz 0.543291 -0.823549
+ 1.268e+11Hz 0.542645 -0.823966
+ 1.269e+11Hz 0.541998 -0.824383
+ 1.27e+11Hz 0.541351 -0.824799
+ 1.271e+11Hz 0.540704 -0.825214
+ 1.272e+11Hz 0.540056 -0.825629
+ 1.273e+11Hz 0.539408 -0.826044
+ 1.274e+11Hz 0.53876 -0.826457
+ 1.275e+11Hz 0.538111 -0.826871
+ 1.276e+11Hz 0.537462 -0.827284
+ 1.277e+11Hz 0.536813 -0.827696
+ 1.278e+11Hz 0.536164 -0.828108
+ 1.279e+11Hz 0.535514 -0.82852
+ 1.28e+11Hz 0.534864 -0.828931
+ 1.281e+11Hz 0.534213 -0.829341
+ 1.282e+11Hz 0.533562 -0.829751
+ 1.283e+11Hz 0.532911 -0.830161
+ 1.284e+11Hz 0.53226 -0.83057
+ 1.285e+11Hz 0.531608 -0.830978
+ 1.286e+11Hz 0.530956 -0.831386
+ 1.287e+11Hz 0.530304 -0.831794
+ 1.288e+11Hz 0.529652 -0.832201
+ 1.289e+11Hz 0.528999 -0.832607
+ 1.29e+11Hz 0.528346 -0.833013
+ 1.291e+11Hz 0.527692 -0.833419
+ 1.292e+11Hz 0.527038 -0.833824
+ 1.293e+11Hz 0.526384 -0.834228
+ 1.294e+11Hz 0.52573 -0.834632
+ 1.295e+11Hz 0.525075 -0.835036
+ 1.296e+11Hz 0.52442 -0.835439
+ 1.297e+11Hz 0.523764 -0.835841
+ 1.298e+11Hz 0.523109 -0.836244
+ 1.299e+11Hz 0.522453 -0.836645
+ 1.3e+11Hz 0.521796 -0.837046
+ 1.301e+11Hz 0.52114 -0.837447
+ 1.302e+11Hz 0.520483 -0.837847
+ 1.303e+11Hz 0.519826 -0.838246
+ 1.304e+11Hz 0.519168 -0.838645
+ 1.305e+11Hz 0.51851 -0.839044
+ 1.306e+11Hz 0.517852 -0.839442
+ 1.307e+11Hz 0.517193 -0.83984
+ 1.308e+11Hz 0.516535 -0.840237
+ 1.309e+11Hz 0.515875 -0.840634
+ 1.31e+11Hz 0.515216 -0.84103
+ 1.311e+11Hz 0.514556 -0.841425
+ 1.312e+11Hz 0.513896 -0.84182
+ 1.313e+11Hz 0.513236 -0.842215
+ 1.314e+11Hz 0.512575 -0.842609
+ 1.315e+11Hz 0.511914 -0.843003
+ 1.316e+11Hz 0.511252 -0.843396
+ 1.317e+11Hz 0.510591 -0.843789
+ 1.318e+11Hz 0.509928 -0.844181
+ 1.319e+11Hz 0.509266 -0.844572
+ 1.32e+11Hz 0.508603 -0.844964
+ 1.321e+11Hz 0.50794 -0.845354
+ 1.322e+11Hz 0.507277 -0.845744
+ 1.323e+11Hz 0.506613 -0.846134
+ 1.324e+11Hz 0.505949 -0.846523
+ 1.325e+11Hz 0.505285 -0.846912
+ 1.326e+11Hz 0.50462 -0.8473
+ 1.327e+11Hz 0.503955 -0.847688
+ 1.328e+11Hz 0.50329 -0.848075
+ 1.329e+11Hz 0.502624 -0.848461
+ 1.33e+11Hz 0.501958 -0.848847
+ 1.331e+11Hz 0.501292 -0.849233
+ 1.332e+11Hz 0.500625 -0.849618
+ 1.333e+11Hz 0.499958 -0.850003
+ 1.334e+11Hz 0.499291 -0.850387
+ 1.335e+11Hz 0.498623 -0.85077
+ 1.336e+11Hz 0.497955 -0.851154
+ 1.337e+11Hz 0.497287 -0.851536
+ 1.338e+11Hz 0.496618 -0.851918
+ 1.339e+11Hz 0.495949 -0.8523
+ 1.34e+11Hz 0.49528 -0.852681
+ 1.341e+11Hz 0.49461 -0.853061
+ 1.342e+11Hz 0.49394 -0.853441
+ 1.343e+11Hz 0.49327 -0.853821
+ 1.344e+11Hz 0.492599 -0.8542
+ 1.345e+11Hz 0.491928 -0.854578
+ 1.346e+11Hz 0.491257 -0.854956
+ 1.347e+11Hz 0.490585 -0.855333
+ 1.348e+11Hz 0.489913 -0.85571
+ 1.349e+11Hz 0.489241 -0.856087
+ 1.35e+11Hz 0.488568 -0.856462
+ 1.351e+11Hz 0.487895 -0.856838
+ 1.352e+11Hz 0.487222 -0.857212
+ 1.353e+11Hz 0.486548 -0.857587
+ 1.354e+11Hz 0.485874 -0.85796
+ 1.355e+11Hz 0.4852 -0.858334
+ 1.356e+11Hz 0.484525 -0.858706
+ 1.357e+11Hz 0.48385 -0.859078
+ 1.358e+11Hz 0.483175 -0.85945
+ 1.359e+11Hz 0.482499 -0.859821
+ 1.36e+11Hz 0.481823 -0.860191
+ 1.361e+11Hz 0.481147 -0.860561
+ 1.362e+11Hz 0.48047 -0.860931
+ 1.363e+11Hz 0.479793 -0.8613
+ 1.364e+11Hz 0.479116 -0.861668
+ 1.365e+11Hz 0.478438 -0.862036
+ 1.366e+11Hz 0.47776 -0.862403
+ 1.367e+11Hz 0.477082 -0.86277
+ 1.368e+11Hz 0.476403 -0.863136
+ 1.369e+11Hz 0.475724 -0.863501
+ 1.37e+11Hz 0.475044 -0.863866
+ 1.371e+11Hz 0.474365 -0.864231
+ 1.372e+11Hz 0.473685 -0.864595
+ 1.373e+11Hz 0.473004 -0.864958
+ 1.374e+11Hz 0.472323 -0.865321
+ 1.375e+11Hz 0.471642 -0.865683
+ 1.376e+11Hz 0.470961 -0.866045
+ 1.377e+11Hz 0.470279 -0.866406
+ 1.378e+11Hz 0.469597 -0.866767
+ 1.379e+11Hz 0.468915 -0.867127
+ 1.38e+11Hz 0.468232 -0.867486
+ 1.381e+11Hz 0.467549 -0.867845
+ 1.382e+11Hz 0.466866 -0.868203
+ 1.383e+11Hz 0.466182 -0.868561
+ 1.384e+11Hz 0.465498 -0.868918
+ 1.385e+11Hz 0.464814 -0.869275
+ 1.386e+11Hz 0.464129 -0.869631
+ 1.387e+11Hz 0.463444 -0.869986
+ 1.388e+11Hz 0.462759 -0.870341
+ 1.389e+11Hz 0.462073 -0.870696
+ 1.39e+11Hz 0.461387 -0.871049
+ 1.391e+11Hz 0.460701 -0.871403
+ 1.392e+11Hz 0.460014 -0.871755
+ 1.393e+11Hz 0.459328 -0.872107
+ 1.394e+11Hz 0.45864 -0.872459
+ 1.395e+11Hz 0.457953 -0.872809
+ 1.396e+11Hz 0.457265 -0.87316
+ 1.397e+11Hz 0.456577 -0.873509
+ 1.398e+11Hz 0.455888 -0.873858
+ 1.399e+11Hz 0.4552 -0.874207
+ 1.4e+11Hz 0.45451 -0.874555
+ 1.401e+11Hz 0.453821 -0.874902
+ 1.402e+11Hz 0.453131 -0.875249
+ 1.403e+11Hz 0.452441 -0.875595
+ 1.404e+11Hz 0.451751 -0.87594
+ 1.405e+11Hz 0.45106 -0.876285
+ 1.406e+11Hz 0.450369 -0.87663
+ 1.407e+11Hz 0.449678 -0.876974
+ 1.408e+11Hz 0.448987 -0.877317
+ 1.409e+11Hz 0.448295 -0.877659
+ 1.41e+11Hz 0.447603 -0.878001
+ 1.411e+11Hz 0.44691 -0.878343
+ 1.412e+11Hz 0.446218 -0.878683
+ 1.413e+11Hz 0.445524 -0.879023
+ 1.414e+11Hz 0.444831 -0.879363
+ 1.415e+11Hz 0.444138 -0.879702
+ 1.416e+11Hz 0.443444 -0.88004
+ 1.417e+11Hz 0.44275 -0.880378
+ 1.418e+11Hz 0.442055 -0.880715
+ 1.419e+11Hz 0.44136 -0.881052
+ 1.42e+11Hz 0.440665 -0.881388
+ 1.421e+11Hz 0.43997 -0.881723
+ 1.422e+11Hz 0.439274 -0.882058
+ 1.423e+11Hz 0.438578 -0.882392
+ 1.424e+11Hz 0.437882 -0.882725
+ 1.425e+11Hz 0.437186 -0.883058
+ 1.426e+11Hz 0.436489 -0.883391
+ 1.427e+11Hz 0.435792 -0.883722
+ 1.428e+11Hz 0.435095 -0.884053
+ 1.429e+11Hz 0.434397 -0.884384
+ 1.43e+11Hz 0.433699 -0.884714
+ 1.431e+11Hz 0.433001 -0.885043
+ 1.432e+11Hz 0.432303 -0.885371
+ 1.433e+11Hz 0.431604 -0.885699
+ 1.434e+11Hz 0.430906 -0.886027
+ 1.435e+11Hz 0.430206 -0.886354
+ 1.436e+11Hz 0.429507 -0.88668
+ 1.437e+11Hz 0.428807 -0.887005
+ 1.438e+11Hz 0.428107 -0.88733
+ 1.439e+11Hz 0.427407 -0.887655
+ 1.44e+11Hz 0.426707 -0.887978
+ 1.441e+11Hz 0.426006 -0.888301
+ 1.442e+11Hz 0.425305 -0.888624
+ 1.443e+11Hz 0.424604 -0.888946
+ 1.444e+11Hz 0.423903 -0.889267
+ 1.445e+11Hz 0.423201 -0.889588
+ 1.446e+11Hz 0.422499 -0.889908
+ 1.447e+11Hz 0.421797 -0.890227
+ 1.448e+11Hz 0.421094 -0.890546
+ 1.449e+11Hz 0.420392 -0.890864
+ 1.45e+11Hz 0.419689 -0.891182
+ 1.451e+11Hz 0.418986 -0.891499
+ 1.452e+11Hz 0.418282 -0.891815
+ 1.453e+11Hz 0.417579 -0.892131
+ 1.454e+11Hz 0.416875 -0.892446
+ 1.455e+11Hz 0.416171 -0.89276
+ 1.456e+11Hz 0.415466 -0.893074
+ 1.457e+11Hz 0.414762 -0.893387
+ 1.458e+11Hz 0.414057 -0.8937
+ 1.459e+11Hz 0.413352 -0.894012
+ 1.46e+11Hz 0.412647 -0.894323
+ 1.461e+11Hz 0.411941 -0.894634
+ 1.462e+11Hz 0.411235 -0.894944
+ 1.463e+11Hz 0.410529 -0.895254
+ 1.464e+11Hz 0.409823 -0.895563
+ 1.465e+11Hz 0.409117 -0.895871
+ 1.466e+11Hz 0.40841 -0.896179
+ 1.467e+11Hz 0.407703 -0.896486
+ 1.468e+11Hz 0.406996 -0.896793
+ 1.469e+11Hz 0.406289 -0.897099
+ 1.47e+11Hz 0.405581 -0.897404
+ 1.471e+11Hz 0.404874 -0.897709
+ 1.472e+11Hz 0.404166 -0.898013
+ 1.473e+11Hz 0.403458 -0.898316
+ 1.474e+11Hz 0.402749 -0.898619
+ 1.475e+11Hz 0.402041 -0.898922
+ 1.476e+11Hz 0.401332 -0.899223
+ 1.477e+11Hz 0.400623 -0.899524
+ 1.478e+11Hz 0.399914 -0.899825
+ 1.479e+11Hz 0.399204 -0.900125
+ 1.48e+11Hz 0.398494 -0.900424
+ 1.481e+11Hz 0.397785 -0.900723
+ 1.482e+11Hz 0.397074 -0.901021
+ 1.483e+11Hz 0.396364 -0.901318
+ 1.484e+11Hz 0.395654 -0.901615
+ 1.485e+11Hz 0.394943 -0.901911
+ 1.486e+11Hz 0.394232 -0.902207
+ 1.487e+11Hz 0.393521 -0.902502
+ 1.488e+11Hz 0.39281 -0.902796
+ 1.489e+11Hz 0.392098 -0.90309
+ 1.49e+11Hz 0.391386 -0.903383
+ 1.491e+11Hz 0.390675 -0.903676
+ 1.492e+11Hz 0.389962 -0.903968
+ 1.493e+11Hz 0.38925 -0.904259
+ 1.494e+11Hz 0.388538 -0.90455
+ 1.495e+11Hz 0.387825 -0.90484
+ 1.496e+11Hz 0.387112 -0.90513
+ 1.497e+11Hz 0.386399 -0.905419
+ 1.498e+11Hz 0.385685 -0.905707
+ 1.499e+11Hz 0.384972 -0.905995
+ 1.5e+11Hz 0.384258 -0.906282
+ 1.501e+11Hz 0.383544 -0.906569
+ 1.502e+11Hz 0.38283 -0.906855
+ 1.503e+11Hz 0.382116 -0.907141
+ 1.504e+11Hz 0.381401 -0.907425
+ 1.505e+11Hz 0.380686 -0.90771
+ 1.506e+11Hz 0.379972 -0.907993
+ 1.507e+11Hz 0.379256 -0.908276
+ 1.508e+11Hz 0.378541 -0.908559
+ 1.509e+11Hz 0.377826 -0.908841
+ 1.51e+11Hz 0.37711 -0.909122
+ 1.511e+11Hz 0.376394 -0.909403
+ 1.512e+11Hz 0.375678 -0.909683
+ 1.513e+11Hz 0.374962 -0.909962
+ 1.514e+11Hz 0.374245 -0.910241
+ 1.515e+11Hz 0.373528 -0.91052
+ 1.516e+11Hz 0.372811 -0.910797
+ 1.517e+11Hz 0.372094 -0.911074
+ 1.518e+11Hz 0.371377 -0.911351
+ 1.519e+11Hz 0.37066 -0.911627
+ 1.52e+11Hz 0.369942 -0.911902
+ 1.521e+11Hz 0.369224 -0.912177
+ 1.522e+11Hz 0.368506 -0.912451
+ 1.523e+11Hz 0.367788 -0.912725
+ 1.524e+11Hz 0.367069 -0.912998
+ 1.525e+11Hz 0.366351 -0.91327
+ 1.526e+11Hz 0.365632 -0.913542
+ 1.527e+11Hz 0.364913 -0.913813
+ 1.528e+11Hz 0.364193 -0.914084
+ 1.529e+11Hz 0.363474 -0.914354
+ 1.53e+11Hz 0.362754 -0.914623
+ 1.531e+11Hz 0.362034 -0.914892
+ 1.532e+11Hz 0.361314 -0.915161
+ 1.533e+11Hz 0.360594 -0.915428
+ 1.534e+11Hz 0.359874 -0.915695
+ 1.535e+11Hz 0.359153 -0.915962
+ 1.536e+11Hz 0.358432 -0.916228
+ 1.537e+11Hz 0.357711 -0.916493
+ 1.538e+11Hz 0.35699 -0.916758
+ 1.539e+11Hz 0.356269 -0.917022
+ 1.54e+11Hz 0.355547 -0.917285
+ 1.541e+11Hz 0.354825 -0.917548
+ 1.542e+11Hz 0.354103 -0.91781
+ 1.543e+11Hz 0.353381 -0.918072
+ 1.544e+11Hz 0.352659 -0.918333
+ 1.545e+11Hz 0.351936 -0.918594
+ 1.546e+11Hz 0.351213 -0.918854
+ 1.547e+11Hz 0.35049 -0.919113
+ 1.548e+11Hz 0.349767 -0.919372
+ 1.549e+11Hz 0.349044 -0.91963
+ 1.55e+11Hz 0.34832 -0.919888
+ 1.551e+11Hz 0.347596 -0.920144
+ 1.552e+11Hz 0.346872 -0.920401
+ 1.553e+11Hz 0.346148 -0.920657
+ 1.554e+11Hz 0.345424 -0.920912
+ 1.555e+11Hz 0.344699 -0.921166
+ 1.556e+11Hz 0.343974 -0.92142
+ 1.557e+11Hz 0.343249 -0.921673
+ 1.558e+11Hz 0.342524 -0.921926
+ 1.559e+11Hz 0.341799 -0.922178
+ 1.56e+11Hz 0.341073 -0.92243
+ 1.561e+11Hz 0.340348 -0.922681
+ 1.562e+11Hz 0.339622 -0.922931
+ 1.563e+11Hz 0.338895 -0.923181
+ 1.564e+11Hz 0.338169 -0.92343
+ 1.565e+11Hz 0.337443 -0.923678
+ 1.566e+11Hz 0.336716 -0.923926
+ 1.567e+11Hz 0.335989 -0.924173
+ 1.568e+11Hz 0.335262 -0.92442
+ 1.569e+11Hz 0.334535 -0.924666
+ 1.57e+11Hz 0.333807 -0.924911
+ 1.571e+11Hz 0.333079 -0.925156
+ 1.572e+11Hz 0.332351 -0.9254
+ 1.573e+11Hz 0.331623 -0.925643
+ 1.574e+11Hz 0.330895 -0.925886
+ 1.575e+11Hz 0.330167 -0.926129
+ 1.576e+11Hz 0.329438 -0.92637
+ 1.577e+11Hz 0.328709 -0.926611
+ 1.578e+11Hz 0.32798 -0.926852
+ 1.579e+11Hz 0.327251 -0.927091
+ 1.58e+11Hz 0.326521 -0.927331
+ 1.581e+11Hz 0.325792 -0.927569
+ 1.582e+11Hz 0.325062 -0.927807
+ 1.583e+11Hz 0.324332 -0.928044
+ 1.584e+11Hz 0.323602 -0.928281
+ 1.585e+11Hz 0.322872 -0.928517
+ 1.586e+11Hz 0.322141 -0.928752
+ 1.587e+11Hz 0.32141 -0.928987
+ 1.588e+11Hz 0.320679 -0.929221
+ 1.589e+11Hz 0.319948 -0.929454
+ 1.59e+11Hz 0.319217 -0.929687
+ 1.591e+11Hz 0.318486 -0.929919
+ 1.592e+11Hz 0.317754 -0.930151
+ 1.593e+11Hz 0.317022 -0.930382
+ 1.594e+11Hz 0.31629 -0.930612
+ 1.595e+11Hz 0.315558 -0.930842
+ 1.596e+11Hz 0.314826 -0.931071
+ 1.597e+11Hz 0.314093 -0.931299
+ 1.598e+11Hz 0.313361 -0.931526
+ 1.599e+11Hz 0.312628 -0.931753
+ 1.6e+11Hz 0.311895 -0.93198
+ 1.601e+11Hz 0.311162 -0.932206
+ 1.602e+11Hz 0.310428 -0.932431
+ 1.603e+11Hz 0.309695 -0.932655
+ 1.604e+11Hz 0.308961 -0.932879
+ 1.605e+11Hz 0.308227 -0.933102
+ 1.606e+11Hz 0.307493 -0.933324
+ 1.607e+11Hz 0.306759 -0.933546
+ 1.608e+11Hz 0.306025 -0.933767
+ 1.609e+11Hz 0.305291 -0.933988
+ 1.61e+11Hz 0.304556 -0.934207
+ 1.611e+11Hz 0.303821 -0.934426
+ 1.612e+11Hz 0.303086 -0.934645
+ 1.613e+11Hz 0.302351 -0.934863
+ 1.614e+11Hz 0.301616 -0.93508
+ 1.615e+11Hz 0.300881 -0.935296
+ 1.616e+11Hz 0.300145 -0.935512
+ 1.617e+11Hz 0.299409 -0.935727
+ 1.618e+11Hz 0.298674 -0.935942
+ 1.619e+11Hz 0.297938 -0.936155
+ 1.62e+11Hz 0.297202 -0.936369
+ 1.621e+11Hz 0.296465 -0.936581
+ 1.622e+11Hz 0.295729 -0.936793
+ 1.623e+11Hz 0.294993 -0.937004
+ 1.624e+11Hz 0.294256 -0.937214
+ 1.625e+11Hz 0.293519 -0.937424
+ 1.626e+11Hz 0.292782 -0.937633
+ 1.627e+11Hz 0.292046 -0.937842
+ 1.628e+11Hz 0.291308 -0.938049
+ 1.629e+11Hz 0.290571 -0.938256
+ 1.63e+11Hz 0.289834 -0.938463
+ 1.631e+11Hz 0.289096 -0.938668
+ 1.632e+11Hz 0.288359 -0.938873
+ 1.633e+11Hz 0.287621 -0.939078
+ 1.634e+11Hz 0.286883 -0.939281
+ 1.635e+11Hz 0.286145 -0.939484
+ 1.636e+11Hz 0.285407 -0.939687
+ 1.637e+11Hz 0.284669 -0.939888
+ 1.638e+11Hz 0.283931 -0.940089
+ 1.639e+11Hz 0.283193 -0.940289
+ 1.64e+11Hz 0.282455 -0.940489
+ 1.641e+11Hz 0.281716 -0.940688
+ 1.642e+11Hz 0.280977 -0.940886
+ 1.643e+11Hz 0.280239 -0.941084
+ 1.644e+11Hz 0.2795 -0.941281
+ 1.645e+11Hz 0.278761 -0.941477
+ 1.646e+11Hz 0.278022 -0.941672
+ 1.647e+11Hz 0.277283 -0.941867
+ 1.648e+11Hz 0.276544 -0.942061
+ 1.649e+11Hz 0.275805 -0.942255
+ 1.65e+11Hz 0.275066 -0.942447
+ 1.651e+11Hz 0.274327 -0.94264
+ 1.652e+11Hz 0.273587 -0.942831
+ 1.653e+11Hz 0.272848 -0.943022
+ 1.654e+11Hz 0.272108 -0.943212
+ 1.655e+11Hz 0.271369 -0.943401
+ 1.656e+11Hz 0.270629 -0.94359
+ 1.657e+11Hz 0.269889 -0.943778
+ 1.658e+11Hz 0.26915 -0.943965
+ 1.659e+11Hz 0.26841 -0.944152
+ 1.66e+11Hz 0.26767 -0.944338
+ 1.661e+11Hz 0.26693 -0.944523
+ 1.662e+11Hz 0.26619 -0.944708
+ 1.663e+11Hz 0.26545 -0.944892
+ 1.664e+11Hz 0.26471 -0.945075
+ 1.665e+11Hz 0.26397 -0.945258
+ 1.666e+11Hz 0.26323 -0.94544
+ 1.667e+11Hz 0.26249 -0.945621
+ 1.668e+11Hz 0.26175 -0.945802
+ 1.669e+11Hz 0.26101 -0.945982
+ 1.67e+11Hz 0.26027 -0.946161
+ 1.671e+11Hz 0.259529 -0.946339
+ 1.672e+11Hz 0.258789 -0.946517
+ 1.673e+11Hz 0.258049 -0.946695
+ 1.674e+11Hz 0.257309 -0.946871
+ 1.675e+11Hz 0.256568 -0.947047
+ 1.676e+11Hz 0.255828 -0.947223
+ 1.677e+11Hz 0.255088 -0.947397
+ 1.678e+11Hz 0.254348 -0.947571
+ 1.679e+11Hz 0.253607 -0.947744
+ 1.68e+11Hz 0.252867 -0.947917
+ 1.681e+11Hz 0.252127 -0.948089
+ 1.682e+11Hz 0.251386 -0.94826
+ 1.683e+11Hz 0.250646 -0.948431
+ 1.684e+11Hz 0.249906 -0.948601
+ 1.685e+11Hz 0.249165 -0.948771
+ 1.686e+11Hz 0.248425 -0.948939
+ 1.687e+11Hz 0.247685 -0.949108
+ 1.688e+11Hz 0.246944 -0.949275
+ 1.689e+11Hz 0.246204 -0.949442
+ 1.69e+11Hz 0.245464 -0.949608
+ 1.691e+11Hz 0.244724 -0.949774
+ 1.692e+11Hz 0.243983 -0.949939
+ 1.693e+11Hz 0.243243 -0.950103
+ 1.694e+11Hz 0.242503 -0.950266
+ 1.695e+11Hz 0.241763 -0.950429
+ 1.696e+11Hz 0.241023 -0.950592
+ 1.697e+11Hz 0.240283 -0.950754
+ 1.698e+11Hz 0.239543 -0.950915
+ 1.699e+11Hz 0.238803 -0.951075
+ 1.7e+11Hz 0.238063 -0.951235
+ 1.701e+11Hz 0.237323 -0.951394
+ 1.702e+11Hz 0.236583 -0.951553
+ 1.703e+11Hz 0.235843 -0.951711
+ 1.704e+11Hz 0.235103 -0.951869
+ 1.705e+11Hz 0.234363 -0.952025
+ 1.706e+11Hz 0.233623 -0.952182
+ 1.707e+11Hz 0.232884 -0.952337
+ 1.708e+11Hz 0.232144 -0.952492
+ 1.709e+11Hz 0.231404 -0.952647
+ 1.71e+11Hz 0.230665 -0.952801
+ 1.711e+11Hz 0.229925 -0.952954
+ 1.712e+11Hz 0.229185 -0.953106
+ 1.713e+11Hz 0.228446 -0.953258
+ 1.714e+11Hz 0.227706 -0.95341
+ 1.715e+11Hz 0.226967 -0.953561
+ 1.716e+11Hz 0.226228 -0.953711
+ 1.717e+11Hz 0.225488 -0.953861
+ 1.718e+11Hz 0.224749 -0.95401
+ 1.719e+11Hz 0.22401 -0.954158
+ 1.72e+11Hz 0.223271 -0.954306
+ 1.721e+11Hz 0.222532 -0.954453
+ 1.722e+11Hz 0.221793 -0.9546
+ 1.723e+11Hz 0.221054 -0.954747
+ 1.724e+11Hz 0.220315 -0.954892
+ 1.725e+11Hz 0.219576 -0.955037
+ 1.726e+11Hz 0.218837 -0.955182
+ 1.727e+11Hz 0.218098 -0.955326
+ 1.728e+11Hz 0.21736 -0.955469
+ 1.729e+11Hz 0.216621 -0.955612
+ 1.73e+11Hz 0.215882 -0.955754
+ 1.731e+11Hz 0.215144 -0.955896
+ 1.732e+11Hz 0.214405 -0.956037
+ 1.733e+11Hz 0.213667 -0.956178
+ 1.734e+11Hz 0.212929 -0.956318
+ 1.735e+11Hz 0.21219 -0.956458
+ 1.736e+11Hz 0.211452 -0.956597
+ 1.737e+11Hz 0.210714 -0.956735
+ 1.738e+11Hz 0.209976 -0.956873
+ 1.739e+11Hz 0.209237 -0.95701
+ 1.74e+11Hz 0.208499 -0.957147
+ 1.741e+11Hz 0.207761 -0.957284
+ 1.742e+11Hz 0.207023 -0.957419
+ 1.743e+11Hz 0.206286 -0.957555
+ 1.744e+11Hz 0.205548 -0.957689
+ 1.745e+11Hz 0.20481 -0.957824
+ 1.746e+11Hz 0.204072 -0.957957
+ 1.747e+11Hz 0.203335 -0.958091
+ 1.748e+11Hz 0.202597 -0.958223
+ 1.749e+11Hz 0.201859 -0.958356
+ 1.75e+11Hz 0.201122 -0.958487
+ 1.751e+11Hz 0.200384 -0.958618
+ 1.752e+11Hz 0.199647 -0.958749
+ 1.753e+11Hz 0.19891 -0.958879
+ 1.754e+11Hz 0.198172 -0.959009
+ 1.755e+11Hz 0.197435 -0.959138
+ 1.756e+11Hz 0.196698 -0.959267
+ 1.757e+11Hz 0.195961 -0.959395
+ 1.758e+11Hz 0.195223 -0.959523
+ 1.759e+11Hz 0.194486 -0.95965
+ 1.76e+11Hz 0.193749 -0.959776
+ 1.761e+11Hz 0.193012 -0.959903
+ 1.762e+11Hz 0.192275 -0.960028
+ 1.763e+11Hz 0.191538 -0.960154
+ 1.764e+11Hz 0.190801 -0.960278
+ 1.765e+11Hz 0.190064 -0.960402
+ 1.766e+11Hz 0.189328 -0.960526
+ 1.767e+11Hz 0.188591 -0.96065
+ 1.768e+11Hz 0.187854 -0.960772
+ 1.769e+11Hz 0.187117 -0.960895
+ 1.77e+11Hz 0.186381 -0.961017
+ 1.771e+11Hz 0.185644 -0.961138
+ 1.772e+11Hz 0.184907 -0.961259
+ 1.773e+11Hz 0.184171 -0.961379
+ 1.774e+11Hz 0.183434 -0.961499
+ 1.775e+11Hz 0.182697 -0.961619
+ 1.776e+11Hz 0.181961 -0.961738
+ 1.777e+11Hz 0.181224 -0.961856
+ 1.778e+11Hz 0.180488 -0.961974
+ 1.779e+11Hz 0.179751 -0.962092
+ 1.78e+11Hz 0.179015 -0.962209
+ 1.781e+11Hz 0.178278 -0.962326
+ 1.782e+11Hz 0.177542 -0.962442
+ 1.783e+11Hz 0.176805 -0.962558
+ 1.784e+11Hz 0.176069 -0.962673
+ 1.785e+11Hz 0.175333 -0.962788
+ 1.786e+11Hz 0.174596 -0.962902
+ 1.787e+11Hz 0.17386 -0.963016
+ 1.788e+11Hz 0.173123 -0.96313
+ 1.789e+11Hz 0.172387 -0.963243
+ 1.79e+11Hz 0.171651 -0.963355
+ 1.791e+11Hz 0.170914 -0.963468
+ 1.792e+11Hz 0.170178 -0.963579
+ 1.793e+11Hz 0.169441 -0.96369
+ 1.794e+11Hz 0.168705 -0.963801
+ 1.795e+11Hz 0.167968 -0.963911
+ 1.796e+11Hz 0.167232 -0.964021
+ 1.797e+11Hz 0.166496 -0.964131
+ 1.798e+11Hz 0.165759 -0.96424
+ 1.799e+11Hz 0.165023 -0.964348
+ 1.8e+11Hz 0.164286 -0.964456
+ 1.801e+11Hz 0.16355 -0.964564
+ 1.802e+11Hz 0.162813 -0.964671
+ 1.803e+11Hz 0.162077 -0.964778
+ 1.804e+11Hz 0.16134 -0.964884
+ 1.805e+11Hz 0.160604 -0.96499
+ 1.806e+11Hz 0.159867 -0.965095
+ 1.807e+11Hz 0.15913 -0.9652
+ 1.808e+11Hz 0.158394 -0.965304
+ 1.809e+11Hz 0.157657 -0.965408
+ 1.81e+11Hz 0.15692 -0.965512
+ 1.811e+11Hz 0.156184 -0.965615
+ 1.812e+11Hz 0.155447 -0.965718
+ 1.813e+11Hz 0.15471 -0.96582
+ 1.814e+11Hz 0.153973 -0.965921
+ 1.815e+11Hz 0.153236 -0.966023
+ 1.816e+11Hz 0.152499 -0.966124
+ 1.817e+11Hz 0.151762 -0.966224
+ 1.818e+11Hz 0.151025 -0.966324
+ 1.819e+11Hz 0.150288 -0.966423
+ 1.82e+11Hz 0.149551 -0.966522
+ 1.821e+11Hz 0.148814 -0.966621
+ 1.822e+11Hz 0.148077 -0.966719
+ 1.823e+11Hz 0.14734 -0.966817
+ 1.824e+11Hz 0.146602 -0.966914
+ 1.825e+11Hz 0.145865 -0.967011
+ 1.826e+11Hz 0.145128 -0.967107
+ 1.827e+11Hz 0.14439 -0.967203
+ 1.828e+11Hz 0.143653 -0.967298
+ 1.829e+11Hz 0.142915 -0.967393
+ 1.83e+11Hz 0.142178 -0.967488
+ 1.831e+11Hz 0.14144 -0.967582
+ 1.832e+11Hz 0.140702 -0.967675
+ 1.833e+11Hz 0.139965 -0.967768
+ 1.834e+11Hz 0.139227 -0.967861
+ 1.835e+11Hz 0.138489 -0.967953
+ 1.836e+11Hz 0.137751 -0.968045
+ 1.837e+11Hz 0.137013 -0.968136
+ 1.838e+11Hz 0.136275 -0.968227
+ 1.839e+11Hz 0.135537 -0.968317
+ 1.84e+11Hz 0.134799 -0.968407
+ 1.841e+11Hz 0.13406 -0.968496
+ 1.842e+11Hz 0.133322 -0.968585
+ 1.843e+11Hz 0.132584 -0.968673
+ 1.844e+11Hz 0.131845 -0.968761
+ 1.845e+11Hz 0.131107 -0.968849
+ 1.846e+11Hz 0.130368 -0.968936
+ 1.847e+11Hz 0.129629 -0.969022
+ 1.848e+11Hz 0.128891 -0.969109
+ 1.849e+11Hz 0.128152 -0.969194
+ 1.85e+11Hz 0.127413 -0.969279
+ 1.851e+11Hz 0.126674 -0.969364
+ 1.852e+11Hz 0.125935 -0.969448
+ 1.853e+11Hz 0.125196 -0.969532
+ 1.854e+11Hz 0.124457 -0.969615
+ 1.855e+11Hz 0.123717 -0.969698
+ 1.856e+11Hz 0.122978 -0.96978
+ 1.857e+11Hz 0.122239 -0.969862
+ 1.858e+11Hz 0.121499 -0.969943
+ 1.859e+11Hz 0.120759 -0.970024
+ 1.86e+11Hz 0.12002 -0.970104
+ 1.861e+11Hz 0.11928 -0.970184
+ 1.862e+11Hz 0.11854 -0.970263
+ 1.863e+11Hz 0.1178 -0.970342
+ 1.864e+11Hz 0.11706 -0.97042
+ 1.865e+11Hz 0.11632 -0.970498
+ 1.866e+11Hz 0.11558 -0.970576
+ 1.867e+11Hz 0.11484 -0.970652
+ 1.868e+11Hz 0.1141 -0.970729
+ 1.869e+11Hz 0.113359 -0.970805
+ 1.87e+11Hz 0.112619 -0.97088
+ 1.871e+11Hz 0.111878 -0.970955
+ 1.872e+11Hz 0.111138 -0.971029
+ 1.873e+11Hz 0.110397 -0.971103
+ 1.874e+11Hz 0.109656 -0.971177
+ 1.875e+11Hz 0.108915 -0.971249
+ 1.876e+11Hz 0.108175 -0.971322
+ 1.877e+11Hz 0.107434 -0.971394
+ 1.878e+11Hz 0.106692 -0.971465
+ 1.879e+11Hz 0.105951 -0.971536
+ 1.88e+11Hz 0.10521 -0.971606
+ 1.881e+11Hz 0.104469 -0.971676
+ 1.882e+11Hz 0.103727 -0.971745
+ 1.883e+11Hz 0.102986 -0.971814
+ 1.884e+11Hz 0.102244 -0.971883
+ 1.885e+11Hz 0.101503 -0.97195
+ 1.886e+11Hz 0.100761 -0.972018
+ 1.887e+11Hz 0.100019 -0.972084
+ 1.888e+11Hz 0.0992772 -0.972151
+ 1.889e+11Hz 0.0985352 -0.972216
+ 1.89e+11Hz 0.0977932 -0.972282
+ 1.891e+11Hz 0.0970511 -0.972346
+ 1.892e+11Hz 0.0963089 -0.972411
+ 1.893e+11Hz 0.0955666 -0.972474
+ 1.894e+11Hz 0.0948242 -0.972537
+ 1.895e+11Hz 0.0940818 -0.9726
+ 1.896e+11Hz 0.0933393 -0.972662
+ 1.897e+11Hz 0.0925967 -0.972724
+ 1.898e+11Hz 0.0918541 -0.972785
+ 1.899e+11Hz 0.0911114 -0.972845
+ 1.9e+11Hz 0.0903686 -0.972905
+ 1.901e+11Hz 0.0896257 -0.972965
+ 1.902e+11Hz 0.0888827 -0.973024
+ 1.903e+11Hz 0.0881397 -0.973082
+ 1.904e+11Hz 0.0873966 -0.97314
+ 1.905e+11Hz 0.0866534 -0.973198
+ 1.906e+11Hz 0.0859102 -0.973254
+ 1.907e+11Hz 0.0851669 -0.973311
+ 1.908e+11Hz 0.0844235 -0.973367
+ 1.909e+11Hz 0.08368 -0.973422
+ 1.91e+11Hz 0.0829365 -0.973477
+ 1.911e+11Hz 0.0821929 -0.973531
+ 1.912e+11Hz 0.0814492 -0.973584
+ 1.913e+11Hz 0.0807055 -0.973638
+ 1.914e+11Hz 0.0799617 -0.97369
+ 1.915e+11Hz 0.0792178 -0.973742
+ 1.916e+11Hz 0.0784739 -0.973794
+ 1.917e+11Hz 0.0777299 -0.973845
+ 1.918e+11Hz 0.0769858 -0.973895
+ 1.919e+11Hz 0.0762416 -0.973945
+ 1.92e+11Hz 0.0754974 -0.973995
+ 1.921e+11Hz 0.0747532 -0.974043
+ 1.922e+11Hz 0.0740088 -0.974092
+ 1.923e+11Hz 0.0732644 -0.97414
+ 1.924e+11Hz 0.0725199 -0.974187
+ 1.925e+11Hz 0.0717754 -0.974233
+ 1.926e+11Hz 0.0710308 -0.97428
+ 1.927e+11Hz 0.0702861 -0.974325
+ 1.928e+11Hz 0.0695414 -0.97437
+ 1.929e+11Hz 0.0687966 -0.974415
+ 1.93e+11Hz 0.0680518 -0.974459
+ 1.931e+11Hz 0.0673068 -0.974502
+ 1.932e+11Hz 0.0665619 -0.974545
+ 1.933e+11Hz 0.0658168 -0.974588
+ 1.934e+11Hz 0.0650717 -0.974629
+ 1.935e+11Hz 0.0643266 -0.974671
+ 1.936e+11Hz 0.0635814 -0.974711
+ 1.937e+11Hz 0.0628361 -0.974752
+ 1.938e+11Hz 0.0620907 -0.974791
+ 1.939e+11Hz 0.0613453 -0.97483
+ 1.94e+11Hz 0.0605999 -0.974869
+ 1.941e+11Hz 0.0598544 -0.974907
+ 1.942e+11Hz 0.0591088 -0.974944
+ 1.943e+11Hz 0.0583632 -0.974981
+ 1.944e+11Hz 0.0576175 -0.975018
+ 1.945e+11Hz 0.0568717 -0.975054
+ 1.946e+11Hz 0.0561259 -0.975089
+ 1.947e+11Hz 0.0553801 -0.975123
+ 1.948e+11Hz 0.0546342 -0.975158
+ 1.949e+11Hz 0.0538882 -0.975191
+ 1.95e+11Hz 0.0531422 -0.975224
+ 1.951e+11Hz 0.0523961 -0.975257
+ 1.952e+11Hz 0.05165 -0.975289
+ 1.953e+11Hz 0.0509038 -0.97532
+ 1.954e+11Hz 0.0501575 -0.975351
+ 1.955e+11Hz 0.0494112 -0.975381
+ 1.956e+11Hz 0.0486649 -0.975411
+ 1.957e+11Hz 0.0479185 -0.97544
+ 1.958e+11Hz 0.047172 -0.975469
+ 1.959e+11Hz 0.0464255 -0.975497
+ 1.96e+11Hz 0.045679 -0.975525
+ 1.961e+11Hz 0.0449323 -0.975552
+ 1.962e+11Hz 0.0441857 -0.975578
+ 1.963e+11Hz 0.043439 -0.975604
+ 1.964e+11Hz 0.0426922 -0.975629
+ 1.965e+11Hz 0.0419454 -0.975654
+ 1.966e+11Hz 0.0411985 -0.975678
+ 1.967e+11Hz 0.0404515 -0.975702
+ 1.968e+11Hz 0.0397046 -0.975725
+ 1.969e+11Hz 0.0389575 -0.975748
+ 1.97e+11Hz 0.0382104 -0.97577
+ 1.971e+11Hz 0.0374633 -0.975791
+ 1.972e+11Hz 0.0367161 -0.975812
+ 1.973e+11Hz 0.0359689 -0.975832
+ 1.974e+11Hz 0.0352216 -0.975852
+ 1.975e+11Hz 0.0344743 -0.975871
+ 1.976e+11Hz 0.0337269 -0.97589
+ 1.977e+11Hz 0.0329794 -0.975908
+ 1.978e+11Hz 0.032232 -0.975925
+ 1.979e+11Hz 0.0314844 -0.975942
+ 1.98e+11Hz 0.0307368 -0.975958
+ 1.981e+11Hz 0.0299892 -0.975974
+ 1.982e+11Hz 0.0292415 -0.975989
+ 1.983e+11Hz 0.0284938 -0.976004
+ 1.984e+11Hz 0.027746 -0.976018
+ 1.985e+11Hz 0.0269982 -0.976031
+ 1.986e+11Hz 0.0262503 -0.976044
+ 1.987e+11Hz 0.0255024 -0.976057
+ 1.988e+11Hz 0.0247544 -0.976068
+ 1.989e+11Hz 0.0240064 -0.97608
+ 1.99e+11Hz 0.0232584 -0.97609
+ 1.991e+11Hz 0.0225103 -0.9761
+ 1.992e+11Hz 0.0217621 -0.97611
+ 1.993e+11Hz 0.0210139 -0.976119
+ 1.994e+11Hz 0.0202657 -0.976127
+ 1.995e+11Hz 0.0195174 -0.976135
+ 1.996e+11Hz 0.018769 -0.976142
+ 1.997e+11Hz 0.0180206 -0.976148
+ 1.998e+11Hz 0.0172722 -0.976154
+ 1.999e+11Hz 0.0165238 -0.97616
+ 2e+11Hz 0.0157752 -0.976165
+ 2.001e+11Hz 0.0150267 -0.976169
+ 2.002e+11Hz 0.0142781 -0.976173
+ 2.003e+11Hz 0.0135295 -0.976176
+ 2.004e+11Hz 0.0127808 -0.976178
+ 2.005e+11Hz 0.0120321 -0.97618
+ 2.006e+11Hz 0.0112833 -0.976181
+ 2.007e+11Hz 0.0105345 -0.976182
+ 2.008e+11Hz 0.00978566 -0.976182
+ 2.009e+11Hz 0.00903679 -0.976182
+ 2.01e+11Hz 0.00828787 -0.976181
+ 2.011e+11Hz 0.00753892 -0.976179
+ 2.012e+11Hz 0.00678993 -0.976177
+ 2.013e+11Hz 0.00604091 -0.976174
+ 2.014e+11Hz 0.00529185 -0.97617
+ 2.015e+11Hz 0.00454275 -0.976166
+ 2.016e+11Hz 0.00379363 -0.976162
+ 2.017e+11Hz 0.00304447 -0.976156
+ 2.018e+11Hz 0.00229528 -0.97615
+ 2.019e+11Hz 0.00154605 -0.976144
+ 2.02e+11Hz 0.000796802 -0.976137
+ 2.021e+11Hz 4.7521e-05 -0.976129
+ 2.022e+11Hz -0.000701788 -0.976121
+ 2.023e+11Hz -0.00145112 -0.976112
+ 2.024e+11Hz -0.00220049 -0.976102
+ 2.025e+11Hz -0.00294987 -0.976092
+ 2.026e+11Hz -0.00369929 -0.976081
+ 2.027e+11Hz -0.00444872 -0.97607
+ 2.028e+11Hz -0.00519818 -0.976058
+ 2.029e+11Hz -0.00594765 -0.976045
+ 2.03e+11Hz -0.00669715 -0.976032
+ 2.031e+11Hz -0.00744666 -0.976018
+ 2.032e+11Hz -0.00819619 -0.976004
+ 2.033e+11Hz -0.00894573 -0.975988
+ 2.034e+11Hz -0.00969529 -0.975973
+ 2.035e+11Hz -0.0104449 -0.975956
+ 2.036e+11Hz -0.0111944 -0.975939
+ 2.037e+11Hz -0.011944 -0.975922
+ 2.038e+11Hz -0.0126936 -0.975903
+ 2.039e+11Hz -0.0134432 -0.975884
+ 2.04e+11Hz -0.0141928 -0.975865
+ 2.041e+11Hz -0.0149425 -0.975845
+ 2.042e+11Hz -0.0156921 -0.975824
+ 2.043e+11Hz -0.0164417 -0.975802
+ 2.044e+11Hz -0.0171913 -0.97578
+ 2.045e+11Hz -0.0179409 -0.975758
+ 2.046e+11Hz -0.0186905 -0.975734
+ 2.047e+11Hz -0.0194401 -0.97571
+ 2.048e+11Hz -0.0201897 -0.975686
+ 2.049e+11Hz -0.0209393 -0.97566
+ 2.05e+11Hz -0.0216888 -0.975634
+ 2.051e+11Hz -0.0224384 -0.975608
+ 2.052e+11Hz -0.0231879 -0.975581
+ 2.053e+11Hz -0.0239374 -0.975553
+ 2.054e+11Hz -0.0246869 -0.975524
+ 2.055e+11Hz -0.0254363 -0.975495
+ 2.056e+11Hz -0.0261858 -0.975465
+ 2.057e+11Hz -0.0269352 -0.975435
+ 2.058e+11Hz -0.0276845 -0.975403
+ 2.059e+11Hz -0.0284339 -0.975372
+ 2.06e+11Hz -0.0291832 -0.975339
+ 2.061e+11Hz -0.0299325 -0.975306
+ 2.062e+11Hz -0.0306817 -0.975272
+ 2.063e+11Hz -0.0314309 -0.975238
+ 2.064e+11Hz -0.03218 -0.975203
+ 2.065e+11Hz -0.0329291 -0.975167
+ 2.066e+11Hz -0.0336781 -0.975131
+ 2.067e+11Hz -0.0344271 -0.975094
+ 2.068e+11Hz -0.035176 -0.975056
+ 2.069e+11Hz -0.0359249 -0.975017
+ 2.07e+11Hz -0.0366737 -0.974978
+ 2.071e+11Hz -0.0374225 -0.974939
+ 2.072e+11Hz -0.0381711 -0.974898
+ 2.073e+11Hz -0.0389197 -0.974857
+ 2.074e+11Hz -0.0396683 -0.974816
+ 2.075e+11Hz -0.0404167 -0.974773
+ 2.076e+11Hz -0.0411651 -0.97473
+ 2.077e+11Hz -0.0419134 -0.974686
+ 2.078e+11Hz -0.0426616 -0.974642
+ 2.079e+11Hz -0.0434098 -0.974597
+ 2.08e+11Hz -0.0441578 -0.974551
+ 2.081e+11Hz -0.0449058 -0.974505
+ 2.082e+11Hz -0.0456536 -0.974458
+ 2.083e+11Hz -0.0464014 -0.97441
+ 2.084e+11Hz -0.047149 -0.974362
+ 2.085e+11Hz -0.0478966 -0.974313
+ 2.086e+11Hz -0.048644 -0.974263
+ 2.087e+11Hz -0.0493913 -0.974213
+ 2.088e+11Hz -0.0501385 -0.974162
+ 2.089e+11Hz -0.0508856 -0.974111
+ 2.09e+11Hz -0.0516326 -0.974058
+ 2.091e+11Hz -0.0523794 -0.974005
+ 2.092e+11Hz -0.0531262 -0.973952
+ 2.093e+11Hz -0.0538728 -0.973897
+ 2.094e+11Hz -0.0546192 -0.973843
+ 2.095e+11Hz -0.0553656 -0.973787
+ 2.096e+11Hz -0.0561117 -0.973731
+ 2.097e+11Hz -0.0568578 -0.973674
+ 2.098e+11Hz -0.0576037 -0.973616
+ 2.099e+11Hz -0.0583494 -0.973558
+ 2.1e+11Hz -0.059095 -0.973499
+ 2.101e+11Hz -0.0598405 -0.97344
+ 2.102e+11Hz -0.0605858 -0.97338
+ 2.103e+11Hz -0.0613309 -0.973319
+ 2.104e+11Hz -0.0620758 -0.973257
+ 2.105e+11Hz -0.0628206 -0.973195
+ 2.106e+11Hz -0.0635652 -0.973133
+ 2.107e+11Hz -0.0643097 -0.973069
+ 2.108e+11Hz -0.065054 -0.973005
+ 2.109e+11Hz -0.0657981 -0.972941
+ 2.11e+11Hz -0.066542 -0.972875
+ 2.111e+11Hz -0.0672857 -0.97281
+ 2.112e+11Hz -0.0680292 -0.972743
+ 2.113e+11Hz -0.0687726 -0.972676
+ 2.114e+11Hz -0.0695157 -0.972608
+ 2.115e+11Hz -0.0702587 -0.97254
+ 2.116e+11Hz -0.0710014 -0.972471
+ 2.117e+11Hz -0.071744 -0.972401
+ 2.118e+11Hz -0.0724863 -0.972331
+ 2.119e+11Hz -0.0732284 -0.97226
+ 2.12e+11Hz -0.0739704 -0.972189
+ 2.121e+11Hz -0.0747121 -0.972116
+ 2.122e+11Hz -0.0754535 -0.972044
+ 2.123e+11Hz -0.0761948 -0.97197
+ 2.124e+11Hz -0.0769359 -0.971897
+ 2.125e+11Hz -0.0776767 -0.971822
+ 2.126e+11Hz -0.0784173 -0.971747
+ 2.127e+11Hz -0.0791577 -0.971671
+ 2.128e+11Hz -0.0798978 -0.971595
+ 2.129e+11Hz -0.0806377 -0.971518
+ 2.13e+11Hz -0.0813774 -0.971441
+ 2.131e+11Hz -0.0821168 -0.971363
+ 2.132e+11Hz -0.082856 -0.971284
+ 2.133e+11Hz -0.0835949 -0.971205
+ 2.134e+11Hz -0.0843336 -0.971125
+ 2.135e+11Hz -0.0850721 -0.971045
+ 2.136e+11Hz -0.0858103 -0.970964
+ 2.137e+11Hz -0.0865482 -0.970883
+ 2.138e+11Hz -0.0872859 -0.970801
+ 2.139e+11Hz -0.0880233 -0.970718
+ 2.14e+11Hz -0.0887605 -0.970635
+ 2.141e+11Hz -0.0894975 -0.970552
+ 2.142e+11Hz -0.0902341 -0.970468
+ 2.143e+11Hz -0.0909705 -0.970383
+ 2.144e+11Hz -0.0917067 -0.970298
+ 2.145e+11Hz -0.0924426 -0.970212
+ 2.146e+11Hz -0.0931782 -0.970126
+ 2.147e+11Hz -0.0939135 -0.970039
+ 2.148e+11Hz -0.0946486 -0.969952
+ 2.149e+11Hz -0.0953834 -0.969864
+ 2.15e+11Hz -0.096118 -0.969776
+ 2.151e+11Hz -0.0968523 -0.969687
+ 2.152e+11Hz -0.0975863 -0.969597
+ 2.153e+11Hz -0.09832 -0.969508
+ 2.154e+11Hz -0.0990535 -0.969417
+ 2.155e+11Hz -0.0997867 -0.969327
+ 2.156e+11Hz -0.10052 -0.969235
+ 2.157e+11Hz -0.101252 -0.969144
+ 2.158e+11Hz -0.101985 -0.969051
+ 2.159e+11Hz -0.102717 -0.968959
+ 2.16e+11Hz -0.103449 -0.968866
+ 2.161e+11Hz -0.10418 -0.968772
+ 2.162e+11Hz -0.104911 -0.968678
+ 2.163e+11Hz -0.105642 -0.968583
+ 2.164e+11Hz -0.106373 -0.968488
+ 2.165e+11Hz -0.107104 -0.968393
+ 2.166e+11Hz -0.107834 -0.968297
+ 2.167e+11Hz -0.108564 -0.968201
+ 2.168e+11Hz -0.109293 -0.968104
+ 2.169e+11Hz -0.110023 -0.968007
+ 2.17e+11Hz -0.110752 -0.96791
+ 2.171e+11Hz -0.111481 -0.967812
+ 2.172e+11Hz -0.112209 -0.967713
+ 2.173e+11Hz -0.112937 -0.967615
+ 2.174e+11Hz -0.113666 -0.967515
+ 2.175e+11Hz -0.114393 -0.967416
+ 2.176e+11Hz -0.115121 -0.967316
+ 2.177e+11Hz -0.115848 -0.967216
+ 2.178e+11Hz -0.116575 -0.967115
+ 2.179e+11Hz -0.117302 -0.967014
+ 2.18e+11Hz -0.118028 -0.966912
+ 2.181e+11Hz -0.118754 -0.96681
+ 2.182e+11Hz -0.11948 -0.966708
+ 2.183e+11Hz -0.120206 -0.966606
+ 2.184e+11Hz -0.120932 -0.966503
+ 2.185e+11Hz -0.121657 -0.966399
+ 2.186e+11Hz -0.122382 -0.966296
+ 2.187e+11Hz -0.123106 -0.966192
+ 2.188e+11Hz -0.123831 -0.966087
+ 2.189e+11Hz -0.124555 -0.965983
+ 2.19e+11Hz -0.125279 -0.965878
+ 2.191e+11Hz -0.126003 -0.965772
+ 2.192e+11Hz -0.126727 -0.965667
+ 2.193e+11Hz -0.12745 -0.965561
+ 2.194e+11Hz -0.128173 -0.965454
+ 2.195e+11Hz -0.128896 -0.965348
+ 2.196e+11Hz -0.129619 -0.965241
+ 2.197e+11Hz -0.130341 -0.965134
+ 2.198e+11Hz -0.131063 -0.965026
+ 2.199e+11Hz -0.131786 -0.964918
+ 2.2e+11Hz -0.132507 -0.96481
+ 2.201e+11Hz -0.133229 -0.964702
+ 2.202e+11Hz -0.133951 -0.964593
+ 2.203e+11Hz -0.134672 -0.964484
+ 2.204e+11Hz -0.135393 -0.964375
+ 2.205e+11Hz -0.136114 -0.964265
+ 2.206e+11Hz -0.136835 -0.964155
+ 2.207e+11Hz -0.137555 -0.964045
+ 2.208e+11Hz -0.138275 -0.963935
+ 2.209e+11Hz -0.138996 -0.963824
+ 2.21e+11Hz -0.139716 -0.963713
+ 2.211e+11Hz -0.140436 -0.963602
+ 2.212e+11Hz -0.141155 -0.963491
+ 2.213e+11Hz -0.141875 -0.963379
+ 2.214e+11Hz -0.142594 -0.963267
+ 2.215e+11Hz -0.143314 -0.963155
+ 2.216e+11Hz -0.144033 -0.963042
+ 2.217e+11Hz -0.144752 -0.96293
+ 2.218e+11Hz -0.145471 -0.962817
+ 2.219e+11Hz -0.14619 -0.962703
+ 2.22e+11Hz -0.146908 -0.96259
+ 2.221e+11Hz -0.147627 -0.962476
+ 2.222e+11Hz -0.148346 -0.962362
+ 2.223e+11Hz -0.149064 -0.962248
+ 2.224e+11Hz -0.149782 -0.962134
+ 2.225e+11Hz -0.1505 -0.962019
+ 2.226e+11Hz -0.151219 -0.961904
+ 2.227e+11Hz -0.151937 -0.961789
+ 2.228e+11Hz -0.152655 -0.961673
+ 2.229e+11Hz -0.153372 -0.961558
+ 2.23e+11Hz -0.15409 -0.961442
+ 2.231e+11Hz -0.154808 -0.961326
+ 2.232e+11Hz -0.155526 -0.96121
+ 2.233e+11Hz -0.156243 -0.961093
+ 2.234e+11Hz -0.156961 -0.960976
+ 2.235e+11Hz -0.157679 -0.960859
+ 2.236e+11Hz -0.158396 -0.960742
+ 2.237e+11Hz -0.159114 -0.960625
+ 2.238e+11Hz -0.159831 -0.960507
+ 2.239e+11Hz -0.160549 -0.960389
+ 2.24e+11Hz -0.161266 -0.960271
+ 2.241e+11Hz -0.161984 -0.960152
+ 2.242e+11Hz -0.162701 -0.960034
+ 2.243e+11Hz -0.163419 -0.959915
+ 2.244e+11Hz -0.164136 -0.959796
+ 2.245e+11Hz -0.164854 -0.959677
+ 2.246e+11Hz -0.165571 -0.959557
+ 2.247e+11Hz -0.166289 -0.959437
+ 2.248e+11Hz -0.167006 -0.959317
+ 2.249e+11Hz -0.167724 -0.959197
+ 2.25e+11Hz -0.168442 -0.959076
+ 2.251e+11Hz -0.169159 -0.958955
+ 2.252e+11Hz -0.169877 -0.958834
+ 2.253e+11Hz -0.170595 -0.958713
+ 2.254e+11Hz -0.171313 -0.958592
+ 2.255e+11Hz -0.172031 -0.95847
+ 2.256e+11Hz -0.172749 -0.958348
+ 2.257e+11Hz -0.173467 -0.958225
+ 2.258e+11Hz -0.174185 -0.958103
+ 2.259e+11Hz -0.174904 -0.95798
+ 2.26e+11Hz -0.175622 -0.957857
+ 2.261e+11Hz -0.176341 -0.957734
+ 2.262e+11Hz -0.177059 -0.95761
+ 2.263e+11Hz -0.177778 -0.957486
+ 2.264e+11Hz -0.178497 -0.957362
+ 2.265e+11Hz -0.179216 -0.957238
+ 2.266e+11Hz -0.179935 -0.957113
+ 2.267e+11Hz -0.180654 -0.956988
+ 2.268e+11Hz -0.181374 -0.956862
+ 2.269e+11Hz -0.182093 -0.956737
+ 2.27e+11Hz -0.182813 -0.956611
+ 2.271e+11Hz -0.183533 -0.956485
+ 2.272e+11Hz -0.184252 -0.956358
+ 2.273e+11Hz -0.184973 -0.956231
+ 2.274e+11Hz -0.185693 -0.956104
+ 2.275e+11Hz -0.186413 -0.955977
+ 2.276e+11Hz -0.187134 -0.955849
+ 2.277e+11Hz -0.187855 -0.955721
+ 2.278e+11Hz -0.188576 -0.955592
+ 2.279e+11Hz -0.189297 -0.955464
+ 2.28e+11Hz -0.190018 -0.955335
+ 2.281e+11Hz -0.19074 -0.955205
+ 2.282e+11Hz -0.191461 -0.955075
+ 2.283e+11Hz -0.192183 -0.954945
+ 2.284e+11Hz -0.192905 -0.954815
+ 2.285e+11Hz -0.193627 -0.954684
+ 2.286e+11Hz -0.19435 -0.954552
+ 2.287e+11Hz -0.195073 -0.954421
+ 2.288e+11Hz -0.195796 -0.954289
+ 2.289e+11Hz -0.196519 -0.954156
+ 2.29e+11Hz -0.197242 -0.954023
+ 2.291e+11Hz -0.197965 -0.95389
+ 2.292e+11Hz -0.198689 -0.953757
+ 2.293e+11Hz -0.199413 -0.953623
+ 2.294e+11Hz -0.200137 -0.953488
+ 2.295e+11Hz -0.200862 -0.953353
+ 2.296e+11Hz -0.201587 -0.953218
+ 2.297e+11Hz -0.202311 -0.953082
+ 2.298e+11Hz -0.203037 -0.952946
+ 2.299e+11Hz -0.203762 -0.95281
+ 2.3e+11Hz -0.204487 -0.952673
+ 2.301e+11Hz -0.205213 -0.952535
+ 2.302e+11Hz -0.205939 -0.952397
+ 2.303e+11Hz -0.206666 -0.952259
+ 2.304e+11Hz -0.207392 -0.95212
+ 2.305e+11Hz -0.208119 -0.95198
+ 2.306e+11Hz -0.208846 -0.951841
+ 2.307e+11Hz -0.209573 -0.9517
+ 2.308e+11Hz -0.210301 -0.951559
+ 2.309e+11Hz -0.211029 -0.951418
+ 2.31e+11Hz -0.211757 -0.951276
+ 2.311e+11Hz -0.212485 -0.951134
+ 2.312e+11Hz -0.213213 -0.950991
+ 2.313e+11Hz -0.213942 -0.950848
+ 2.314e+11Hz -0.214671 -0.950704
+ 2.315e+11Hz -0.2154 -0.950559
+ 2.316e+11Hz -0.21613 -0.950414
+ 2.317e+11Hz -0.21686 -0.950268
+ 2.318e+11Hz -0.21759 -0.950122
+ 2.319e+11Hz -0.21832 -0.949976
+ 2.32e+11Hz -0.21905 -0.949828
+ 2.321e+11Hz -0.219781 -0.94968
+ 2.322e+11Hz -0.220512 -0.949532
+ 2.323e+11Hz -0.221243 -0.949383
+ 2.324e+11Hz -0.221974 -0.949233
+ 2.325e+11Hz -0.222706 -0.949083
+ 2.326e+11Hz -0.223438 -0.948932
+ 2.327e+11Hz -0.22417 -0.948781
+ 2.328e+11Hz -0.224902 -0.948629
+ 2.329e+11Hz -0.225635 -0.948476
+ 2.33e+11Hz -0.226368 -0.948323
+ 2.331e+11Hz -0.227101 -0.948169
+ 2.332e+11Hz -0.227834 -0.948014
+ 2.333e+11Hz -0.228568 -0.947859
+ 2.334e+11Hz -0.229301 -0.947703
+ 2.335e+11Hz -0.230035 -0.947546
+ 2.336e+11Hz -0.230769 -0.947389
+ 2.337e+11Hz -0.231504 -0.947231
+ 2.338e+11Hz -0.232238 -0.947073
+ 2.339e+11Hz -0.232973 -0.946913
+ 2.34e+11Hz -0.233708 -0.946753
+ 2.341e+11Hz -0.234443 -0.946593
+ 2.342e+11Hz -0.235178 -0.946431
+ 2.343e+11Hz -0.235914 -0.946269
+ 2.344e+11Hz -0.23665 -0.946107
+ 2.345e+11Hz -0.237385 -0.945943
+ 2.346e+11Hz -0.238122 -0.945779
+ 2.347e+11Hz -0.238858 -0.945614
+ 2.348e+11Hz -0.239594 -0.945448
+ 2.349e+11Hz -0.240331 -0.945282
+ 2.35e+11Hz -0.241068 -0.945115
+ 2.351e+11Hz -0.241805 -0.944947
+ 2.352e+11Hz -0.242542 -0.944778
+ 2.353e+11Hz -0.243279 -0.944609
+ 2.354e+11Hz -0.244016 -0.944439
+ 2.355e+11Hz -0.244754 -0.944268
+ 2.356e+11Hz -0.245491 -0.944096
+ 2.357e+11Hz -0.246229 -0.943924
+ 2.358e+11Hz -0.246967 -0.943751
+ 2.359e+11Hz -0.247705 -0.943577
+ 2.36e+11Hz -0.248443 -0.943402
+ 2.361e+11Hz -0.249182 -0.943227
+ 2.362e+11Hz -0.24992 -0.94305
+ 2.363e+11Hz -0.250659 -0.942873
+ 2.364e+11Hz -0.251397 -0.942695
+ 2.365e+11Hz -0.252136 -0.942517
+ 2.366e+11Hz -0.252875 -0.942337
+ 2.367e+11Hz -0.253614 -0.942157
+ 2.368e+11Hz -0.254353 -0.941976
+ 2.369e+11Hz -0.255092 -0.941794
+ 2.37e+11Hz -0.255831 -0.941611
+ 2.371e+11Hz -0.25657 -0.941427
+ 2.372e+11Hz -0.257309 -0.941243
+ 2.373e+11Hz -0.258049 -0.941058
+ 2.374e+11Hz -0.258788 -0.940872
+ 2.375e+11Hz -0.259527 -0.940685
+ 2.376e+11Hz -0.260267 -0.940497
+ 2.377e+11Hz -0.261006 -0.940309
+ 2.378e+11Hz -0.261746 -0.94012
+ 2.379e+11Hz -0.262485 -0.93993
+ 2.38e+11Hz -0.263225 -0.939739
+ 2.381e+11Hz -0.263964 -0.939547
+ 2.382e+11Hz -0.264704 -0.939354
+ 2.383e+11Hz -0.265443 -0.939161
+ 2.384e+11Hz -0.266183 -0.938966
+ 2.385e+11Hz -0.266923 -0.938771
+ 2.386e+11Hz -0.267662 -0.938575
+ 2.387e+11Hz -0.268402 -0.938378
+ 2.388e+11Hz -0.269141 -0.938181
+ 2.389e+11Hz -0.26988 -0.937982
+ 2.39e+11Hz -0.27062 -0.937783
+ 2.391e+11Hz -0.271359 -0.937582
+ 2.392e+11Hz -0.272098 -0.937381
+ 2.393e+11Hz -0.272838 -0.937179
+ 2.394e+11Hz -0.273577 -0.936976
+ 2.395e+11Hz -0.274316 -0.936773
+ 2.396e+11Hz -0.275055 -0.936568
+ 2.397e+11Hz -0.275794 -0.936363
+ 2.398e+11Hz -0.276533 -0.936157
+ 2.399e+11Hz -0.277272 -0.93595
+ 2.4e+11Hz -0.27801 -0.935742
+ 2.401e+11Hz -0.278749 -0.935533
+ 2.402e+11Hz -0.279487 -0.935324
+ 2.403e+11Hz -0.280226 -0.935113
+ 2.404e+11Hz -0.280964 -0.934902
+ 2.405e+11Hz -0.281702 -0.93469
+ 2.406e+11Hz -0.28244 -0.934477
+ 2.407e+11Hz -0.283178 -0.934263
+ 2.408e+11Hz -0.283916 -0.934048
+ 2.409e+11Hz -0.284653 -0.933833
+ 2.41e+11Hz -0.285391 -0.933617
+ 2.411e+11Hz -0.286128 -0.933399
+ 2.412e+11Hz -0.286865 -0.933181
+ 2.413e+11Hz -0.287602 -0.932963
+ 2.414e+11Hz -0.288339 -0.932743
+ 2.415e+11Hz -0.289076 -0.932522
+ 2.416e+11Hz -0.289812 -0.932301
+ 2.417e+11Hz -0.290549 -0.932079
+ 2.418e+11Hz -0.291285 -0.931856
+ 2.419e+11Hz -0.292021 -0.931632
+ 2.42e+11Hz -0.292756 -0.931407
+ 2.421e+11Hz -0.293492 -0.931182
+ 2.422e+11Hz -0.294227 -0.930956
+ 2.423e+11Hz -0.294962 -0.930728
+ 2.424e+11Hz -0.295697 -0.930501
+ 2.425e+11Hz -0.296432 -0.930272
+ 2.426e+11Hz -0.297166 -0.930042
+ 2.427e+11Hz -0.297901 -0.929812
+ 2.428e+11Hz -0.298635 -0.929581
+ 2.429e+11Hz -0.299368 -0.929349
+ 2.43e+11Hz -0.300102 -0.929116
+ 2.431e+11Hz -0.300835 -0.928882
+ 2.432e+11Hz -0.301568 -0.928648
+ 2.433e+11Hz -0.302301 -0.928413
+ 2.434e+11Hz -0.303034 -0.928177
+ 2.435e+11Hz -0.303766 -0.92794
+ 2.436e+11Hz -0.304498 -0.927703
+ 2.437e+11Hz -0.30523 -0.927464
+ 2.438e+11Hz -0.305962 -0.927225
+ 2.439e+11Hz -0.306693 -0.926985
+ 2.44e+11Hz -0.307424 -0.926745
+ 2.441e+11Hz -0.308155 -0.926503
+ 2.442e+11Hz -0.308885 -0.926261
+ 2.443e+11Hz -0.309616 -0.926018
+ 2.444e+11Hz -0.310345 -0.925774
+ 2.445e+11Hz -0.311075 -0.92553
+ 2.446e+11Hz -0.311805 -0.925285
+ 2.447e+11Hz -0.312534 -0.925039
+ 2.448e+11Hz -0.313262 -0.924792
+ 2.449e+11Hz -0.313991 -0.924545
+ 2.45e+11Hz -0.314719 -0.924296
+ 2.451e+11Hz -0.315447 -0.924047
+ 2.452e+11Hz -0.316175 -0.923798
+ 2.453e+11Hz -0.316902 -0.923547
+ 2.454e+11Hz -0.317629 -0.923296
+ 2.455e+11Hz -0.318356 -0.923044
+ 2.456e+11Hz -0.319082 -0.922791
+ 2.457e+11Hz -0.319808 -0.922538
+ 2.458e+11Hz -0.320534 -0.922284
+ 2.459e+11Hz -0.321259 -0.922029
+ 2.46e+11Hz -0.321985 -0.921774
+ 2.461e+11Hz -0.32271 -0.921517
+ 2.462e+11Hz -0.323434 -0.92126
+ 2.463e+11Hz -0.324158 -0.921003
+ 2.464e+11Hz -0.324882 -0.920744
+ 2.465e+11Hz -0.325606 -0.920485
+ 2.466e+11Hz -0.326329 -0.920225
+ 2.467e+11Hz -0.327052 -0.919965
+ 2.468e+11Hz -0.327775 -0.919704
+ 2.469e+11Hz -0.328497 -0.919442
+ 2.47e+11Hz -0.329219 -0.919179
+ 2.471e+11Hz -0.329941 -0.918916
+ 2.472e+11Hz -0.330662 -0.918652
+ 2.473e+11Hz -0.331383 -0.918388
+ 2.474e+11Hz -0.332103 -0.918122
+ 2.475e+11Hz -0.332824 -0.917856
+ 2.476e+11Hz -0.333544 -0.91759
+ 2.477e+11Hz -0.334264 -0.917322
+ 2.478e+11Hz -0.334983 -0.917054
+ 2.479e+11Hz -0.335702 -0.916786
+ 2.48e+11Hz -0.336421 -0.916516
+ 2.481e+11Hz -0.337139 -0.916247
+ 2.482e+11Hz -0.337857 -0.915976
+ 2.483e+11Hz -0.338575 -0.915705
+ 2.484e+11Hz -0.339292 -0.915433
+ 2.485e+11Hz -0.340009 -0.91516
+ 2.486e+11Hz -0.340726 -0.914887
+ 2.487e+11Hz -0.341442 -0.914613
+ 2.488e+11Hz -0.342158 -0.914338
+ 2.489e+11Hz -0.342874 -0.914063
+ 2.49e+11Hz -0.343589 -0.913787
+ 2.491e+11Hz -0.344304 -0.913511
+ 2.492e+11Hz -0.345019 -0.913234
+ 2.493e+11Hz -0.345733 -0.912956
+ 2.494e+11Hz -0.346447 -0.912678
+ 2.495e+11Hz -0.347161 -0.912399
+ 2.496e+11Hz -0.347874 -0.912119
+ 2.497e+11Hz -0.348587 -0.911839
+ 2.498e+11Hz -0.3493 -0.911558
+ 2.499e+11Hz -0.350012 -0.911276
+ 2.5e+11Hz -0.350724 -0.910994
+ 2.501e+11Hz -0.351436 -0.910712
+ 2.502e+11Hz -0.352147 -0.910428
+ 2.503e+11Hz -0.352858 -0.910144
+ 2.504e+11Hz -0.353569 -0.909859
+ 2.505e+11Hz -0.354279 -0.909574
+ 2.506e+11Hz -0.354989 -0.909288
+ 2.507e+11Hz -0.355699 -0.909002
+ 2.508e+11Hz -0.356408 -0.908715
+ 2.509e+11Hz -0.357117 -0.908427
+ 2.51e+11Hz -0.357826 -0.908139
+ 2.511e+11Hz -0.358534 -0.90785
+ 2.512e+11Hz -0.359242 -0.90756
+ 2.513e+11Hz -0.35995 -0.90727
+ 2.514e+11Hz -0.360657 -0.906979
+ 2.515e+11Hz -0.361364 -0.906688
+ 2.516e+11Hz -0.36207 -0.906396
+ 2.517e+11Hz -0.362777 -0.906103
+ 2.518e+11Hz -0.363483 -0.90581
+ 2.519e+11Hz -0.364188 -0.905516
+ 2.52e+11Hz -0.364894 -0.905221
+ 2.521e+11Hz -0.365598 -0.904926
+ 2.522e+11Hz -0.366303 -0.904631
+ 2.523e+11Hz -0.367007 -0.904334
+ 2.524e+11Hz -0.367711 -0.904038
+ 2.525e+11Hz -0.368415 -0.90374
+ 2.526e+11Hz -0.369118 -0.903442
+ 2.527e+11Hz -0.369821 -0.903143
+ 2.528e+11Hz -0.370523 -0.902844
+ 2.529e+11Hz -0.371226 -0.902544
+ 2.53e+11Hz -0.371928 -0.902244
+ 2.531e+11Hz -0.372629 -0.901943
+ 2.532e+11Hz -0.37333 -0.901641
+ 2.533e+11Hz -0.374031 -0.901339
+ 2.534e+11Hz -0.374732 -0.901036
+ 2.535e+11Hz -0.375432 -0.900732
+ 2.536e+11Hz -0.376131 -0.900428
+ 2.537e+11Hz -0.376831 -0.900123
+ 2.538e+11Hz -0.37753 -0.899818
+ 2.539e+11Hz -0.378229 -0.899512
+ 2.54e+11Hz -0.378927 -0.899206
+ 2.541e+11Hz -0.379625 -0.898899
+ 2.542e+11Hz -0.380323 -0.898591
+ 2.543e+11Hz -0.38102 -0.898283
+ 2.544e+11Hz -0.381717 -0.897974
+ 2.545e+11Hz -0.382414 -0.897664
+ 2.546e+11Hz -0.38311 -0.897354
+ 2.547e+11Hz -0.383806 -0.897044
+ 2.548e+11Hz -0.384502 -0.896732
+ 2.549e+11Hz -0.385197 -0.896421
+ 2.55e+11Hz -0.385892 -0.896108
+ 2.551e+11Hz -0.386586 -0.895795
+ 2.552e+11Hz -0.38728 -0.895481
+ 2.553e+11Hz -0.387974 -0.895167
+ 2.554e+11Hz -0.388667 -0.894852
+ 2.555e+11Hz -0.38936 -0.894537
+ 2.556e+11Hz -0.390053 -0.894221
+ 2.557e+11Hz -0.390745 -0.893904
+ 2.558e+11Hz -0.391437 -0.893587
+ 2.559e+11Hz -0.392128 -0.893269
+ 2.56e+11Hz -0.392819 -0.892951
+ 2.561e+11Hz -0.39351 -0.892632
+ 2.562e+11Hz -0.3942 -0.892312
+ 2.563e+11Hz -0.39489 -0.891992
+ 2.564e+11Hz -0.39558 -0.891672
+ 2.565e+11Hz -0.396269 -0.89135
+ 2.566e+11Hz -0.396958 -0.891028
+ 2.567e+11Hz -0.397646 -0.890706
+ 2.568e+11Hz -0.398334 -0.890383
+ 2.569e+11Hz -0.399022 -0.890059
+ 2.57e+11Hz -0.399709 -0.889735
+ 2.571e+11Hz -0.400396 -0.88941
+ 2.572e+11Hz -0.401082 -0.889085
+ 2.573e+11Hz -0.401768 -0.888759
+ 2.574e+11Hz -0.402454 -0.888432
+ 2.575e+11Hz -0.403139 -0.888105
+ 2.576e+11Hz -0.403824 -0.887778
+ 2.577e+11Hz -0.404508 -0.887449
+ 2.578e+11Hz -0.405192 -0.887121
+ 2.579e+11Hz -0.405875 -0.886791
+ 2.58e+11Hz -0.406558 -0.886461
+ 2.581e+11Hz -0.407241 -0.886131
+ 2.582e+11Hz -0.407923 -0.8858
+ 2.583e+11Hz -0.408605 -0.885468
+ 2.584e+11Hz -0.409286 -0.885136
+ 2.585e+11Hz -0.409967 -0.884803
+ 2.586e+11Hz -0.410648 -0.88447
+ 2.587e+11Hz -0.411328 -0.884136
+ 2.588e+11Hz -0.412007 -0.883802
+ 2.589e+11Hz -0.412686 -0.883467
+ 2.59e+11Hz -0.413365 -0.883131
+ 2.591e+11Hz -0.414043 -0.882795
+ 2.592e+11Hz -0.414721 -0.882458
+ 2.593e+11Hz -0.415398 -0.882121
+ 2.594e+11Hz -0.416075 -0.881784
+ 2.595e+11Hz -0.416752 -0.881446
+ 2.596e+11Hz -0.417428 -0.881107
+ 2.597e+11Hz -0.418103 -0.880768
+ 2.598e+11Hz -0.418778 -0.880428
+ 2.599e+11Hz -0.419453 -0.880088
+ 2.6e+11Hz -0.420127 -0.879747
+ 2.601e+11Hz -0.420801 -0.879405
+ 2.602e+11Hz -0.421474 -0.879064
+ 2.603e+11Hz -0.422146 -0.878721
+ 2.604e+11Hz -0.422819 -0.878379
+ 2.605e+11Hz -0.42349 -0.878035
+ 2.606e+11Hz -0.424162 -0.877691
+ 2.607e+11Hz -0.424832 -0.877347
+ 2.608e+11Hz -0.425503 -0.877002
+ 2.609e+11Hz -0.426173 -0.876657
+ 2.61e+11Hz -0.426842 -0.876311
+ 2.611e+11Hz -0.427511 -0.875965
+ 2.612e+11Hz -0.428179 -0.875618
+ 2.613e+11Hz -0.428847 -0.875271
+ 2.614e+11Hz -0.429514 -0.874923
+ 2.615e+11Hz -0.430181 -0.874575
+ 2.616e+11Hz -0.430847 -0.874227
+ 2.617e+11Hz -0.431513 -0.873878
+ 2.618e+11Hz -0.432179 -0.873528
+ 2.619e+11Hz -0.432843 -0.873178
+ 2.62e+11Hz -0.433508 -0.872828
+ 2.621e+11Hz -0.434172 -0.872477
+ 2.622e+11Hz -0.434835 -0.872126
+ 2.623e+11Hz -0.435498 -0.871774
+ 2.624e+11Hz -0.43616 -0.871422
+ 2.625e+11Hz -0.436822 -0.87107
+ 2.626e+11Hz -0.437484 -0.870717
+ 2.627e+11Hz -0.438144 -0.870364
+ 2.628e+11Hz -0.438805 -0.87001
+ 2.629e+11Hz -0.439465 -0.869656
+ 2.63e+11Hz -0.440124 -0.869301
+ 2.631e+11Hz -0.440783 -0.868947
+ 2.632e+11Hz -0.441441 -0.868591
+ 2.633e+11Hz -0.442099 -0.868236
+ 2.634e+11Hz -0.442756 -0.86788
+ 2.635e+11Hz -0.443413 -0.867523
+ 2.636e+11Hz -0.444069 -0.867167
+ 2.637e+11Hz -0.444725 -0.86681
+ 2.638e+11Hz -0.44538 -0.866452
+ 2.639e+11Hz -0.446035 -0.866094
+ 2.64e+11Hz -0.44669 -0.865736
+ 2.641e+11Hz -0.447343 -0.865378
+ 2.642e+11Hz -0.447997 -0.865019
+ 2.643e+11Hz -0.448649 -0.86466
+ 2.644e+11Hz -0.449302 -0.8643
+ 2.645e+11Hz -0.449954 -0.863941
+ 2.646e+11Hz -0.450605 -0.863581
+ 2.647e+11Hz -0.451256 -0.86322
+ 2.648e+11Hz -0.451906 -0.86286
+ 2.649e+11Hz -0.452556 -0.862499
+ 2.65e+11Hz -0.453205 -0.862137
+ 2.651e+11Hz -0.453854 -0.861776
+ 2.652e+11Hz -0.454503 -0.861414
+ 2.653e+11Hz -0.455151 -0.861052
+ 2.654e+11Hz -0.455798 -0.86069
+ 2.655e+11Hz -0.456445 -0.860327
+ 2.656e+11Hz -0.457092 -0.859964
+ 2.657e+11Hz -0.457738 -0.859601
+ 2.658e+11Hz -0.458384 -0.859238
+ 2.659e+11Hz -0.459029 -0.858874
+ 2.66e+11Hz -0.459673 -0.85851
+ 2.661e+11Hz -0.460318 -0.858146
+ 2.662e+11Hz -0.460962 -0.857782
+ 2.663e+11Hz -0.461605 -0.857418
+ 2.664e+11Hz -0.462248 -0.857053
+ 2.665e+11Hz -0.46289 -0.856688
+ 2.666e+11Hz -0.463532 -0.856323
+ 2.667e+11Hz -0.464174 -0.855957
+ 2.668e+11Hz -0.464815 -0.855592
+ 2.669e+11Hz -0.465456 -0.855226
+ 2.67e+11Hz -0.466097 -0.85486
+ 2.671e+11Hz -0.466737 -0.854494
+ 2.672e+11Hz -0.467376 -0.854128
+ 2.673e+11Hz -0.468015 -0.853761
+ 2.674e+11Hz -0.468654 -0.853395
+ 2.675e+11Hz -0.469293 -0.853028
+ 2.676e+11Hz -0.469931 -0.852661
+ 2.677e+11Hz -0.470568 -0.852293
+ 2.678e+11Hz -0.471205 -0.851926
+ 2.679e+11Hz -0.471842 -0.851559
+ 2.68e+11Hz -0.472479 -0.851191
+ 2.681e+11Hz -0.473115 -0.850823
+ 2.682e+11Hz -0.473751 -0.850455
+ 2.683e+11Hz -0.474386 -0.850087
+ 2.684e+11Hz -0.475022 -0.849719
+ 2.685e+11Hz -0.475656 -0.849351
+ 2.686e+11Hz -0.476291 -0.848982
+ 2.687e+11Hz -0.476925 -0.848613
+ 2.688e+11Hz -0.477559 -0.848245
+ 2.689e+11Hz -0.478193 -0.847876
+ 2.69e+11Hz -0.478826 -0.847507
+ 2.691e+11Hz -0.479459 -0.847138
+ 2.692e+11Hz -0.480091 -0.846768
+ 2.693e+11Hz -0.480724 -0.846399
+ 2.694e+11Hz -0.481356 -0.846029
+ 2.695e+11Hz -0.481988 -0.84566
+ 2.696e+11Hz -0.482619 -0.84529
+ 2.697e+11Hz -0.483251 -0.84492
+ 2.698e+11Hz -0.483882 -0.84455
+ 2.699e+11Hz -0.484513 -0.84418
+ 2.7e+11Hz -0.485143 -0.84381
+ 2.701e+11Hz -0.485774 -0.84344
+ 2.702e+11Hz -0.486404 -0.843069
+ 2.703e+11Hz -0.487034 -0.842699
+ 2.704e+11Hz -0.487664 -0.842328
+ 2.705e+11Hz -0.488293 -0.841957
+ 2.706e+11Hz -0.488923 -0.841586
+ 2.707e+11Hz -0.489552 -0.841215
+ 2.708e+11Hz -0.490181 -0.840844
+ 2.709e+11Hz -0.49081 -0.840473
+ 2.71e+11Hz -0.491439 -0.840102
+ 2.711e+11Hz -0.492067 -0.83973
+ 2.712e+11Hz -0.492696 -0.839359
+ 2.713e+11Hz -0.493324 -0.838987
+ 2.714e+11Hz -0.493952 -0.838615
+ 2.715e+11Hz -0.49458 -0.838243
+ 2.716e+11Hz -0.495208 -0.837871
+ 2.717e+11Hz -0.495836 -0.837499
+ 2.718e+11Hz -0.496464 -0.837127
+ 2.719e+11Hz -0.497092 -0.836754
+ 2.72e+11Hz -0.497719 -0.836382
+ 2.721e+11Hz -0.498347 -0.836009
+ 2.722e+11Hz -0.498974 -0.835636
+ 2.723e+11Hz -0.499601 -0.835263
+ 2.724e+11Hz -0.500229 -0.83489
+ 2.725e+11Hz -0.500856 -0.834517
+ 2.726e+11Hz -0.501483 -0.834144
+ 2.727e+11Hz -0.50211 -0.83377
+ 2.728e+11Hz -0.502738 -0.833396
+ 2.729e+11Hz -0.503365 -0.833022
+ 2.73e+11Hz -0.503992 -0.832648
+ 2.731e+11Hz -0.504619 -0.832274
+ 2.732e+11Hz -0.505246 -0.8319
+ 2.733e+11Hz -0.505873 -0.831525
+ 2.734e+11Hz -0.5065 -0.83115
+ 2.735e+11Hz -0.507127 -0.830775
+ 2.736e+11Hz -0.507755 -0.8304
+ 2.737e+11Hz -0.508382 -0.830025
+ 2.738e+11Hz -0.509009 -0.829649
+ 2.739e+11Hz -0.509636 -0.829273
+ 2.74e+11Hz -0.510264 -0.828897
+ 2.741e+11Hz -0.510891 -0.828521
+ 2.742e+11Hz -0.511519 -0.828145
+ 2.743e+11Hz -0.512146 -0.827768
+ 2.744e+11Hz -0.512774 -0.827391
+ 2.745e+11Hz -0.513401 -0.827014
+ 2.746e+11Hz -0.514029 -0.826636
+ 2.747e+11Hz -0.514657 -0.826259
+ 2.748e+11Hz -0.515285 -0.825881
+ 2.749e+11Hz -0.515913 -0.825502
+ 2.75e+11Hz -0.516541 -0.825124
+ 2.751e+11Hz -0.517169 -0.824745
+ 2.752e+11Hz -0.517798 -0.824366
+ 2.753e+11Hz -0.518426 -0.823987
+ 2.754e+11Hz -0.519055 -0.823607
+ 2.755e+11Hz -0.519683 -0.823227
+ 2.756e+11Hz -0.520312 -0.822846
+ 2.757e+11Hz -0.520941 -0.822466
+ 2.758e+11Hz -0.52157 -0.822084
+ 2.759e+11Hz -0.522199 -0.821703
+ 2.76e+11Hz -0.522829 -0.821321
+ 2.761e+11Hz -0.523458 -0.820939
+ 2.762e+11Hz -0.524088 -0.820556
+ 2.763e+11Hz -0.524718 -0.820174
+ 2.764e+11Hz -0.525348 -0.81979
+ 2.765e+11Hz -0.525978 -0.819406
+ 2.766e+11Hz -0.526608 -0.819022
+ 2.767e+11Hz -0.527238 -0.818638
+ 2.768e+11Hz -0.527869 -0.818253
+ 2.769e+11Hz -0.5285 -0.817867
+ 2.77e+11Hz -0.529131 -0.817481
+ 2.771e+11Hz -0.529762 -0.817095
+ 2.772e+11Hz -0.530393 -0.816708
+ 2.773e+11Hz -0.531024 -0.816321
+ 2.774e+11Hz -0.531656 -0.815933
+ 2.775e+11Hz -0.532287 -0.815545
+ 2.776e+11Hz -0.532919 -0.815156
+ 2.777e+11Hz -0.533551 -0.814767
+ 2.778e+11Hz -0.534184 -0.814377
+ 2.779e+11Hz -0.534816 -0.813987
+ 2.78e+11Hz -0.535448 -0.813596
+ 2.781e+11Hz -0.536081 -0.813205
+ 2.782e+11Hz -0.536714 -0.812813
+ 2.783e+11Hz -0.537347 -0.81242
+ 2.784e+11Hz -0.53798 -0.812027
+ 2.785e+11Hz -0.538613 -0.811633
+ 2.786e+11Hz -0.539247 -0.811239
+ 2.787e+11Hz -0.53988 -0.810844
+ 2.788e+11Hz -0.540514 -0.810449
+ 2.789e+11Hz -0.541148 -0.810053
+ 2.79e+11Hz -0.541782 -0.809656
+ 2.791e+11Hz -0.542416 -0.809258
+ 2.792e+11Hz -0.54305 -0.80886
+ 2.793e+11Hz -0.543685 -0.808462
+ 2.794e+11Hz -0.544319 -0.808062
+ 2.795e+11Hz -0.544954 -0.807662
+ 2.796e+11Hz -0.545589 -0.807262
+ 2.797e+11Hz -0.546224 -0.80686
+ 2.798e+11Hz -0.546859 -0.806458
+ 2.799e+11Hz -0.547494 -0.806055
+ 2.8e+11Hz -0.548129 -0.805652
+ 2.801e+11Hz -0.548765 -0.805248
+ 2.802e+11Hz -0.5494 -0.804843
+ 2.803e+11Hz -0.550036 -0.804437
+ 2.804e+11Hz -0.550671 -0.804031
+ 2.805e+11Hz -0.551307 -0.803623
+ 2.806e+11Hz -0.551943 -0.803215
+ 2.807e+11Hz -0.552579 -0.802807
+ 2.808e+11Hz -0.553215 -0.802397
+ 2.809e+11Hz -0.553851 -0.801987
+ 2.81e+11Hz -0.554487 -0.801576
+ 2.811e+11Hz -0.555123 -0.801164
+ 2.812e+11Hz -0.555759 -0.800751
+ 2.813e+11Hz -0.556395 -0.800338
+ 2.814e+11Hz -0.557031 -0.799923
+ 2.815e+11Hz -0.557667 -0.799508
+ 2.816e+11Hz -0.558303 -0.799092
+ 2.817e+11Hz -0.55894 -0.798675
+ 2.818e+11Hz -0.559576 -0.798258
+ 2.819e+11Hz -0.560212 -0.797839
+ 2.82e+11Hz -0.560848 -0.79742
+ 2.821e+11Hz -0.561484 -0.797
+ 2.822e+11Hz -0.56212 -0.796579
+ 2.823e+11Hz -0.562756 -0.796157
+ 2.824e+11Hz -0.563392 -0.795734
+ 2.825e+11Hz -0.564028 -0.79531
+ 2.826e+11Hz -0.564664 -0.794885
+ 2.827e+11Hz -0.5653 -0.79446
+ 2.828e+11Hz -0.565935 -0.794033
+ 2.829e+11Hz -0.566571 -0.793606
+ 2.83e+11Hz -0.567207 -0.793178
+ 2.831e+11Hz -0.567842 -0.792749
+ 2.832e+11Hz -0.568477 -0.792319
+ 2.833e+11Hz -0.569112 -0.791888
+ 2.834e+11Hz -0.569747 -0.791456
+ 2.835e+11Hz -0.570382 -0.791023
+ 2.836e+11Hz -0.571017 -0.790589
+ 2.837e+11Hz -0.571651 -0.790155
+ 2.838e+11Hz -0.572285 -0.789719
+ 2.839e+11Hz -0.572919 -0.789283
+ 2.84e+11Hz -0.573553 -0.788845
+ 2.841e+11Hz -0.574187 -0.788407
+ 2.842e+11Hz -0.57482 -0.787968
+ 2.843e+11Hz -0.575454 -0.787527
+ 2.844e+11Hz -0.576087 -0.787086
+ 2.845e+11Hz -0.57672 -0.786644
+ 2.846e+11Hz -0.577352 -0.786201
+ 2.847e+11Hz -0.577984 -0.785757
+ 2.848e+11Hz -0.578616 -0.785312
+ 2.849e+11Hz -0.579248 -0.784866
+ 2.85e+11Hz -0.579879 -0.784419
+ 2.851e+11Hz -0.58051 -0.783972
+ 2.852e+11Hz -0.581141 -0.783523
+ 2.853e+11Hz -0.581772 -0.783073
+ 2.854e+11Hz -0.582402 -0.782623
+ 2.855e+11Hz -0.583032 -0.782171
+ 2.856e+11Hz -0.583661 -0.781719
+ 2.857e+11Hz -0.58429 -0.781265
+ 2.858e+11Hz -0.584919 -0.780811
+ 2.859e+11Hz -0.585547 -0.780356
+ 2.86e+11Hz -0.586175 -0.779899
+ 2.861e+11Hz -0.586802 -0.779442
+ 2.862e+11Hz -0.58743 -0.778984
+ 2.863e+11Hz -0.588056 -0.778525
+ 2.864e+11Hz -0.588683 -0.778065
+ 2.865e+11Hz -0.589308 -0.777605
+ 2.866e+11Hz -0.589934 -0.777143
+ 2.867e+11Hz -0.590559 -0.77668
+ 2.868e+11Hz -0.591183 -0.776217
+ 2.869e+11Hz -0.591807 -0.775752
+ 2.87e+11Hz -0.592431 -0.775287
+ 2.871e+11Hz -0.593054 -0.77482
+ 2.872e+11Hz -0.593677 -0.774353
+ 2.873e+11Hz -0.594299 -0.773885
+ 2.874e+11Hz -0.59492 -0.773416
+ 2.875e+11Hz -0.595541 -0.772947
+ 2.876e+11Hz -0.596162 -0.772476
+ 2.877e+11Hz -0.596782 -0.772004
+ 2.878e+11Hz -0.597401 -0.771532
+ 2.879e+11Hz -0.59802 -0.771059
+ 2.88e+11Hz -0.598638 -0.770585
+ 2.881e+11Hz -0.599256 -0.77011
+ 2.882e+11Hz -0.599873 -0.769634
+ 2.883e+11Hz -0.60049 -0.769157
+ 2.884e+11Hz -0.601106 -0.76868
+ 2.885e+11Hz -0.601722 -0.768201
+ 2.886e+11Hz -0.602336 -0.767722
+ 2.887e+11Hz -0.602951 -0.767242
+ 2.888e+11Hz -0.603564 -0.766762
+ 2.889e+11Hz -0.604177 -0.76628
+ 2.89e+11Hz -0.60479 -0.765798
+ 2.891e+11Hz -0.605402 -0.765315
+ 2.892e+11Hz -0.606013 -0.764831
+ 2.893e+11Hz -0.606623 -0.764346
+ 2.894e+11Hz -0.607233 -0.763861
+ 2.895e+11Hz -0.607843 -0.763374
+ 2.896e+11Hz -0.608451 -0.762888
+ 2.897e+11Hz -0.609059 -0.7624
+ 2.898e+11Hz -0.609666 -0.761911
+ 2.899e+11Hz -0.610273 -0.761422
+ 2.9e+11Hz -0.610879 -0.760932
+ 2.901e+11Hz -0.611484 -0.760442
+ 2.902e+11Hz -0.612089 -0.759951
+ 2.903e+11Hz -0.612693 -0.759459
+ 2.904e+11Hz -0.613296 -0.758966
+ 2.905e+11Hz -0.613899 -0.758473
+ 2.906e+11Hz -0.614501 -0.757978
+ 2.907e+11Hz -0.615102 -0.757484
+ 2.908e+11Hz -0.615703 -0.756988
+ 2.909e+11Hz -0.616302 -0.756492
+ 2.91e+11Hz -0.616902 -0.755996
+ 2.911e+11Hz -0.6175 -0.755498
+ 2.912e+11Hz -0.618098 -0.755
+ 2.913e+11Hz -0.618695 -0.754502
+ 2.914e+11Hz -0.619291 -0.754003
+ 2.915e+11Hz -0.619887 -0.753503
+ 2.916e+11Hz -0.620482 -0.753003
+ 2.917e+11Hz -0.621076 -0.752502
+ 2.918e+11Hz -0.62167 -0.752
+ 2.919e+11Hz -0.622262 -0.751498
+ 2.92e+11Hz -0.622855 -0.750995
+ 2.921e+11Hz -0.623446 -0.750492
+ 2.922e+11Hz -0.624037 -0.749988
+ 2.923e+11Hz -0.624627 -0.749484
+ 2.924e+11Hz -0.625216 -0.748979
+ 2.925e+11Hz -0.625805 -0.748473
+ 2.926e+11Hz -0.626392 -0.747967
+ 2.927e+11Hz -0.62698 -0.747461
+ 2.928e+11Hz -0.627566 -0.746954
+ 2.929e+11Hz -0.628152 -0.746446
+ 2.93e+11Hz -0.628737 -0.745938
+ 2.931e+11Hz -0.629322 -0.74543
+ 2.932e+11Hz -0.629905 -0.744921
+ 2.933e+11Hz -0.630488 -0.744411
+ 2.934e+11Hz -0.631071 -0.743901
+ 2.935e+11Hz -0.631652 -0.743391
+ 2.936e+11Hz -0.632233 -0.74288
+ 2.937e+11Hz -0.632813 -0.742369
+ 2.938e+11Hz -0.633393 -0.741857
+ 2.939e+11Hz -0.633972 -0.741345
+ 2.94e+11Hz -0.63455 -0.740832
+ 2.941e+11Hz -0.635128 -0.740319
+ 2.942e+11Hz -0.635705 -0.739805
+ 2.943e+11Hz -0.636281 -0.739291
+ 2.944e+11Hz -0.636856 -0.738777
+ 2.945e+11Hz -0.637431 -0.738262
+ 2.946e+11Hz -0.638005 -0.737747
+ 2.947e+11Hz -0.638579 -0.737231
+ 2.948e+11Hz -0.639152 -0.736716
+ 2.949e+11Hz -0.639724 -0.736199
+ 2.95e+11Hz -0.640296 -0.735682
+ 2.951e+11Hz -0.640867 -0.735165
+ 2.952e+11Hz -0.641437 -0.734648
+ 2.953e+11Hz -0.642007 -0.73413
+ 2.954e+11Hz -0.642576 -0.733612
+ 2.955e+11Hz -0.643144 -0.733093
+ 2.956e+11Hz -0.643712 -0.732574
+ 2.957e+11Hz -0.644279 -0.732055
+ 2.958e+11Hz -0.644846 -0.731535
+ 2.959e+11Hz -0.645412 -0.731015
+ 2.96e+11Hz -0.645978 -0.730494
+ 2.961e+11Hz -0.646542 -0.729974
+ 2.962e+11Hz -0.647107 -0.729452
+ 2.963e+11Hz -0.64767 -0.728931
+ 2.964e+11Hz -0.648233 -0.728409
+ 2.965e+11Hz -0.648796 -0.727887
+ 2.966e+11Hz -0.649358 -0.727364
+ 2.967e+11Hz -0.649919 -0.726842
+ 2.968e+11Hz -0.65048 -0.726318
+ 2.969e+11Hz -0.65104 -0.725795
+ 2.97e+11Hz -0.651599 -0.725271
+ 2.971e+11Hz -0.652158 -0.724747
+ 2.972e+11Hz -0.652717 -0.724222
+ 2.973e+11Hz -0.653275 -0.723698
+ 2.974e+11Hz -0.653832 -0.723172
+ 2.975e+11Hz -0.654389 -0.722647
+ 2.976e+11Hz -0.654946 -0.722121
+ 2.977e+11Hz -0.655501 -0.721595
+ 2.978e+11Hz -0.656057 -0.721069
+ 2.979e+11Hz -0.656612 -0.720542
+ 2.98e+11Hz -0.657166 -0.720015
+ 2.981e+11Hz -0.65772 -0.719487
+ 2.982e+11Hz -0.658273 -0.718959
+ 2.983e+11Hz -0.658826 -0.718431
+ 2.984e+11Hz -0.659378 -0.717903
+ 2.985e+11Hz -0.659929 -0.717374
+ 2.986e+11Hz -0.660481 -0.716845
+ 2.987e+11Hz -0.661031 -0.716316
+ 2.988e+11Hz -0.661582 -0.715786
+ 2.989e+11Hz -0.662131 -0.715256
+ 2.99e+11Hz -0.662681 -0.714725
+ 2.991e+11Hz -0.66323 -0.714194
+ 2.992e+11Hz -0.663778 -0.713663
+ 2.993e+11Hz -0.664326 -0.713132
+ 2.994e+11Hz -0.664873 -0.7126
+ 2.995e+11Hz -0.66542 -0.712068
+ 2.996e+11Hz -0.665967 -0.711535
+ 2.997e+11Hz -0.666513 -0.711002
+ 2.998e+11Hz -0.667058 -0.710469
+ 2.999e+11Hz -0.667603 -0.709936
+ 3e+11Hz -0.668148 -0.709402
+ ]

A22 %vd(20 3) %vd(22, 3) xfer4
.model xfer4 xfer R_I=true table=[
+ 0Hz 0.0047718 0
+ 1e+08Hz 0.00477202 3.3416e-06
+ 2e+08Hz 0.00477265 6.6748e-06
+ 3e+08Hz 0.0047737 9.99121e-06
+ 4e+08Hz 0.00477517 1.32825e-05
+ 5e+08Hz 0.00477706 1.65402e-05
+ 6e+08Hz 0.00477937 1.9756e-05
+ 7e+08Hz 0.0047821 2.29215e-05
+ 8e+08Hz 0.00478524 2.60286e-05
+ 9e+08Hz 0.0047888 2.90688e-05
+ 1e+09Hz 0.00479277 3.20341e-05
+ 1.1e+09Hz 0.00479716 3.49161e-05
+ 1.2e+09Hz 0.00480195 3.77067e-05
+ 1.3e+09Hz 0.00480715 4.03978e-05
+ 1.4e+09Hz 0.00481276 4.29814e-05
+ 1.5e+09Hz 0.00481877 4.54495e-05
+ 1.6e+09Hz 0.00482518 4.77941e-05
+ 1.7e+09Hz 0.00483198 5.00074e-05
+ 1.8e+09Hz 0.00483919 5.20816e-05
+ 1.9e+09Hz 0.00484678 5.40089e-05
+ 2e+09Hz 0.00485476 5.57818e-05
+ 2.1e+09Hz 0.00486313 5.73926e-05
+ 2.2e+09Hz 0.00487188 5.88339e-05
+ 2.3e+09Hz 0.00488101 6.00983e-05
+ 2.4e+09Hz 0.00489051 6.11784e-05
+ 2.5e+09Hz 0.00490038 6.20672e-05
+ 2.6e+09Hz 0.00491061 6.27574e-05
+ 2.7e+09Hz 0.00492121 6.32421e-05
+ 2.8e+09Hz 0.00493216 6.35144e-05
+ 2.9e+09Hz 0.00494347 6.35675e-05
+ 3e+09Hz 0.00495512 6.33948e-05
+ 3.1e+09Hz 0.00496711 6.29896e-05
+ 3.2e+09Hz 0.00497945 6.23456e-05
+ 3.3e+09Hz 0.00499211 6.14564e-05
+ 3.4e+09Hz 0.0050051 6.03159e-05
+ 3.5e+09Hz 0.00501841 5.89179e-05
+ 3.6e+09Hz 0.00503204 5.72566e-05
+ 3.7e+09Hz 0.00504598 5.53262e-05
+ 3.8e+09Hz 0.00506022 5.3121e-05
+ 3.9e+09Hz 0.00507476 5.06354e-05
+ 4e+09Hz 0.00508959 4.78642e-05
+ 4.1e+09Hz 0.00510471 4.48019e-05
+ 4.2e+09Hz 0.00512011 4.14436e-05
+ 4.3e+09Hz 0.00513579 3.77843e-05
+ 4.4e+09Hz 0.00515173 3.38191e-05
+ 4.5e+09Hz 0.00516793 2.95435e-05
+ 4.6e+09Hz 0.00518439 2.49528e-05
+ 4.7e+09Hz 0.0052011 2.00428e-05
+ 4.8e+09Hz 0.00521804 1.48093e-05
+ 4.9e+09Hz 0.00523522 9.24808e-06
+ 5e+09Hz 0.00525263 3.3554e-06
+ 5.1e+09Hz 0.00527026 -2.87253e-06
+ 5.2e+09Hz 0.00528811 -9.43928e-06
+ 5.3e+09Hz 0.00530616 -1.63483e-05
+ 5.4e+09Hz 0.00532441 -2.36027e-05
+ 5.5e+09Hz 0.00534285 -3.12058e-05
+ 5.6e+09Hz 0.00536148 -3.91605e-05
+ 5.7e+09Hz 0.00538029 -4.74694e-05
+ 5.8e+09Hz 0.00539927 -5.61353e-05
+ 5.9e+09Hz 0.00541841 -6.51606e-05
+ 6e+09Hz 0.00543771 -7.45476e-05
+ 6.1e+09Hz 0.00545716 -8.42984e-05
+ 6.2e+09Hz 0.00547675 -9.44149e-05
+ 6.3e+09Hz 0.00549648 -0.000104899
+ 6.4e+09Hz 0.00551633 -0.000115753
+ 6.5e+09Hz 0.0055363 -0.000126977
+ 6.6e+09Hz 0.00555639 -0.000138573
+ 6.7e+09Hz 0.00557658 -0.000150542
+ 6.8e+09Hz 0.00559687 -0.000162886
+ 6.9e+09Hz 0.00561724 -0.000175605
+ 7e+09Hz 0.00563771 -0.0001887
+ 7.1e+09Hz 0.00565825 -0.00020217
+ 7.2e+09Hz 0.00567885 -0.000216018
+ 7.3e+09Hz 0.00569952 -0.000230243
+ 7.4e+09Hz 0.00572024 -0.000244844
+ 7.5e+09Hz 0.00574101 -0.000259822
+ 7.6e+09Hz 0.00576182 -0.000275178
+ 7.7e+09Hz 0.00578266 -0.000290909
+ 7.8e+09Hz 0.00580352 -0.000307016
+ 7.9e+09Hz 0.00582441 -0.000323498
+ 8e+09Hz 0.0058453 -0.000340355
+ 8.1e+09Hz 0.0058662 -0.000357584
+ 8.2e+09Hz 0.00588709 -0.000375186
+ 8.3e+09Hz 0.00590798 -0.000393159
+ 8.4e+09Hz 0.00592884 -0.000411502
+ 8.5e+09Hz 0.00594969 -0.000430212
+ 8.6e+09Hz 0.0059705 -0.000449289
+ 8.7e+09Hz 0.00599128 -0.00046873
+ 8.8e+09Hz 0.00601201 -0.000488534
+ 8.9e+09Hz 0.0060327 -0.000508699
+ 9e+09Hz 0.00605332 -0.000529222
+ 9.1e+09Hz 0.00607388 -0.000550101
+ 9.2e+09Hz 0.00609438 -0.000571334
+ 9.3e+09Hz 0.0061148 -0.000592918
+ 9.4e+09Hz 0.00613513 -0.00061485
+ 9.5e+09Hz 0.00615538 -0.000637128
+ 9.6e+09Hz 0.00617553 -0.000659749
+ 9.7e+09Hz 0.00619559 -0.00068271
+ 9.8e+09Hz 0.00621554 -0.000706007
+ 9.9e+09Hz 0.00623537 -0.000729638
+ 1e+10Hz 0.00625509 -0.0007536
+ 1.01e+10Hz 0.00627469 -0.000777888
+ 1.02e+10Hz 0.00629416 -0.000802499
+ 1.03e+10Hz 0.0063135 -0.00082743
+ 1.04e+10Hz 0.0063327 -0.000852677
+ 1.05e+10Hz 0.00635175 -0.000878236
+ 1.06e+10Hz 0.00637065 -0.000904103
+ 1.07e+10Hz 0.00638941 -0.000930275
+ 1.08e+10Hz 0.006408 -0.000956747
+ 1.09e+10Hz 0.00642643 -0.000983515
+ 1.1e+10Hz 0.00644469 -0.00101058
+ 1.11e+10Hz 0.00646278 -0.00103792
+ 1.12e+10Hz 0.00648069 -0.00106555
+ 1.13e+10Hz 0.00649842 -0.00109346
+ 1.14e+10Hz 0.00651597 -0.00112165
+ 1.15e+10Hz 0.00653332 -0.0011501
+ 1.16e+10Hz 0.00655049 -0.00117882
+ 1.17e+10Hz 0.00656745 -0.0012078
+ 1.18e+10Hz 0.00658422 -0.00123704
+ 1.19e+10Hz 0.00660078 -0.00126653
+ 1.2e+10Hz 0.00661713 -0.00129626
+ 1.21e+10Hz 0.00663328 -0.00132624
+ 1.22e+10Hz 0.0066492 -0.00135645
+ 1.23e+10Hz 0.00666491 -0.0013869
+ 1.24e+10Hz 0.0066804 -0.00141757
+ 1.25e+10Hz 0.00669567 -0.00144846
+ 1.26e+10Hz 0.00671071 -0.00147957
+ 1.27e+10Hz 0.00672552 -0.00151089
+ 1.28e+10Hz 0.0067401 -0.00154242
+ 1.29e+10Hz 0.00675444 -0.00157415
+ 1.3e+10Hz 0.00676855 -0.00160607
+ 1.31e+10Hz 0.00678242 -0.00163819
+ 1.32e+10Hz 0.00679605 -0.00167049
+ 1.33e+10Hz 0.00680944 -0.00170297
+ 1.34e+10Hz 0.00682259 -0.00173563
+ 1.35e+10Hz 0.00683548 -0.00176846
+ 1.36e+10Hz 0.00684813 -0.00180146
+ 1.37e+10Hz 0.00686054 -0.00183461
+ 1.38e+10Hz 0.00687269 -0.00186792
+ 1.39e+10Hz 0.00688459 -0.00190138
+ 1.4e+10Hz 0.00689623 -0.00193498
+ 1.41e+10Hz 0.00690763 -0.00196872
+ 1.42e+10Hz 0.00691877 -0.00200259
+ 1.43e+10Hz 0.00692965 -0.0020366
+ 1.44e+10Hz 0.00694028 -0.00207073
+ 1.45e+10Hz 0.00695065 -0.00210497
+ 1.46e+10Hz 0.00696076 -0.00213933
+ 1.47e+10Hz 0.00697062 -0.0021738
+ 1.48e+10Hz 0.00698022 -0.00220837
+ 1.49e+10Hz 0.00698956 -0.00224303
+ 1.5e+10Hz 0.00699865 -0.00227779
+ 1.51e+10Hz 0.00700747 -0.00231264
+ 1.52e+10Hz 0.00701604 -0.00234757
+ 1.53e+10Hz 0.00702435 -0.00238258
+ 1.54e+10Hz 0.00703241 -0.00241767
+ 1.55e+10Hz 0.00704021 -0.00245282
+ 1.56e+10Hz 0.00704775 -0.00248803
+ 1.57e+10Hz 0.00705504 -0.0025233
+ 1.58e+10Hz 0.00706207 -0.00255863
+ 1.59e+10Hz 0.00706885 -0.00259401
+ 1.6e+10Hz 0.00707538 -0.00262943
+ 1.61e+10Hz 0.00708166 -0.00266489
+ 1.62e+10Hz 0.00708769 -0.00270038
+ 1.63e+10Hz 0.00709347 -0.00273591
+ 1.64e+10Hz 0.007099 -0.00277146
+ 1.65e+10Hz 0.00710429 -0.00280704
+ 1.66e+10Hz 0.00710933 -0.00284263
+ 1.67e+10Hz 0.00711413 -0.00287824
+ 1.68e+10Hz 0.00711869 -0.00291386
+ 1.69e+10Hz 0.007123 -0.00294948
+ 1.7e+10Hz 0.00712709 -0.0029851
+ 1.71e+10Hz 0.00713093 -0.00302072
+ 1.72e+10Hz 0.00713454 -0.00305634
+ 1.73e+10Hz 0.00713792 -0.00309194
+ 1.74e+10Hz 0.00714107 -0.00312753
+ 1.75e+10Hz 0.007144 -0.0031631
+ 1.76e+10Hz 0.0071467 -0.00319865
+ 1.77e+10Hz 0.00714917 -0.00323418
+ 1.78e+10Hz 0.00715143 -0.00326967
+ 1.79e+10Hz 0.00715346 -0.00330514
+ 1.8e+10Hz 0.00715529 -0.00334057
+ 1.81e+10Hz 0.0071569 -0.00337596
+ 1.82e+10Hz 0.0071583 -0.00341131
+ 1.83e+10Hz 0.00715949 -0.00344661
+ 1.84e+10Hz 0.00716048 -0.00348187
+ 1.85e+10Hz 0.00716126 -0.00351707
+ 1.86e+10Hz 0.00716185 -0.00355222
+ 1.87e+10Hz 0.00716224 -0.00358732
+ 1.88e+10Hz 0.00716243 -0.00362236
+ 1.89e+10Hz 0.00716244 -0.00365733
+ 1.9e+10Hz 0.00716225 -0.00369224
+ 1.91e+10Hz 0.00716189 -0.00372709
+ 1.92e+10Hz 0.00716134 -0.00376186
+ 1.93e+10Hz 0.00716061 -0.00379657
+ 1.94e+10Hz 0.00715971 -0.0038312
+ 1.95e+10Hz 0.00715863 -0.00386576
+ 1.96e+10Hz 0.00715739 -0.00390024
+ 1.97e+10Hz 0.00715598 -0.00393464
+ 1.98e+10Hz 0.00715441 -0.00396895
+ 1.99e+10Hz 0.00715267 -0.00400319
+ 2e+10Hz 0.00715079 -0.00403734
+ 2.01e+10Hz 0.00714874 -0.00407141
+ 2.02e+10Hz 0.00714655 -0.00410539
+ 2.03e+10Hz 0.00714421 -0.00413928
+ 2.04e+10Hz 0.00714173 -0.00417308
+ 2.05e+10Hz 0.0071391 -0.00420679
+ 2.06e+10Hz 0.00713634 -0.0042404
+ 2.07e+10Hz 0.00713345 -0.00427393
+ 2.08e+10Hz 0.00713043 -0.00430736
+ 2.09e+10Hz 0.00712727 -0.00434069
+ 2.1e+10Hz 0.007124 -0.00437393
+ 2.11e+10Hz 0.0071206 -0.00440707
+ 2.12e+10Hz 0.00711709 -0.00444012
+ 2.13e+10Hz 0.00711346 -0.00447306
+ 2.14e+10Hz 0.00710972 -0.00450591
+ 2.15e+10Hz 0.00710587 -0.00453866
+ 2.16e+10Hz 0.00710192 -0.00457131
+ 2.17e+10Hz 0.00709786 -0.00460386
+ 2.18e+10Hz 0.00709371 -0.00463632
+ 2.19e+10Hz 0.00708946 -0.00466867
+ 2.2e+10Hz 0.00708512 -0.00470093
+ 2.21e+10Hz 0.00708069 -0.00473308
+ 2.22e+10Hz 0.00707617 -0.00476514
+ 2.23e+10Hz 0.00707157 -0.0047971
+ 2.24e+10Hz 0.00706689 -0.00482896
+ 2.25e+10Hz 0.00706213 -0.00486072
+ 2.26e+10Hz 0.0070573 -0.00489238
+ 2.27e+10Hz 0.00705239 -0.00492395
+ 2.28e+10Hz 0.00704742 -0.00495542
+ 2.29e+10Hz 0.00704238 -0.0049868
+ 2.3e+10Hz 0.00703728 -0.00501808
+ 2.31e+10Hz 0.00703211 -0.00504927
+ 2.32e+10Hz 0.00702689 -0.00508036
+ 2.33e+10Hz 0.00702161 -0.00511136
+ 2.34e+10Hz 0.00701628 -0.00514227
+ 2.35e+10Hz 0.0070109 -0.00517309
+ 2.36e+10Hz 0.00700547 -0.00520382
+ 2.37e+10Hz 0.00699999 -0.00523446
+ 2.38e+10Hz 0.00699447 -0.00526501
+ 2.39e+10Hz 0.00698891 -0.00529548
+ 2.4e+10Hz 0.00698331 -0.00532587
+ 2.41e+10Hz 0.00697767 -0.00535617
+ 2.42e+10Hz 0.006972 -0.00538639
+ 2.43e+10Hz 0.0069663 -0.00541653
+ 2.44e+10Hz 0.00696057 -0.00544659
+ 2.45e+10Hz 0.0069548 -0.00547657
+ 2.46e+10Hz 0.00694902 -0.00550648
+ 2.47e+10Hz 0.0069432 -0.00553631
+ 2.48e+10Hz 0.00693737 -0.00556607
+ 2.49e+10Hz 0.00693151 -0.00559576
+ 2.5e+10Hz 0.00692563 -0.00562538
+ 2.51e+10Hz 0.00691974 -0.00565493
+ 2.52e+10Hz 0.00691383 -0.00568442
+ 2.53e+10Hz 0.0069079 -0.00571384
+ 2.54e+10Hz 0.00690196 -0.0057432
+ 2.55e+10Hz 0.00689601 -0.0057725
+ 2.56e+10Hz 0.00689004 -0.00580175
+ 2.57e+10Hz 0.00688407 -0.00583093
+ 2.58e+10Hz 0.00687809 -0.00586006
+ 2.59e+10Hz 0.0068721 -0.00588914
+ 2.6e+10Hz 0.00686611 -0.00591816
+ 2.61e+10Hz 0.00686011 -0.00594714
+ 2.62e+10Hz 0.0068541 -0.00597607
+ 2.63e+10Hz 0.0068481 -0.00600495
+ 2.64e+10Hz 0.00684208 -0.00603379
+ 2.65e+10Hz 0.00683607 -0.00606259
+ 2.66e+10Hz 0.00683006 -0.00609135
+ 2.67e+10Hz 0.00682404 -0.00612007
+ 2.68e+10Hz 0.00681803 -0.00614876
+ 2.69e+10Hz 0.00681201 -0.00617741
+ 2.7e+10Hz 0.006806 -0.00620604
+ 2.71e+10Hz 0.00679998 -0.00623463
+ 2.72e+10Hz 0.00679397 -0.00626319
+ 2.73e+10Hz 0.00678796 -0.00629173
+ 2.74e+10Hz 0.00678195 -0.00632025
+ 2.75e+10Hz 0.00677594 -0.00634874
+ 2.76e+10Hz 0.00676994 -0.00637721
+ 2.77e+10Hz 0.00676394 -0.00640566
+ 2.78e+10Hz 0.00675793 -0.0064341
+ 2.79e+10Hz 0.00675193 -0.00646252
+ 2.8e+10Hz 0.00674593 -0.00649093
+ 2.81e+10Hz 0.00673994 -0.00651933
+ 2.82e+10Hz 0.00673394 -0.00654773
+ 2.83e+10Hz 0.00672795 -0.00657611
+ 2.84e+10Hz 0.00672195 -0.00660449
+ 2.85e+10Hz 0.00671596 -0.00663286
+ 2.86e+10Hz 0.00670996 -0.00666123
+ 2.87e+10Hz 0.00670396 -0.0066896
+ 2.88e+10Hz 0.00669797 -0.00671798
+ 2.89e+10Hz 0.00669197 -0.00674635
+ 2.9e+10Hz 0.00668596 -0.00677473
+ 2.91e+10Hz 0.00667996 -0.00680312
+ 2.92e+10Hz 0.00667394 -0.00683151
+ 2.93e+10Hz 0.00666793 -0.00685991
+ 2.94e+10Hz 0.00666191 -0.00688833
+ 2.95e+10Hz 0.00665588 -0.00691675
+ 2.96e+10Hz 0.00664984 -0.00694519
+ 2.97e+10Hz 0.00664379 -0.00697364
+ 2.98e+10Hz 0.00663774 -0.00700211
+ 2.99e+10Hz 0.00663167 -0.00703059
+ 3e+10Hz 0.00662559 -0.0070591
+ 3.01e+10Hz 0.0066195 -0.00708762
+ 3.02e+10Hz 0.0066134 -0.00711617
+ 3.03e+10Hz 0.00660728 -0.00714473
+ 3.04e+10Hz 0.00660115 -0.00717332
+ 3.05e+10Hz 0.00659499 -0.00720193
+ 3.06e+10Hz 0.00658882 -0.00723057
+ 3.07e+10Hz 0.00658263 -0.00725924
+ 3.08e+10Hz 0.00657642 -0.00728793
+ 3.09e+10Hz 0.00657018 -0.00731664
+ 3.1e+10Hz 0.00656392 -0.00734539
+ 3.11e+10Hz 0.00655764 -0.00737417
+ 3.12e+10Hz 0.00655133 -0.00740297
+ 3.13e+10Hz 0.00654499 -0.00743181
+ 3.14e+10Hz 0.00653862 -0.00746067
+ 3.15e+10Hz 0.00653223 -0.00748957
+ 3.16e+10Hz 0.0065258 -0.00751851
+ 3.17e+10Hz 0.00651933 -0.00754747
+ 3.18e+10Hz 0.00651284 -0.00757647
+ 3.19e+10Hz 0.0065063 -0.0076055
+ 3.2e+10Hz 0.00649973 -0.00763456
+ 3.21e+10Hz 0.00649312 -0.00766366
+ 3.22e+10Hz 0.00648647 -0.0076928
+ 3.23e+10Hz 0.00647977 -0.00772197
+ 3.24e+10Hz 0.00647304 -0.00775117
+ 3.25e+10Hz 0.00646626 -0.00778041
+ 3.26e+10Hz 0.00645943 -0.00780968
+ 3.27e+10Hz 0.00645255 -0.00783899
+ 3.28e+10Hz 0.00644563 -0.00786834
+ 3.29e+10Hz 0.00643865 -0.00789772
+ 3.3e+10Hz 0.00643162 -0.00792713
+ 3.31e+10Hz 0.00642454 -0.00795658
+ 3.32e+10Hz 0.00641741 -0.00798607
+ 3.33e+10Hz 0.00641021 -0.00801559
+ 3.34e+10Hz 0.00640296 -0.00804514
+ 3.35e+10Hz 0.00639565 -0.00807473
+ 3.36e+10Hz 0.00638828 -0.00810435
+ 3.37e+10Hz 0.00638085 -0.00813401
+ 3.38e+10Hz 0.00637336 -0.0081637
+ 3.39e+10Hz 0.00636579 -0.00819342
+ 3.4e+10Hz 0.00635817 -0.00822317
+ 3.41e+10Hz 0.00635047 -0.00825296
+ 3.42e+10Hz 0.00634271 -0.00828277
+ 3.43e+10Hz 0.00633488 -0.00831262
+ 3.44e+10Hz 0.00632698 -0.00834249
+ 3.45e+10Hz 0.006319 -0.00837239
+ 3.46e+10Hz 0.00631095 -0.00840233
+ 3.47e+10Hz 0.00630283 -0.00843229
+ 3.48e+10Hz 0.00629463 -0.00846227
+ 3.49e+10Hz 0.00628635 -0.00849228
+ 3.5e+10Hz 0.006278 -0.00852232
+ 3.51e+10Hz 0.00626956 -0.00855238
+ 3.52e+10Hz 0.00626105 -0.00858247
+ 3.53e+10Hz 0.00625245 -0.00861258
+ 3.54e+10Hz 0.00624377 -0.0086427
+ 3.55e+10Hz 0.00623501 -0.00867285
+ 3.56e+10Hz 0.00622617 -0.00870302
+ 3.57e+10Hz 0.00621724 -0.00873321
+ 3.58e+10Hz 0.00620822 -0.00876341
+ 3.59e+10Hz 0.00619912 -0.00879363
+ 3.6e+10Hz 0.00618992 -0.00882387
+ 3.61e+10Hz 0.00618064 -0.00885412
+ 3.62e+10Hz 0.00617128 -0.00888438
+ 3.63e+10Hz 0.00616182 -0.00891465
+ 3.64e+10Hz 0.00615227 -0.00894494
+ 3.65e+10Hz 0.00614262 -0.00897523
+ 3.66e+10Hz 0.00613289 -0.00900553
+ 3.67e+10Hz 0.00612307 -0.00903584
+ 3.68e+10Hz 0.00611315 -0.00906616
+ 3.69e+10Hz 0.00610313 -0.00909648
+ 3.7e+10Hz 0.00609303 -0.0091268
+ 3.71e+10Hz 0.00608282 -0.00915712
+ 3.72e+10Hz 0.00607253 -0.00918745
+ 3.73e+10Hz 0.00606213 -0.00921777
+ 3.74e+10Hz 0.00605165 -0.00924809
+ 3.75e+10Hz 0.00604106 -0.00927841
+ 3.76e+10Hz 0.00603038 -0.00930872
+ 3.77e+10Hz 0.0060196 -0.00933903
+ 3.78e+10Hz 0.00600873 -0.00936933
+ 3.79e+10Hz 0.00599776 -0.00939962
+ 3.8e+10Hz 0.00598669 -0.0094299
+ 3.81e+10Hz 0.00597552 -0.00946017
+ 3.82e+10Hz 0.00596426 -0.00949043
+ 3.83e+10Hz 0.0059529 -0.00952067
+ 3.84e+10Hz 0.00594144 -0.0095509
+ 3.85e+10Hz 0.00592989 -0.00958111
+ 3.86e+10Hz 0.00591823 -0.00961131
+ 3.87e+10Hz 0.00590648 -0.00964148
+ 3.88e+10Hz 0.00589464 -0.00967163
+ 3.89e+10Hz 0.00588269 -0.00970177
+ 3.9e+10Hz 0.00587065 -0.00973187
+ 3.91e+10Hz 0.00585851 -0.00976196
+ 3.92e+10Hz 0.00584628 -0.00979201
+ 3.93e+10Hz 0.00583395 -0.00982204
+ 3.94e+10Hz 0.00582152 -0.00985205
+ 3.95e+10Hz 0.005809 -0.00988202
+ 3.96e+10Hz 0.00579639 -0.00991196
+ 3.97e+10Hz 0.00578368 -0.00994187
+ 3.98e+10Hz 0.00577088 -0.00997175
+ 3.99e+10Hz 0.00575798 -0.0100016
+ 4e+10Hz 0.00574499 -0.0100314
+ 4.01e+10Hz 0.00573191 -0.0100612
+ 4.02e+10Hz 0.00571873 -0.0100909
+ 4.03e+10Hz 0.00570547 -0.0101206
+ 4.04e+10Hz 0.00569211 -0.0101502
+ 4.05e+10Hz 0.00567866 -0.0101798
+ 4.06e+10Hz 0.00566513 -0.0102094
+ 4.07e+10Hz 0.0056515 -0.0102389
+ 4.08e+10Hz 0.00563779 -0.0102684
+ 4.09e+10Hz 0.00562399 -0.0102979
+ 4.1e+10Hz 0.00561011 -0.0103272
+ 4.11e+10Hz 0.00559614 -0.0103566
+ 4.12e+10Hz 0.00558208 -0.0103859
+ 4.13e+10Hz 0.00556794 -0.0104151
+ 4.14e+10Hz 0.00555372 -0.0104443
+ 4.15e+10Hz 0.00553941 -0.0104734
+ 4.16e+10Hz 0.00552503 -0.0105025
+ 4.17e+10Hz 0.00551056 -0.0105316
+ 4.18e+10Hz 0.00549601 -0.0105605
+ 4.19e+10Hz 0.00548139 -0.0105895
+ 4.2e+10Hz 0.00546669 -0.0106183
+ 4.21e+10Hz 0.00545191 -0.0106472
+ 4.22e+10Hz 0.00543705 -0.0106759
+ 4.23e+10Hz 0.00542212 -0.0107046
+ 4.24e+10Hz 0.00540712 -0.0107333
+ 4.25e+10Hz 0.00539205 -0.0107619
+ 4.26e+10Hz 0.0053769 -0.0107904
+ 4.27e+10Hz 0.00536168 -0.0108189
+ 4.28e+10Hz 0.0053464 -0.0108473
+ 4.29e+10Hz 0.00533104 -0.0108756
+ 4.3e+10Hz 0.00531562 -0.0109039
+ 4.31e+10Hz 0.00530013 -0.0109321
+ 4.32e+10Hz 0.00528458 -0.0109603
+ 4.33e+10Hz 0.00526896 -0.0109884
+ 4.34e+10Hz 0.00525328 -0.0110164
+ 4.35e+10Hz 0.00523754 -0.0110444
+ 4.36e+10Hz 0.00522174 -0.0110723
+ 4.37e+10Hz 0.00520587 -0.0111001
+ 4.38e+10Hz 0.00518995 -0.0111279
+ 4.39e+10Hz 0.00517397 -0.0111556
+ 4.4e+10Hz 0.00515794 -0.0111833
+ 4.41e+10Hz 0.00514185 -0.0112109
+ 4.42e+10Hz 0.0051257 -0.0112384
+ 4.43e+10Hz 0.00510951 -0.0112659
+ 4.44e+10Hz 0.00509326 -0.0112933
+ 4.45e+10Hz 0.00507696 -0.0113206
+ 4.46e+10Hz 0.00506061 -0.0113479
+ 4.47e+10Hz 0.00504421 -0.0113751
+ 4.48e+10Hz 0.00502776 -0.0114022
+ 4.49e+10Hz 0.00501127 -0.0114293
+ 4.5e+10Hz 0.00499473 -0.0114563
+ 4.51e+10Hz 0.00497815 -0.0114833
+ 4.52e+10Hz 0.00496152 -0.0115102
+ 4.53e+10Hz 0.00494485 -0.011537
+ 4.54e+10Hz 0.00492814 -0.0115637
+ 4.55e+10Hz 0.00491139 -0.0115904
+ 4.56e+10Hz 0.0048946 -0.0116171
+ 4.57e+10Hz 0.00487777 -0.0116436
+ 4.58e+10Hz 0.00486091 -0.0116701
+ 4.59e+10Hz 0.004844 -0.0116966
+ 4.6e+10Hz 0.00482706 -0.0117229
+ 4.61e+10Hz 0.00481009 -0.0117493
+ 4.62e+10Hz 0.00479308 -0.0117755
+ 4.63e+10Hz 0.00477604 -0.0118017
+ 4.64e+10Hz 0.00475897 -0.0118279
+ 4.65e+10Hz 0.00474187 -0.0118539
+ 4.66e+10Hz 0.00472473 -0.01188
+ 4.67e+10Hz 0.00470757 -0.0119059
+ 4.68e+10Hz 0.00469037 -0.0119318
+ 4.69e+10Hz 0.00467315 -0.0119577
+ 4.7e+10Hz 0.0046559 -0.0119834
+ 4.71e+10Hz 0.00463863 -0.0120092
+ 4.72e+10Hz 0.00462133 -0.0120349
+ 4.73e+10Hz 0.004604 -0.0120605
+ 4.74e+10Hz 0.00458665 -0.012086
+ 4.75e+10Hz 0.00456928 -0.0121115
+ 4.76e+10Hz 0.00455188 -0.012137
+ 4.77e+10Hz 0.00453446 -0.0121624
+ 4.78e+10Hz 0.00451701 -0.0121878
+ 4.79e+10Hz 0.00449955 -0.0122131
+ 4.8e+10Hz 0.00448206 -0.0122383
+ 4.81e+10Hz 0.00446456 -0.0122635
+ 4.82e+10Hz 0.00444703 -0.0122887
+ 4.83e+10Hz 0.00442948 -0.0123138
+ 4.84e+10Hz 0.00441192 -0.0123388
+ 4.85e+10Hz 0.00439433 -0.0123638
+ 4.86e+10Hz 0.00437673 -0.0123888
+ 4.87e+10Hz 0.00435911 -0.0124137
+ 4.88e+10Hz 0.00434147 -0.0124386
+ 4.89e+10Hz 0.00432381 -0.0124634
+ 4.9e+10Hz 0.00430614 -0.0124882
+ 4.91e+10Hz 0.00428845 -0.0125129
+ 4.92e+10Hz 0.00427074 -0.0125376
+ 4.93e+10Hz 0.00425302 -0.0125623
+ 4.94e+10Hz 0.00423528 -0.0125869
+ 4.95e+10Hz 0.00421752 -0.0126114
+ 4.96e+10Hz 0.00419975 -0.012636
+ 4.97e+10Hz 0.00418197 -0.0126605
+ 4.98e+10Hz 0.00416416 -0.0126849
+ 4.99e+10Hz 0.00414634 -0.0127094
+ 5e+10Hz 0.00412851 -0.0127337
+ 5.01e+10Hz 0.00411066 -0.0127581
+ 5.02e+10Hz 0.00409279 -0.0127824
+ 5.03e+10Hz 0.00407491 -0.0128067
+ 5.04e+10Hz 0.00405702 -0.0128309
+ 5.05e+10Hz 0.00403911 -0.0128552
+ 5.06e+10Hz 0.00402118 -0.0128793
+ 5.07e+10Hz 0.00400323 -0.0129035
+ 5.08e+10Hz 0.00398527 -0.0129276
+ 5.09e+10Hz 0.0039673 -0.0129517
+ 5.1e+10Hz 0.0039493 -0.0129758
+ 5.11e+10Hz 0.00393129 -0.0129998
+ 5.12e+10Hz 0.00391327 -0.0130238
+ 5.13e+10Hz 0.00389523 -0.0130478
+ 5.14e+10Hz 0.00387717 -0.0130718
+ 5.15e+10Hz 0.00385909 -0.0130957
+ 5.16e+10Hz 0.00384099 -0.0131196
+ 5.17e+10Hz 0.00382288 -0.0131435
+ 5.18e+10Hz 0.00380475 -0.0131673
+ 5.19e+10Hz 0.00378659 -0.0131912
+ 5.2e+10Hz 0.00376842 -0.013215
+ 5.21e+10Hz 0.00375023 -0.0132388
+ 5.22e+10Hz 0.00373202 -0.0132625
+ 5.23e+10Hz 0.00371379 -0.0132863
+ 5.24e+10Hz 0.00369554 -0.01331
+ 5.25e+10Hz 0.00367727 -0.0133337
+ 5.26e+10Hz 0.00365898 -0.0133574
+ 5.27e+10Hz 0.00364066 -0.013381
+ 5.28e+10Hz 0.00362232 -0.0134047
+ 5.29e+10Hz 0.00360396 -0.0134283
+ 5.3e+10Hz 0.00358558 -0.0134519
+ 5.31e+10Hz 0.00356717 -0.0134755
+ 5.32e+10Hz 0.00354873 -0.0134991
+ 5.33e+10Hz 0.00353027 -0.0135226
+ 5.34e+10Hz 0.00351179 -0.0135462
+ 5.35e+10Hz 0.00349328 -0.0135697
+ 5.36e+10Hz 0.00347474 -0.0135932
+ 5.37e+10Hz 0.00345617 -0.0136167
+ 5.38e+10Hz 0.00343758 -0.0136402
+ 5.39e+10Hz 0.00341896 -0.0136636
+ 5.4e+10Hz 0.00340031 -0.0136871
+ 5.41e+10Hz 0.00338162 -0.0137105
+ 5.42e+10Hz 0.00336291 -0.0137339
+ 5.43e+10Hz 0.00334417 -0.0137573
+ 5.44e+10Hz 0.0033254 -0.0137807
+ 5.45e+10Hz 0.00330659 -0.0138041
+ 5.46e+10Hz 0.00328775 -0.0138274
+ 5.47e+10Hz 0.00326888 -0.0138507
+ 5.48e+10Hz 0.00324997 -0.0138741
+ 5.49e+10Hz 0.00323103 -0.0138974
+ 5.5e+10Hz 0.00321206 -0.0139207
+ 5.51e+10Hz 0.00319305 -0.013944
+ 5.52e+10Hz 0.003174 -0.0139672
+ 5.53e+10Hz 0.00315491 -0.0139905
+ 5.54e+10Hz 0.00313579 -0.0140137
+ 5.55e+10Hz 0.00311663 -0.0140369
+ 5.56e+10Hz 0.00309743 -0.0140601
+ 5.57e+10Hz 0.00307819 -0.0140833
+ 5.58e+10Hz 0.00305891 -0.0141065
+ 5.59e+10Hz 0.00303959 -0.0141296
+ 5.6e+10Hz 0.00302023 -0.0141528
+ 5.61e+10Hz 0.00300083 -0.0141759
+ 5.62e+10Hz 0.00298138 -0.014199
+ 5.63e+10Hz 0.0029619 -0.0142221
+ 5.64e+10Hz 0.00294236 -0.0142452
+ 5.65e+10Hz 0.00292279 -0.0142682
+ 5.66e+10Hz 0.00290317 -0.0142913
+ 5.67e+10Hz 0.0028835 -0.0143143
+ 5.68e+10Hz 0.00286379 -0.0143373
+ 5.69e+10Hz 0.00284404 -0.0143603
+ 5.7e+10Hz 0.00282424 -0.0143832
+ 5.71e+10Hz 0.00280439 -0.0144062
+ 5.72e+10Hz 0.00278449 -0.0144291
+ 5.73e+10Hz 0.00276454 -0.014452
+ 5.74e+10Hz 0.00274455 -0.0144749
+ 5.75e+10Hz 0.00272451 -0.0144978
+ 5.76e+10Hz 0.00270442 -0.0145206
+ 5.77e+10Hz 0.00268427 -0.0145434
+ 5.78e+10Hz 0.00266408 -0.0145662
+ 5.79e+10Hz 0.00264384 -0.014589
+ 5.8e+10Hz 0.00262355 -0.0146117
+ 5.81e+10Hz 0.0026032 -0.0146345
+ 5.82e+10Hz 0.00258281 -0.0146571
+ 5.83e+10Hz 0.00256236 -0.0146798
+ 5.84e+10Hz 0.00254186 -0.0147025
+ 5.85e+10Hz 0.00252131 -0.0147251
+ 5.86e+10Hz 0.00250071 -0.0147477
+ 5.87e+10Hz 0.00248005 -0.0147702
+ 5.88e+10Hz 0.00245934 -0.0147928
+ 5.89e+10Hz 0.00243858 -0.0148153
+ 5.9e+10Hz 0.00241776 -0.0148378
+ 5.91e+10Hz 0.00239689 -0.0148602
+ 5.92e+10Hz 0.00237597 -0.0148826
+ 5.93e+10Hz 0.00235499 -0.014905
+ 5.94e+10Hz 0.00233395 -0.0149274
+ 5.95e+10Hz 0.00231287 -0.0149497
+ 5.96e+10Hz 0.00229172 -0.014972
+ 5.97e+10Hz 0.00227053 -0.0149942
+ 5.98e+10Hz 0.00224928 -0.0150164
+ 5.99e+10Hz 0.00222797 -0.0150386
+ 6e+10Hz 0.00220661 -0.0150607
+ 6.01e+10Hz 0.0021852 -0.0150829
+ 6.02e+10Hz 0.00216373 -0.0151049
+ 6.03e+10Hz 0.0021422 -0.015127
+ 6.04e+10Hz 0.00212063 -0.0151489
+ 6.05e+10Hz 0.00209899 -0.0151709
+ 6.06e+10Hz 0.00207731 -0.0151928
+ 6.07e+10Hz 0.00205556 -0.0152147
+ 6.08e+10Hz 0.00203377 -0.0152365
+ 6.09e+10Hz 0.00201192 -0.0152583
+ 6.1e+10Hz 0.00199002 -0.01528
+ 6.11e+10Hz 0.00196806 -0.0153017
+ 6.12e+10Hz 0.00194605 -0.0153234
+ 6.13e+10Hz 0.00192398 -0.015345
+ 6.14e+10Hz 0.00190187 -0.0153665
+ 6.15e+10Hz 0.0018797 -0.015388
+ 6.16e+10Hz 0.00185747 -0.0154095
+ 6.17e+10Hz 0.0018352 -0.0154309
+ 6.18e+10Hz 0.00181287 -0.0154523
+ 6.19e+10Hz 0.00179049 -0.0154736
+ 6.2e+10Hz 0.00176806 -0.0154949
+ 6.21e+10Hz 0.00174558 -0.0155161
+ 6.22e+10Hz 0.00172305 -0.0155373
+ 6.23e+10Hz 0.00170047 -0.0155584
+ 6.24e+10Hz 0.00167783 -0.0155795
+ 6.25e+10Hz 0.00165515 -0.0156005
+ 6.26e+10Hz 0.00163242 -0.0156214
+ 6.27e+10Hz 0.00160964 -0.0156423
+ 6.28e+10Hz 0.00158682 -0.0156632
+ 6.29e+10Hz 0.00156394 -0.015684
+ 6.3e+10Hz 0.00154102 -0.0157047
+ 6.31e+10Hz 0.00151805 -0.0157254
+ 6.32e+10Hz 0.00149503 -0.015746
+ 6.33e+10Hz 0.00147197 -0.0157666
+ 6.34e+10Hz 0.00144886 -0.0157871
+ 6.35e+10Hz 0.00142571 -0.0158076
+ 6.36e+10Hz 0.00140252 -0.015828
+ 6.37e+10Hz 0.00137928 -0.0158483
+ 6.38e+10Hz 0.001356 -0.0158686
+ 6.39e+10Hz 0.00133267 -0.0158888
+ 6.4e+10Hz 0.0013093 -0.015909
+ 6.41e+10Hz 0.0012859 -0.0159291
+ 6.42e+10Hz 0.00126245 -0.0159491
+ 6.43e+10Hz 0.00123896 -0.0159691
+ 6.44e+10Hz 0.00121543 -0.015989
+ 6.45e+10Hz 0.00119186 -0.0160089
+ 6.46e+10Hz 0.00116826 -0.0160287
+ 6.47e+10Hz 0.00114461 -0.0160484
+ 6.48e+10Hz 0.00112093 -0.016068
+ 6.49e+10Hz 0.00109722 -0.0160876
+ 6.5e+10Hz 0.00107346 -0.0161072
+ 6.51e+10Hz 0.00104968 -0.0161267
+ 6.52e+10Hz 0.00102586 -0.0161461
+ 6.53e+10Hz 0.001002 -0.0161654
+ 6.54e+10Hz 0.000978114 -0.0161847
+ 6.55e+10Hz 0.000954194 -0.0162039
+ 6.56e+10Hz 0.000930242 -0.0162231
+ 6.57e+10Hz 0.000906259 -0.0162422
+ 6.58e+10Hz 0.000882246 -0.0162612
+ 6.59e+10Hz 0.000858204 -0.0162802
+ 6.6e+10Hz 0.000834133 -0.0162991
+ 6.61e+10Hz 0.000810033 -0.0163179
+ 6.62e+10Hz 0.000785906 -0.0163367
+ 6.63e+10Hz 0.000761752 -0.0163554
+ 6.64e+10Hz 0.000737572 -0.016374
+ 6.65e+10Hz 0.000713366 -0.0163926
+ 6.66e+10Hz 0.000689136 -0.0164111
+ 6.67e+10Hz 0.000664881 -0.0164295
+ 6.68e+10Hz 0.000640603 -0.0164479
+ 6.69e+10Hz 0.000616302 -0.0164662
+ 6.7e+10Hz 0.000591979 -0.0164845
+ 6.71e+10Hz 0.000567634 -0.0165026
+ 6.72e+10Hz 0.000543269 -0.0165208
+ 6.73e+10Hz 0.000518883 -0.0165388
+ 6.74e+10Hz 0.000494478 -0.0165568
+ 6.75e+10Hz 0.000470054 -0.0165747
+ 6.76e+10Hz 0.000445611 -0.0165926
+ 6.77e+10Hz 0.000421151 -0.0166104
+ 6.78e+10Hz 0.000396674 -0.0166281
+ 6.79e+10Hz 0.00037218 -0.0166458
+ 6.8e+10Hz 0.00034767 -0.0166634
+ 6.81e+10Hz 0.000323145 -0.016681
+ 6.82e+10Hz 0.000298606 -0.0166985
+ 6.83e+10Hz 0.000274052 -0.0167159
+ 6.84e+10Hz 0.000249484 -0.0167332
+ 6.85e+10Hz 0.000224904 -0.0167505
+ 6.86e+10Hz 0.00020031 -0.0167678
+ 6.87e+10Hz 0.000175705 -0.016785
+ 6.88e+10Hz 0.000151089 -0.0168021
+ 6.89e+10Hz 0.000126461 -0.0168191
+ 6.9e+10Hz 0.000101823 -0.0168361
+ 6.91e+10Hz 7.71752e-05 -0.0168531
+ 6.92e+10Hz 5.25176e-05 -0.01687
+ 6.93e+10Hz 2.7851e-05 -0.0168868
+ 6.94e+10Hz 3.17567e-06 -0.0169035
+ 6.95e+10Hz -2.15078e-05 -0.0169202
+ 6.96e+10Hz -4.61991e-05 -0.0169369
+ 6.97e+10Hz -7.08978e-05 -0.0169535
+ 6.98e+10Hz -9.56035e-05 -0.01697
+ 6.99e+10Hz -0.000120316 -0.0169865
+ 7e+10Hz -0.000145034 -0.0170029
+ 7.01e+10Hz -0.000169759 -0.0170193
+ 7.02e+10Hz -0.000194489 -0.0170356
+ 7.03e+10Hz -0.000219224 -0.0170519
+ 7.04e+10Hz -0.000243964 -0.0170681
+ 7.05e+10Hz -0.000268709 -0.0170842
+ 7.06e+10Hz -0.000293458 -0.0171003
+ 7.07e+10Hz -0.000318212 -0.0171163
+ 7.08e+10Hz -0.000342969 -0.0171323
+ 7.09e+10Hz -0.00036773 -0.0171483
+ 7.1e+10Hz -0.000392494 -0.0171642
+ 7.11e+10Hz -0.000417262 -0.01718
+ 7.12e+10Hz -0.000442032 -0.0171958
+ 7.13e+10Hz -0.000466806 -0.0172116
+ 7.14e+10Hz -0.000491582 -0.0172272
+ 7.15e+10Hz -0.000516361 -0.0172429
+ 7.16e+10Hz -0.000541142 -0.0172585
+ 7.17e+10Hz -0.000565925 -0.017274
+ 7.18e+10Hz -0.000590711 -0.0172895
+ 7.19e+10Hz -0.000615499 -0.017305
+ 7.2e+10Hz -0.000640289 -0.0173204
+ 7.21e+10Hz -0.000665081 -0.0173358
+ 7.22e+10Hz -0.000689875 -0.0173511
+ 7.23e+10Hz -0.000714671 -0.0173664
+ 7.24e+10Hz -0.000739469 -0.0173816
+ 7.25e+10Hz -0.000764269 -0.0173968
+ 7.26e+10Hz -0.000789071 -0.0174119
+ 7.27e+10Hz -0.000813875 -0.017427
+ 7.28e+10Hz -0.000838681 -0.0174421
+ 7.29e+10Hz -0.00086349 -0.0174571
+ 7.3e+10Hz -0.0008883 -0.0174721
+ 7.31e+10Hz -0.000913113 -0.017487
+ 7.32e+10Hz -0.000937929 -0.0175019
+ 7.33e+10Hz -0.000962747 -0.0175168
+ 7.34e+10Hz -0.000987567 -0.0175316
+ 7.35e+10Hz -0.00101239 -0.0175464
+ 7.36e+10Hz -0.00103722 -0.0175611
+ 7.37e+10Hz -0.00106205 -0.0175758
+ 7.38e+10Hz -0.00108688 -0.0175905
+ 7.39e+10Hz -0.00111172 -0.0176051
+ 7.4e+10Hz -0.00113656 -0.0176197
+ 7.41e+10Hz -0.0011614 -0.0176343
+ 7.42e+10Hz -0.00118625 -0.0176488
+ 7.43e+10Hz -0.0012111 -0.0176633
+ 7.44e+10Hz -0.00123596 -0.0176778
+ 7.45e+10Hz -0.00126082 -0.0176922
+ 7.46e+10Hz -0.00128569 -0.0177066
+ 7.47e+10Hz -0.00131056 -0.0177209
+ 7.48e+10Hz -0.00133544 -0.0177352
+ 7.49e+10Hz -0.00136033 -0.0177495
+ 7.5e+10Hz -0.00138522 -0.0177638
+ 7.51e+10Hz -0.00141012 -0.017778
+ 7.52e+10Hz -0.00143503 -0.0177921
+ 7.53e+10Hz -0.00145994 -0.0178063
+ 7.54e+10Hz -0.00148486 -0.0178204
+ 7.55e+10Hz -0.00150979 -0.0178345
+ 7.56e+10Hz -0.00153472 -0.0178486
+ 7.57e+10Hz -0.00155967 -0.0178626
+ 7.58e+10Hz -0.00158463 -0.0178766
+ 7.59e+10Hz -0.00160959 -0.0178905
+ 7.6e+10Hz -0.00163456 -0.0179045
+ 7.61e+10Hz -0.00165955 -0.0179184
+ 7.62e+10Hz -0.00168454 -0.0179322
+ 7.63e+10Hz -0.00170955 -0.0179461
+ 7.64e+10Hz -0.00173457 -0.0179599
+ 7.65e+10Hz -0.0017596 -0.0179737
+ 7.66e+10Hz -0.00178464 -0.0179874
+ 7.67e+10Hz -0.00180969 -0.0180011
+ 7.68e+10Hz -0.00183476 -0.0180148
+ 7.69e+10Hz -0.00185984 -0.0180285
+ 7.7e+10Hz -0.00188493 -0.0180421
+ 7.71e+10Hz -0.00191004 -0.0180557
+ 7.72e+10Hz -0.00193516 -0.0180693
+ 7.73e+10Hz -0.0019603 -0.0180828
+ 7.74e+10Hz -0.00198546 -0.0180963
+ 7.75e+10Hz -0.00201062 -0.0181098
+ 7.76e+10Hz -0.00203581 -0.0181232
+ 7.77e+10Hz -0.00206101 -0.0181366
+ 7.78e+10Hz -0.00208623 -0.01815
+ 7.79e+10Hz -0.00211147 -0.0181634
+ 7.8e+10Hz -0.00213672 -0.0181767
+ 7.81e+10Hz -0.00216199 -0.01819
+ 7.82e+10Hz -0.00218728 -0.0182033
+ 7.83e+10Hz -0.00221259 -0.0182165
+ 7.84e+10Hz -0.00223792 -0.0182297
+ 7.85e+10Hz -0.00226327 -0.0182429
+ 7.86e+10Hz -0.00228864 -0.018256
+ 7.87e+10Hz -0.00231403 -0.0182691
+ 7.88e+10Hz -0.00233944 -0.0182822
+ 7.89e+10Hz -0.00236487 -0.0182952
+ 7.9e+10Hz -0.00239032 -0.0183083
+ 7.91e+10Hz -0.0024158 -0.0183212
+ 7.92e+10Hz -0.00244129 -0.0183342
+ 7.93e+10Hz -0.00246681 -0.0183471
+ 7.94e+10Hz -0.00249235 -0.01836
+ 7.95e+10Hz -0.00251792 -0.0183728
+ 7.96e+10Hz -0.00254351 -0.0183856
+ 7.97e+10Hz -0.00256912 -0.0183984
+ 7.98e+10Hz -0.00259475 -0.0184112
+ 7.99e+10Hz -0.00262041 -0.0184239
+ 8e+10Hz -0.0026461 -0.0184366
+ 8.01e+10Hz -0.00267181 -0.0184492
+ 8.02e+10Hz -0.00269754 -0.0184618
+ 8.03e+10Hz -0.0027233 -0.0184744
+ 8.04e+10Hz -0.00274908 -0.0184869
+ 8.05e+10Hz -0.00277489 -0.0184994
+ 8.06e+10Hz -0.00280073 -0.0185119
+ 8.07e+10Hz -0.00282659 -0.0185243
+ 8.08e+10Hz -0.00285248 -0.0185367
+ 8.09e+10Hz -0.0028784 -0.018549
+ 8.1e+10Hz -0.00290434 -0.0185613
+ 8.11e+10Hz -0.00293031 -0.0185736
+ 8.12e+10Hz -0.0029563 -0.0185858
+ 8.13e+10Hz -0.00298233 -0.018598
+ 8.14e+10Hz -0.00300838 -0.0186101
+ 8.15e+10Hz -0.00303445 -0.0186222
+ 8.16e+10Hz -0.00306056 -0.0186343
+ 8.17e+10Hz -0.00308669 -0.0186463
+ 8.18e+10Hz -0.00311285 -0.0186583
+ 8.19e+10Hz -0.00313904 -0.0186702
+ 8.2e+10Hz -0.00316525 -0.0186821
+ 8.21e+10Hz -0.00319149 -0.018694
+ 8.22e+10Hz -0.00321776 -0.0187058
+ 8.23e+10Hz -0.00324406 -0.0187175
+ 8.24e+10Hz -0.00327039 -0.0187293
+ 8.25e+10Hz -0.00329674 -0.0187409
+ 8.26e+10Hz -0.00332312 -0.0187525
+ 8.27e+10Hz -0.00334953 -0.0187641
+ 8.28e+10Hz -0.00337596 -0.0187756
+ 8.29e+10Hz -0.00340242 -0.0187871
+ 8.3e+10Hz -0.00342892 -0.0187986
+ 8.31e+10Hz -0.00345543 -0.0188099
+ 8.32e+10Hz -0.00348198 -0.0188213
+ 8.33e+10Hz -0.00350855 -0.0188326
+ 8.34e+10Hz -0.00353515 -0.0188438
+ 8.35e+10Hz -0.00356177 -0.018855
+ 8.36e+10Hz -0.00358843 -0.0188661
+ 8.37e+10Hz -0.0036151 -0.0188772
+ 8.38e+10Hz -0.00364181 -0.0188882
+ 8.39e+10Hz -0.00366854 -0.0188992
+ 8.4e+10Hz -0.0036953 -0.0189101
+ 8.41e+10Hz -0.00372208 -0.018921
+ 8.42e+10Hz -0.00374888 -0.0189318
+ 8.43e+10Hz -0.00377572 -0.0189426
+ 8.44e+10Hz -0.00380258 -0.0189533
+ 8.45e+10Hz -0.00382946 -0.0189639
+ 8.46e+10Hz -0.00385636 -0.0189745
+ 8.47e+10Hz -0.00388329 -0.0189851
+ 8.48e+10Hz -0.00391025 -0.0189956
+ 8.49e+10Hz -0.00393723 -0.019006
+ 8.5e+10Hz -0.00396423 -0.0190164
+ 8.51e+10Hz -0.00399125 -0.0190267
+ 8.52e+10Hz -0.0040183 -0.0190369
+ 8.53e+10Hz -0.00404537 -0.0190471
+ 8.54e+10Hz -0.00407246 -0.0190573
+ 8.55e+10Hz -0.00409957 -0.0190674
+ 8.56e+10Hz -0.0041267 -0.0190774
+ 8.57e+10Hz -0.00415385 -0.0190873
+ 8.58e+10Hz -0.00418103 -0.0190972
+ 8.59e+10Hz -0.00420822 -0.0191071
+ 8.6e+10Hz -0.00423543 -0.0191168
+ 8.61e+10Hz -0.00426266 -0.0191266
+ 8.62e+10Hz -0.00428991 -0.0191362
+ 8.63e+10Hz -0.00431718 -0.0191458
+ 8.64e+10Hz -0.00434447 -0.0191554
+ 8.65e+10Hz -0.00437177 -0.0191648
+ 8.66e+10Hz -0.00439909 -0.0191742
+ 8.67e+10Hz -0.00442643 -0.0191836
+ 8.68e+10Hz -0.00445378 -0.0191929
+ 8.69e+10Hz -0.00448115 -0.0192021
+ 8.7e+10Hz -0.00450853 -0.0192112
+ 8.71e+10Hz -0.00453593 -0.0192203
+ 8.72e+10Hz -0.00456334 -0.0192293
+ 8.73e+10Hz -0.00459076 -0.0192383
+ 8.74e+10Hz -0.0046182 -0.0192472
+ 8.75e+10Hz -0.00464565 -0.019256
+ 8.76e+10Hz -0.00467311 -0.0192648
+ 8.77e+10Hz -0.00470059 -0.0192735
+ 8.78e+10Hz -0.00472807 -0.0192822
+ 8.79e+10Hz -0.00475556 -0.0192907
+ 8.8e+10Hz -0.00478307 -0.0192992
+ 8.81e+10Hz -0.00481058 -0.0193077
+ 8.82e+10Hz -0.00483811 -0.0193161
+ 8.83e+10Hz -0.00486564 -0.0193244
+ 8.84e+10Hz -0.00489318 -0.0193326
+ 8.85e+10Hz -0.00492072 -0.0193408
+ 8.86e+10Hz -0.00494828 -0.0193489
+ 8.87e+10Hz -0.00497583 -0.019357
+ 8.88e+10Hz -0.0050034 -0.0193649
+ 8.89e+10Hz -0.00503097 -0.0193729
+ 8.9e+10Hz -0.00505855 -0.0193807
+ 8.91e+10Hz -0.00508613 -0.0193885
+ 8.92e+10Hz -0.00511371 -0.0193962
+ 8.93e+10Hz -0.0051413 -0.0194039
+ 8.94e+10Hz -0.00516888 -0.0194115
+ 8.95e+10Hz -0.00519648 -0.019419
+ 8.96e+10Hz -0.00522407 -0.0194265
+ 8.97e+10Hz -0.00525166 -0.0194338
+ 8.98e+10Hz -0.00527926 -0.0194412
+ 8.99e+10Hz -0.00530685 -0.0194484
+ 9e+10Hz -0.00533445 -0.0194556
+ 9.01e+10Hz -0.00536204 -0.0194628
+ 9.02e+10Hz -0.00538963 -0.0194698
+ 9.03e+10Hz -0.00541723 -0.0194768
+ 9.04e+10Hz -0.00544481 -0.0194838
+ 9.05e+10Hz -0.0054724 -0.0194907
+ 9.06e+10Hz -0.00549998 -0.0194975
+ 9.07e+10Hz -0.00552756 -0.0195042
+ 9.08e+10Hz -0.00555514 -0.0195109
+ 9.09e+10Hz -0.00558271 -0.0195175
+ 9.1e+10Hz -0.00561028 -0.0195241
+ 9.11e+10Hz -0.00563784 -0.0195306
+ 9.12e+10Hz -0.00566539 -0.019537
+ 9.13e+10Hz -0.00569294 -0.0195433
+ 9.14e+10Hz -0.00572048 -0.0195497
+ 9.15e+10Hz -0.00574802 -0.0195559
+ 9.16e+10Hz -0.00577554 -0.0195621
+ 9.17e+10Hz -0.00580306 -0.0195682
+ 9.18e+10Hz -0.00583058 -0.0195742
+ 9.19e+10Hz -0.00585808 -0.0195802
+ 9.2e+10Hz -0.00588557 -0.0195862
+ 9.21e+10Hz -0.00591306 -0.019592
+ 9.22e+10Hz -0.00594053 -0.0195979
+ 9.23e+10Hz -0.005968 -0.0196036
+ 9.24e+10Hz -0.00599545 -0.0196093
+ 9.25e+10Hz -0.0060229 -0.0196149
+ 9.26e+10Hz -0.00605033 -0.0196205
+ 9.27e+10Hz -0.00607776 -0.019626
+ 9.28e+10Hz -0.00610517 -0.0196315
+ 9.29e+10Hz -0.00613257 -0.0196369
+ 9.3e+10Hz -0.00615996 -0.0196422
+ 9.31e+10Hz -0.00618733 -0.0196475
+ 9.32e+10Hz -0.0062147 -0.0196527
+ 9.33e+10Hz -0.00624205 -0.0196579
+ 9.34e+10Hz -0.00626938 -0.019663
+ 9.35e+10Hz -0.00629671 -0.0196681
+ 9.36e+10Hz -0.00632402 -0.0196731
+ 9.37e+10Hz -0.00635132 -0.019678
+ 9.38e+10Hz -0.0063786 -0.0196829
+ 9.39e+10Hz -0.00640587 -0.0196877
+ 9.4e+10Hz -0.00643313 -0.0196925
+ 9.41e+10Hz -0.00646037 -0.0196972
+ 9.42e+10Hz -0.0064876 -0.0197019
+ 9.43e+10Hz -0.00651481 -0.0197065
+ 9.44e+10Hz -0.00654201 -0.0197111
+ 9.45e+10Hz -0.00656919 -0.0197156
+ 9.46e+10Hz -0.00659636 -0.0197201
+ 9.47e+10Hz -0.00662351 -0.0197245
+ 9.48e+10Hz -0.00665065 -0.0197288
+ 9.49e+10Hz -0.00667778 -0.0197331
+ 9.5e+10Hz -0.00670488 -0.0197374
+ 9.51e+10Hz -0.00673198 -0.0197416
+ 9.52e+10Hz -0.00675905 -0.0197457
+ 9.53e+10Hz -0.00678612 -0.0197499
+ 9.54e+10Hz -0.00681316 -0.0197539
+ 9.55e+10Hz -0.0068402 -0.0197579
+ 9.56e+10Hz -0.00686721 -0.0197619
+ 9.57e+10Hz -0.00689421 -0.0197658
+ 9.58e+10Hz -0.0069212 -0.0197696
+ 9.59e+10Hz -0.00694817 -0.0197734
+ 9.6e+10Hz -0.00697512 -0.0197772
+ 9.61e+10Hz -0.00700206 -0.0197809
+ 9.62e+10Hz -0.00702899 -0.0197846
+ 9.63e+10Hz -0.00705589 -0.0197882
+ 9.64e+10Hz -0.00708279 -0.0197918
+ 9.65e+10Hz -0.00710967 -0.0197953
+ 9.66e+10Hz -0.00713653 -0.0197988
+ 9.67e+10Hz -0.00716338 -0.0198023
+ 9.68e+10Hz -0.00719021 -0.0198056
+ 9.69e+10Hz -0.00721703 -0.019809
+ 9.7e+10Hz -0.00724383 -0.0198123
+ 9.71e+10Hz -0.00727062 -0.0198156
+ 9.72e+10Hz -0.0072974 -0.0198188
+ 9.73e+10Hz -0.00732416 -0.0198219
+ 9.74e+10Hz -0.0073509 -0.0198251
+ 9.75e+10Hz -0.00737763 -0.0198281
+ 9.76e+10Hz -0.00740435 -0.0198312
+ 9.77e+10Hz -0.00743105 -0.0198342
+ 9.78e+10Hz -0.00745774 -0.0198371
+ 9.79e+10Hz -0.00748442 -0.01984
+ 9.8e+10Hz -0.00751108 -0.0198429
+ 9.81e+10Hz -0.00753773 -0.0198457
+ 9.82e+10Hz -0.00756437 -0.0198485
+ 9.83e+10Hz -0.00759099 -0.0198513
+ 9.84e+10Hz -0.0076176 -0.0198539
+ 9.85e+10Hz -0.0076442 -0.0198566
+ 9.86e+10Hz -0.00767078 -0.0198592
+ 9.87e+10Hz -0.00769736 -0.0198618
+ 9.88e+10Hz -0.00772392 -0.0198643
+ 9.89e+10Hz -0.00775047 -0.0198668
+ 9.9e+10Hz -0.007777 -0.0198693
+ 9.91e+10Hz -0.00780353 -0.0198717
+ 9.92e+10Hz -0.00783004 -0.019874
+ 9.93e+10Hz -0.00785654 -0.0198763
+ 9.94e+10Hz -0.00788303 -0.0198786
+ 9.95e+10Hz -0.00790951 -0.0198809
+ 9.96e+10Hz -0.00793598 -0.0198831
+ 9.97e+10Hz -0.00796244 -0.0198852
+ 9.98e+10Hz -0.00798889 -0.0198873
+ 9.99e+10Hz -0.00801533 -0.0198894
+ 1e+11Hz -0.00804175 -0.0198914
+ 1.001e+11Hz -0.00806817 -0.0198934
+ 1.002e+11Hz -0.00809458 -0.0198954
+ 1.003e+11Hz -0.00812098 -0.0198973
+ 1.004e+11Hz -0.00814737 -0.0198992
+ 1.005e+11Hz -0.00817375 -0.019901
+ 1.006e+11Hz -0.00820012 -0.0199028
+ 1.007e+11Hz -0.00822648 -0.0199045
+ 1.008e+11Hz -0.00825283 -0.0199063
+ 1.009e+11Hz -0.00827917 -0.0199079
+ 1.01e+11Hz -0.00830551 -0.0199095
+ 1.011e+11Hz -0.00833184 -0.0199111
+ 1.012e+11Hz -0.00835816 -0.0199127
+ 1.013e+11Hz -0.00838447 -0.0199142
+ 1.014e+11Hz -0.00841077 -0.0199156
+ 1.015e+11Hz -0.00843707 -0.019917
+ 1.016e+11Hz -0.00846336 -0.0199184
+ 1.017e+11Hz -0.00848964 -0.0199197
+ 1.018e+11Hz -0.00851591 -0.019921
+ 1.019e+11Hz -0.00854217 -0.0199223
+ 1.02e+11Hz -0.00856843 -0.0199235
+ 1.021e+11Hz -0.00859468 -0.0199246
+ 1.022e+11Hz -0.00862093 -0.0199257
+ 1.023e+11Hz -0.00864717 -0.0199268
+ 1.024e+11Hz -0.0086734 -0.0199278
+ 1.025e+11Hz -0.00869962 -0.0199288
+ 1.026e+11Hz -0.00872584 -0.0199298
+ 1.027e+11Hz -0.00875205 -0.0199307
+ 1.028e+11Hz -0.00877825 -0.0199315
+ 1.029e+11Hz -0.00880445 -0.0199323
+ 1.03e+11Hz -0.00883064 -0.0199331
+ 1.031e+11Hz -0.00885682 -0.0199338
+ 1.032e+11Hz -0.008883 -0.0199345
+ 1.033e+11Hz -0.00890917 -0.0199351
+ 1.034e+11Hz -0.00893534 -0.0199357
+ 1.035e+11Hz -0.00896149 -0.0199363
+ 1.036e+11Hz -0.00898764 -0.0199368
+ 1.037e+11Hz -0.00901379 -0.0199372
+ 1.038e+11Hz -0.00903993 -0.0199376
+ 1.039e+11Hz -0.00906606 -0.019938
+ 1.04e+11Hz -0.00909218 -0.0199383
+ 1.041e+11Hz -0.0091183 -0.0199385
+ 1.042e+11Hz -0.00914441 -0.0199388
+ 1.043e+11Hz -0.00917052 -0.0199389
+ 1.044e+11Hz -0.00919662 -0.019939
+ 1.045e+11Hz -0.00922271 -0.0199391
+ 1.046e+11Hz -0.00924879 -0.0199391
+ 1.047e+11Hz -0.00927487 -0.0199391
+ 1.048e+11Hz -0.00930094 -0.019939
+ 1.049e+11Hz -0.009327 -0.0199389
+ 1.05e+11Hz -0.00935305 -0.0199388
+ 1.051e+11Hz -0.0093791 -0.0199385
+ 1.052e+11Hz -0.00940514 -0.0199383
+ 1.053e+11Hz -0.00943117 -0.019938
+ 1.054e+11Hz -0.00945719 -0.0199376
+ 1.055e+11Hz -0.00948321 -0.0199372
+ 1.056e+11Hz -0.00950921 -0.0199367
+ 1.057e+11Hz -0.00953521 -0.0199362
+ 1.058e+11Hz -0.0095612 -0.0199356
+ 1.059e+11Hz -0.00958718 -0.019935
+ 1.06e+11Hz -0.00961315 -0.0199343
+ 1.061e+11Hz -0.00963911 -0.0199336
+ 1.062e+11Hz -0.00966506 -0.0199328
+ 1.063e+11Hz -0.009691 -0.019932
+ 1.064e+11Hz -0.00971693 -0.0199311
+ 1.065e+11Hz -0.00974285 -0.0199302
+ 1.066e+11Hz -0.00976876 -0.0199292
+ 1.067e+11Hz -0.00979465 -0.0199281
+ 1.068e+11Hz -0.00982054 -0.019927
+ 1.069e+11Hz -0.00984641 -0.0199259
+ 1.07e+11Hz -0.00987228 -0.0199247
+ 1.071e+11Hz -0.00989813 -0.0199234
+ 1.072e+11Hz -0.00992397 -0.0199221
+ 1.073e+11Hz -0.00994979 -0.0199208
+ 1.074e+11Hz -0.0099756 -0.0199194
+ 1.075e+11Hz -0.0100014 -0.0199179
+ 1.076e+11Hz -0.0100272 -0.0199164
+ 1.077e+11Hz -0.010053 -0.0199148
+ 1.078e+11Hz -0.0100787 -0.0199132
+ 1.079e+11Hz -0.0101045 -0.0199115
+ 1.08e+11Hz -0.0101302 -0.0199097
+ 1.081e+11Hz -0.0101559 -0.0199079
+ 1.082e+11Hz -0.0101816 -0.0199061
+ 1.083e+11Hz -0.0102073 -0.0199042
+ 1.084e+11Hz -0.0102329 -0.0199022
+ 1.085e+11Hz -0.0102586 -0.0199002
+ 1.086e+11Hz -0.0102842 -0.0198981
+ 1.087e+11Hz -0.0103098 -0.019896
+ 1.088e+11Hz -0.0103354 -0.0198938
+ 1.089e+11Hz -0.010361 -0.0198916
+ 1.09e+11Hz -0.0103865 -0.0198893
+ 1.091e+11Hz -0.0104121 -0.0198869
+ 1.092e+11Hz -0.0104376 -0.0198845
+ 1.093e+11Hz -0.0104631 -0.0198821
+ 1.094e+11Hz -0.0104886 -0.0198796
+ 1.095e+11Hz -0.010514 -0.019877
+ 1.096e+11Hz -0.0105394 -0.0198744
+ 1.097e+11Hz -0.0105648 -0.0198717
+ 1.098e+11Hz -0.0105902 -0.0198689
+ 1.099e+11Hz -0.0106156 -0.0198661
+ 1.1e+11Hz -0.0106409 -0.0198633
+ 1.101e+11Hz -0.0106663 -0.0198604
+ 1.102e+11Hz -0.0106916 -0.0198574
+ 1.103e+11Hz -0.0107168 -0.0198544
+ 1.104e+11Hz -0.0107421 -0.0198513
+ 1.105e+11Hz -0.0107673 -0.0198482
+ 1.106e+11Hz -0.0107925 -0.019845
+ 1.107e+11Hz -0.0108177 -0.0198418
+ 1.108e+11Hz -0.0108428 -0.0198385
+ 1.109e+11Hz -0.0108679 -0.0198351
+ 1.11e+11Hz -0.010893 -0.0198317
+ 1.111e+11Hz -0.0109181 -0.0198283
+ 1.112e+11Hz -0.0109431 -0.0198248
+ 1.113e+11Hz -0.0109681 -0.0198212
+ 1.114e+11Hz -0.0109931 -0.0198176
+ 1.115e+11Hz -0.0110181 -0.0198139
+ 1.116e+11Hz -0.011043 -0.0198102
+ 1.117e+11Hz -0.0110679 -0.0198064
+ 1.118e+11Hz -0.0110927 -0.0198026
+ 1.119e+11Hz -0.0111176 -0.0197987
+ 1.12e+11Hz -0.0111424 -0.0197947
+ 1.121e+11Hz -0.0111671 -0.0197908
+ 1.122e+11Hz -0.0111919 -0.0197867
+ 1.123e+11Hz -0.0112166 -0.0197826
+ 1.124e+11Hz -0.0112412 -0.0197785
+ 1.125e+11Hz -0.0112659 -0.0197743
+ 1.126e+11Hz -0.0112905 -0.01977
+ 1.127e+11Hz -0.011315 -0.0197657
+ 1.128e+11Hz -0.0113396 -0.0197614
+ 1.129e+11Hz -0.0113641 -0.019757
+ 1.13e+11Hz -0.0113886 -0.0197525
+ 1.131e+11Hz -0.011413 -0.019748
+ 1.132e+11Hz -0.0114374 -0.0197435
+ 1.133e+11Hz -0.0114618 -0.0197389
+ 1.134e+11Hz -0.0114861 -0.0197342
+ 1.135e+11Hz -0.0115104 -0.0197295
+ 1.136e+11Hz -0.0115346 -0.0197248
+ 1.137e+11Hz -0.0115588 -0.01972
+ 1.138e+11Hz -0.011583 -0.0197151
+ 1.139e+11Hz -0.0116072 -0.0197102
+ 1.14e+11Hz -0.0116313 -0.0197053
+ 1.141e+11Hz -0.0116553 -0.0197003
+ 1.142e+11Hz -0.0116794 -0.0196953
+ 1.143e+11Hz -0.0117034 -0.0196902
+ 1.144e+11Hz -0.0117273 -0.0196851
+ 1.145e+11Hz -0.0117512 -0.0196799
+ 1.146e+11Hz -0.0117751 -0.0196747
+ 1.147e+11Hz -0.011799 -0.0196695
+ 1.148e+11Hz -0.0118228 -0.0196642
+ 1.149e+11Hz -0.0118465 -0.0196588
+ 1.15e+11Hz -0.0118702 -0.0196534
+ 1.151e+11Hz -0.0118939 -0.019648
+ 1.152e+11Hz -0.0119176 -0.0196425
+ 1.153e+11Hz -0.0119412 -0.019637
+ 1.154e+11Hz -0.0119647 -0.0196315
+ 1.155e+11Hz -0.0119883 -0.0196259
+ 1.156e+11Hz -0.0120117 -0.0196202
+ 1.157e+11Hz -0.0120352 -0.0196146
+ 1.158e+11Hz -0.0120586 -0.0196088
+ 1.159e+11Hz -0.0120819 -0.0196031
+ 1.16e+11Hz -0.0121053 -0.0195973
+ 1.161e+11Hz -0.0121285 -0.0195914
+ 1.162e+11Hz -0.0121518 -0.0195856
+ 1.163e+11Hz -0.012175 -0.0195797
+ 1.164e+11Hz -0.0121981 -0.0195737
+ 1.165e+11Hz -0.0122212 -0.0195677
+ 1.166e+11Hz -0.0122443 -0.0195617
+ 1.167e+11Hz -0.0122673 -0.0195556
+ 1.168e+11Hz -0.0122903 -0.0195495
+ 1.169e+11Hz -0.0123133 -0.0195434
+ 1.17e+11Hz -0.0123362 -0.0195372
+ 1.171e+11Hz -0.012359 -0.019531
+ 1.172e+11Hz -0.0123819 -0.0195248
+ 1.173e+11Hz -0.0124047 -0.0195185
+ 1.174e+11Hz -0.0124274 -0.0195122
+ 1.175e+11Hz -0.0124501 -0.0195059
+ 1.176e+11Hz -0.0124728 -0.0194995
+ 1.177e+11Hz -0.0124954 -0.0194931
+ 1.178e+11Hz -0.012518 -0.0194866
+ 1.179e+11Hz -0.0125405 -0.0194802
+ 1.18e+11Hz -0.012563 -0.0194737
+ 1.181e+11Hz -0.0125854 -0.0194671
+ 1.182e+11Hz -0.0126079 -0.0194606
+ 1.183e+11Hz -0.0126302 -0.019454
+ 1.184e+11Hz -0.0126526 -0.0194473
+ 1.185e+11Hz -0.0126749 -0.0194407
+ 1.186e+11Hz -0.0126971 -0.019434
+ 1.187e+11Hz -0.0127193 -0.0194273
+ 1.188e+11Hz -0.0127415 -0.0194205
+ 1.189e+11Hz -0.0127636 -0.0194137
+ 1.19e+11Hz -0.0127857 -0.0194069
+ 1.191e+11Hz -0.0128078 -0.0194001
+ 1.192e+11Hz -0.0128298 -0.0193932
+ 1.193e+11Hz -0.0128518 -0.0193863
+ 1.194e+11Hz -0.0128737 -0.0193794
+ 1.195e+11Hz -0.0128956 -0.0193725
+ 1.196e+11Hz -0.0129175 -0.0193655
+ 1.197e+11Hz -0.0129393 -0.0193585
+ 1.198e+11Hz -0.0129611 -0.0193515
+ 1.199e+11Hz -0.0129828 -0.0193444
+ 1.2e+11Hz -0.0130045 -0.0193373
+ 1.201e+11Hz -0.0130262 -0.0193302
+ 1.202e+11Hz -0.0130478 -0.0193231
+ 1.203e+11Hz -0.0130694 -0.0193159
+ 1.204e+11Hz -0.0130909 -0.0193088
+ 1.205e+11Hz -0.0131125 -0.0193016
+ 1.206e+11Hz -0.0131339 -0.0192943
+ 1.207e+11Hz -0.0131554 -0.0192871
+ 1.208e+11Hz -0.0131768 -0.0192798
+ 1.209e+11Hz -0.0131982 -0.0192725
+ 1.21e+11Hz -0.0132195 -0.0192651
+ 1.211e+11Hz -0.0132408 -0.0192578
+ 1.212e+11Hz -0.013262 -0.0192504
+ 1.213e+11Hz -0.0132833 -0.019243
+ 1.214e+11Hz -0.0133045 -0.0192356
+ 1.215e+11Hz -0.0133256 -0.0192281
+ 1.216e+11Hz -0.0133467 -0.0192206
+ 1.217e+11Hz -0.0133678 -0.0192131
+ 1.218e+11Hz -0.0133889 -0.0192056
+ 1.219e+11Hz -0.0134099 -0.0191981
+ 1.22e+11Hz -0.0134309 -0.0191905
+ 1.221e+11Hz -0.0134518 -0.0191829
+ 1.222e+11Hz -0.0134727 -0.0191753
+ 1.223e+11Hz -0.0134936 -0.0191676
+ 1.224e+11Hz -0.0135144 -0.01916
+ 1.225e+11Hz -0.0135353 -0.0191523
+ 1.226e+11Hz -0.013556 -0.0191446
+ 1.227e+11Hz -0.0135768 -0.0191369
+ 1.228e+11Hz -0.0135975 -0.0191291
+ 1.229e+11Hz -0.0136182 -0.0191213
+ 1.23e+11Hz -0.0136388 -0.0191135
+ 1.231e+11Hz -0.0136594 -0.0191057
+ 1.232e+11Hz -0.01368 -0.0190978
+ 1.233e+11Hz -0.0137006 -0.0190899
+ 1.234e+11Hz -0.0137211 -0.0190821
+ 1.235e+11Hz -0.0137416 -0.0190741
+ 1.236e+11Hz -0.013762 -0.0190662
+ 1.237e+11Hz -0.0137825 -0.0190582
+ 1.238e+11Hz -0.0138028 -0.0190502
+ 1.239e+11Hz -0.0138232 -0.0190422
+ 1.24e+11Hz -0.0138435 -0.0190342
+ 1.241e+11Hz -0.0138638 -0.0190261
+ 1.242e+11Hz -0.0138841 -0.019018
+ 1.243e+11Hz -0.0139043 -0.0190099
+ 1.244e+11Hz -0.0139246 -0.0190018
+ 1.245e+11Hz -0.0139447 -0.0189936
+ 1.246e+11Hz -0.0139649 -0.0189854
+ 1.247e+11Hz -0.013985 -0.0189772
+ 1.248e+11Hz -0.0140051 -0.018969
+ 1.249e+11Hz -0.0140251 -0.0189607
+ 1.25e+11Hz -0.0140452 -0.0189524
+ 1.251e+11Hz -0.0140652 -0.0189441
+ 1.252e+11Hz -0.0140851 -0.0189358
+ 1.253e+11Hz -0.0141051 -0.0189274
+ 1.254e+11Hz -0.014125 -0.018919
+ 1.255e+11Hz -0.0141448 -0.0189106
+ 1.256e+11Hz -0.0141647 -0.0189022
+ 1.257e+11Hz -0.0141845 -0.0188937
+ 1.258e+11Hz -0.0142043 -0.0188852
+ 1.259e+11Hz -0.0142241 -0.0188767
+ 1.26e+11Hz -0.0142438 -0.0188681
+ 1.261e+11Hz -0.0142635 -0.0188596
+ 1.262e+11Hz -0.0142831 -0.018851
+ 1.263e+11Hz -0.0143028 -0.0188423
+ 1.264e+11Hz -0.0143224 -0.0188337
+ 1.265e+11Hz -0.014342 -0.018825
+ 1.266e+11Hz -0.0143615 -0.0188163
+ 1.267e+11Hz -0.014381 -0.0188076
+ 1.268e+11Hz -0.0144005 -0.0187988
+ 1.269e+11Hz -0.01442 -0.01879
+ 1.27e+11Hz -0.0144394 -0.0187812
+ 1.271e+11Hz -0.0144588 -0.0187724
+ 1.272e+11Hz -0.0144781 -0.0187635
+ 1.273e+11Hz -0.0144975 -0.0187546
+ 1.274e+11Hz -0.0145168 -0.0187456
+ 1.275e+11Hz -0.014536 -0.0187367
+ 1.276e+11Hz -0.0145553 -0.0187277
+ 1.277e+11Hz -0.0145745 -0.0187187
+ 1.278e+11Hz -0.0145937 -0.0187096
+ 1.279e+11Hz -0.0146128 -0.0187005
+ 1.28e+11Hz -0.0146319 -0.0186914
+ 1.281e+11Hz -0.014651 -0.0186823
+ 1.282e+11Hz -0.01467 -0.0186731
+ 1.283e+11Hz -0.014689 -0.0186639
+ 1.284e+11Hz -0.014708 -0.0186547
+ 1.285e+11Hz -0.014727 -0.0186454
+ 1.286e+11Hz -0.0147459 -0.0186362
+ 1.287e+11Hz -0.0147648 -0.0186268
+ 1.288e+11Hz -0.0147836 -0.0186175
+ 1.289e+11Hz -0.0148024 -0.0186081
+ 1.29e+11Hz -0.0148212 -0.0185987
+ 1.291e+11Hz -0.0148399 -0.0185892
+ 1.292e+11Hz -0.0148587 -0.0185798
+ 1.293e+11Hz -0.0148773 -0.0185703
+ 1.294e+11Hz -0.014896 -0.0185607
+ 1.295e+11Hz -0.0149146 -0.0185512
+ 1.296e+11Hz -0.0149331 -0.0185416
+ 1.297e+11Hz -0.0149517 -0.0185319
+ 1.298e+11Hz -0.0149701 -0.0185223
+ 1.299e+11Hz -0.0149886 -0.0185126
+ 1.3e+11Hz -0.015007 -0.0185028
+ 1.301e+11Hz -0.0150254 -0.0184931
+ 1.302e+11Hz -0.0150437 -0.0184833
+ 1.303e+11Hz -0.015062 -0.0184735
+ 1.304e+11Hz -0.0150803 -0.0184636
+ 1.305e+11Hz -0.0150985 -0.0184537
+ 1.306e+11Hz -0.0151167 -0.0184438
+ 1.307e+11Hz -0.0151349 -0.0184339
+ 1.308e+11Hz -0.015153 -0.0184239
+ 1.309e+11Hz -0.015171 -0.0184139
+ 1.31e+11Hz -0.0151891 -0.0184039
+ 1.311e+11Hz -0.0152071 -0.0183938
+ 1.312e+11Hz -0.015225 -0.0183837
+ 1.313e+11Hz -0.0152429 -0.0183735
+ 1.314e+11Hz -0.0152608 -0.0183634
+ 1.315e+11Hz -0.0152786 -0.0183532
+ 1.316e+11Hz -0.0152963 -0.0183429
+ 1.317e+11Hz -0.0153141 -0.0183327
+ 1.318e+11Hz -0.0153318 -0.0183224
+ 1.319e+11Hz -0.0153494 -0.0183121
+ 1.32e+11Hz -0.015367 -0.0183017
+ 1.321e+11Hz -0.0153846 -0.0182913
+ 1.322e+11Hz -0.0154021 -0.0182809
+ 1.323e+11Hz -0.0154195 -0.0182705
+ 1.324e+11Hz -0.0154369 -0.01826
+ 1.325e+11Hz -0.0154543 -0.0182495
+ 1.326e+11Hz -0.0154716 -0.018239
+ 1.327e+11Hz -0.0154889 -0.0182284
+ 1.328e+11Hz -0.0155061 -0.0182178
+ 1.329e+11Hz -0.0155233 -0.0182072
+ 1.33e+11Hz -0.0155404 -0.0181966
+ 1.331e+11Hz -0.0155575 -0.0181859
+ 1.332e+11Hz -0.0155745 -0.0181752
+ 1.333e+11Hz -0.0155915 -0.0181645
+ 1.334e+11Hz -0.0156085 -0.0181537
+ 1.335e+11Hz -0.0156253 -0.0181429
+ 1.336e+11Hz -0.0156422 -0.0181321
+ 1.337e+11Hz -0.0156589 -0.0181212
+ 1.338e+11Hz -0.0156757 -0.0181104
+ 1.339e+11Hz -0.0156923 -0.0180995
+ 1.34e+11Hz -0.015709 -0.0180886
+ 1.341e+11Hz -0.0157255 -0.0180776
+ 1.342e+11Hz -0.0157421 -0.0180666
+ 1.343e+11Hz -0.0157585 -0.0180556
+ 1.344e+11Hz -0.0157749 -0.0180446
+ 1.345e+11Hz -0.0157913 -0.0180336
+ 1.346e+11Hz -0.0158076 -0.0180225
+ 1.347e+11Hz -0.0158238 -0.0180114
+ 1.348e+11Hz -0.01584 -0.0180003
+ 1.349e+11Hz -0.0158562 -0.0179892
+ 1.35e+11Hz -0.0158723 -0.017978
+ 1.351e+11Hz -0.0158883 -0.0179668
+ 1.352e+11Hz -0.0159043 -0.0179556
+ 1.353e+11Hz -0.0159202 -0.0179444
+ 1.354e+11Hz -0.015936 -0.0179332
+ 1.355e+11Hz -0.0159518 -0.0179219
+ 1.356e+11Hz -0.0159676 -0.0179106
+ 1.357e+11Hz -0.0159833 -0.0178993
+ 1.358e+11Hz -0.0159989 -0.017888
+ 1.359e+11Hz -0.0160145 -0.0178766
+ 1.36e+11Hz -0.01603 -0.0178653
+ 1.361e+11Hz -0.0160454 -0.0178539
+ 1.362e+11Hz -0.0160608 -0.0178425
+ 1.363e+11Hz -0.0160761 -0.0178311
+ 1.364e+11Hz -0.0160914 -0.0178197
+ 1.365e+11Hz -0.0161066 -0.0178082
+ 1.366e+11Hz -0.0161218 -0.0177968
+ 1.367e+11Hz -0.0161369 -0.0177853
+ 1.368e+11Hz -0.0161519 -0.0177738
+ 1.369e+11Hz -0.0161669 -0.0177623
+ 1.37e+11Hz -0.0161818 -0.0177508
+ 1.371e+11Hz -0.0161967 -0.0177393
+ 1.372e+11Hz -0.0162115 -0.0177278
+ 1.373e+11Hz -0.0162262 -0.0177162
+ 1.374e+11Hz -0.0162409 -0.0177047
+ 1.375e+11Hz -0.0162555 -0.0176931
+ 1.376e+11Hz -0.0162701 -0.0176816
+ 1.377e+11Hz -0.0162845 -0.01767
+ 1.378e+11Hz -0.016299 -0.0176584
+ 1.379e+11Hz -0.0163133 -0.0176468
+ 1.38e+11Hz -0.0163277 -0.0176352
+ 1.381e+11Hz -0.0163419 -0.0176236
+ 1.382e+11Hz -0.0163561 -0.0176119
+ 1.383e+11Hz -0.0163702 -0.0176003
+ 1.384e+11Hz -0.0163843 -0.0175887
+ 1.385e+11Hz -0.0163983 -0.0175771
+ 1.386e+11Hz -0.0164122 -0.0175654
+ 1.387e+11Hz -0.0164261 -0.0175538
+ 1.388e+11Hz -0.0164399 -0.0175421
+ 1.389e+11Hz -0.0164537 -0.0175305
+ 1.39e+11Hz -0.0164674 -0.0175188
+ 1.391e+11Hz -0.016481 -0.0175072
+ 1.392e+11Hz -0.0164946 -0.0174955
+ 1.393e+11Hz -0.0165081 -0.0174839
+ 1.394e+11Hz -0.0165215 -0.0174722
+ 1.395e+11Hz -0.0165349 -0.0174606
+ 1.396e+11Hz -0.0165482 -0.0174489
+ 1.397e+11Hz -0.0165615 -0.0174373
+ 1.398e+11Hz -0.0165747 -0.0174256
+ 1.399e+11Hz -0.0165879 -0.017414
+ 1.4e+11Hz -0.0166009 -0.0174024
+ 1.401e+11Hz -0.016614 -0.0173907
+ 1.402e+11Hz -0.0166269 -0.0173791
+ 1.403e+11Hz -0.0166398 -0.0173675
+ 1.404e+11Hz -0.0166527 -0.0173559
+ 1.405e+11Hz -0.0166655 -0.0173443
+ 1.406e+11Hz -0.0166782 -0.0173327
+ 1.407e+11Hz -0.0166908 -0.0173211
+ 1.408e+11Hz -0.0167035 -0.0173095
+ 1.409e+11Hz -0.016716 -0.0172979
+ 1.41e+11Hz -0.0167285 -0.0172863
+ 1.411e+11Hz -0.0167409 -0.0172748
+ 1.412e+11Hz -0.0167533 -0.0172632
+ 1.413e+11Hz -0.0167656 -0.0172517
+ 1.414e+11Hz -0.0167779 -0.0172402
+ 1.415e+11Hz -0.01679 -0.0172286
+ 1.416e+11Hz -0.0168022 -0.0172171
+ 1.417e+11Hz -0.0168143 -0.0172056
+ 1.418e+11Hz -0.0168263 -0.0171942
+ 1.419e+11Hz -0.0168383 -0.0171827
+ 1.42e+11Hz -0.0168502 -0.0171712
+ 1.421e+11Hz -0.016862 -0.0171598
+ 1.422e+11Hz -0.0168738 -0.0171484
+ 1.423e+11Hz -0.0168856 -0.017137
+ 1.424e+11Hz -0.0168973 -0.0171256
+ 1.425e+11Hz -0.0169089 -0.0171142
+ 1.426e+11Hz -0.0169205 -0.0171028
+ 1.427e+11Hz -0.016932 -0.0170915
+ 1.428e+11Hz -0.0169435 -0.0170801
+ 1.429e+11Hz -0.0169549 -0.0170688
+ 1.43e+11Hz -0.0169662 -0.0170575
+ 1.431e+11Hz -0.0169775 -0.0170463
+ 1.432e+11Hz -0.0169888 -0.017035
+ 1.433e+11Hz -0.017 -0.0170238
+ 1.434e+11Hz -0.0170112 -0.0170125
+ 1.435e+11Hz -0.0170223 -0.0170013
+ 1.436e+11Hz -0.0170333 -0.0169902
+ 1.437e+11Hz -0.0170443 -0.016979
+ 1.438e+11Hz -0.0170553 -0.0169679
+ 1.439e+11Hz -0.0170661 -0.0169567
+ 1.44e+11Hz -0.017077 -0.0169456
+ 1.441e+11Hz -0.0170878 -0.0169346
+ 1.442e+11Hz -0.0170985 -0.0169235
+ 1.443e+11Hz -0.0171092 -0.0169125
+ 1.444e+11Hz -0.0171199 -0.0169015
+ 1.445e+11Hz -0.0171305 -0.0168905
+ 1.446e+11Hz -0.017141 -0.0168795
+ 1.447e+11Hz -0.0171515 -0.0168686
+ 1.448e+11Hz -0.017162 -0.0168576
+ 1.449e+11Hz -0.0171724 -0.0168468
+ 1.45e+11Hz -0.0171828 -0.0168359
+ 1.451e+11Hz -0.0171931 -0.016825
+ 1.452e+11Hz -0.0172033 -0.0168142
+ 1.453e+11Hz -0.0172136 -0.0168034
+ 1.454e+11Hz -0.0172238 -0.0167926
+ 1.455e+11Hz -0.0172339 -0.0167819
+ 1.456e+11Hz -0.017244 -0.0167712
+ 1.457e+11Hz -0.017254 -0.0167605
+ 1.458e+11Hz -0.017264 -0.0167498
+ 1.459e+11Hz -0.017274 -0.0167391
+ 1.46e+11Hz -0.0172839 -0.0167285
+ 1.461e+11Hz -0.0172938 -0.0167179
+ 1.462e+11Hz -0.0173036 -0.0167073
+ 1.463e+11Hz -0.0173134 -0.0166968
+ 1.464e+11Hz -0.0173231 -0.0166863
+ 1.465e+11Hz -0.0173328 -0.0166758
+ 1.466e+11Hz -0.0173425 -0.0166653
+ 1.467e+11Hz -0.0173521 -0.0166549
+ 1.468e+11Hz -0.0173617 -0.0166445
+ 1.469e+11Hz -0.0173712 -0.0166341
+ 1.47e+11Hz -0.0173807 -0.0166237
+ 1.471e+11Hz -0.0173902 -0.0166134
+ 1.472e+11Hz -0.0173996 -0.0166031
+ 1.473e+11Hz -0.017409 -0.0165928
+ 1.474e+11Hz -0.0174183 -0.0165826
+ 1.475e+11Hz -0.0174276 -0.0165723
+ 1.476e+11Hz -0.0174369 -0.0165622
+ 1.477e+11Hz -0.0174461 -0.016552
+ 1.478e+11Hz -0.0174553 -0.0165419
+ 1.479e+11Hz -0.0174644 -0.0165317
+ 1.48e+11Hz -0.0174736 -0.0165217
+ 1.481e+11Hz -0.0174826 -0.0165116
+ 1.482e+11Hz -0.0174917 -0.0165016
+ 1.483e+11Hz -0.0175007 -0.0164916
+ 1.484e+11Hz -0.0175096 -0.0164816
+ 1.485e+11Hz -0.0175186 -0.0164717
+ 1.486e+11Hz -0.0175275 -0.0164618
+ 1.487e+11Hz -0.0175363 -0.0164519
+ 1.488e+11Hz -0.0175451 -0.0164421
+ 1.489e+11Hz -0.0175539 -0.0164322
+ 1.49e+11Hz -0.0175627 -0.0164224
+ 1.491e+11Hz -0.0175714 -0.0164127
+ 1.492e+11Hz -0.0175801 -0.016403
+ 1.493e+11Hz -0.0175887 -0.0163932
+ 1.494e+11Hz -0.0175973 -0.0163836
+ 1.495e+11Hz -0.0176059 -0.0163739
+ 1.496e+11Hz -0.0176144 -0.0163643
+ 1.497e+11Hz -0.0176229 -0.0163547
+ 1.498e+11Hz -0.0176314 -0.0163452
+ 1.499e+11Hz -0.0176399 -0.0163356
+ 1.5e+11Hz -0.0176483 -0.0163261
+ 1.501e+11Hz -0.0176566 -0.0163167
+ 1.502e+11Hz -0.017665 -0.0163072
+ 1.503e+11Hz -0.0176733 -0.0162978
+ 1.504e+11Hz -0.0176816 -0.0162885
+ 1.505e+11Hz -0.0176898 -0.0162791
+ 1.506e+11Hz -0.017698 -0.0162698
+ 1.507e+11Hz -0.0177062 -0.0162605
+ 1.508e+11Hz -0.0177144 -0.0162513
+ 1.509e+11Hz -0.0177225 -0.016242
+ 1.51e+11Hz -0.0177305 -0.0162329
+ 1.511e+11Hz -0.0177386 -0.0162237
+ 1.512e+11Hz -0.0177466 -0.0162146
+ 1.513e+11Hz -0.0177546 -0.0162055
+ 1.514e+11Hz -0.0177626 -0.0161964
+ 1.515e+11Hz -0.0177705 -0.0161874
+ 1.516e+11Hz -0.0177784 -0.0161784
+ 1.517e+11Hz -0.0177862 -0.0161694
+ 1.518e+11Hz -0.0177941 -0.0161605
+ 1.519e+11Hz -0.0178019 -0.0161516
+ 1.52e+11Hz -0.0178096 -0.0161427
+ 1.521e+11Hz -0.0178174 -0.0161338
+ 1.522e+11Hz -0.0178251 -0.016125
+ 1.523e+11Hz -0.0178327 -0.0161163
+ 1.524e+11Hz -0.0178404 -0.0161075
+ 1.525e+11Hz -0.017848 -0.0160988
+ 1.526e+11Hz -0.0178556 -0.0160901
+ 1.527e+11Hz -0.0178631 -0.0160815
+ 1.528e+11Hz -0.0178707 -0.0160729
+ 1.529e+11Hz -0.0178781 -0.0160643
+ 1.53e+11Hz -0.0178856 -0.0160558
+ 1.531e+11Hz -0.017893 -0.0160473
+ 1.532e+11Hz -0.0179004 -0.0160388
+ 1.533e+11Hz -0.0179078 -0.0160304
+ 1.534e+11Hz -0.0179152 -0.016022
+ 1.535e+11Hz -0.0179225 -0.0160137
+ 1.536e+11Hz -0.0179298 -0.0160053
+ 1.537e+11Hz -0.017937 -0.0159971
+ 1.538e+11Hz -0.0179442 -0.0159888
+ 1.539e+11Hz -0.0179514 -0.0159806
+ 1.54e+11Hz -0.0179586 -0.0159724
+ 1.541e+11Hz -0.0179657 -0.0159643
+ 1.542e+11Hz -0.0179728 -0.0159562
+ 1.543e+11Hz -0.0179799 -0.0159481
+ 1.544e+11Hz -0.017987 -0.0159401
+ 1.545e+11Hz -0.017994 -0.0159321
+ 1.546e+11Hz -0.018001 -0.0159242
+ 1.547e+11Hz -0.018008 -0.0159163
+ 1.548e+11Hz -0.0180149 -0.0159084
+ 1.549e+11Hz -0.0180218 -0.0159006
+ 1.55e+11Hz -0.0180287 -0.0158928
+ 1.551e+11Hz -0.0180355 -0.0158851
+ 1.552e+11Hz -0.0180424 -0.0158774
+ 1.553e+11Hz -0.0180492 -0.0158697
+ 1.554e+11Hz -0.0180559 -0.0158621
+ 1.555e+11Hz -0.0180627 -0.0158546
+ 1.556e+11Hz -0.0180694 -0.015847
+ 1.557e+11Hz -0.0180761 -0.0158396
+ 1.558e+11Hz -0.0180828 -0.0158321
+ 1.559e+11Hz -0.0180894 -0.0158247
+ 1.56e+11Hz -0.018096 -0.0158174
+ 1.561e+11Hz -0.0181026 -0.0158101
+ 1.562e+11Hz -0.0181092 -0.0158028
+ 1.563e+11Hz -0.0181157 -0.0157956
+ 1.564e+11Hz -0.0181222 -0.0157885
+ 1.565e+11Hz -0.0181287 -0.0157814
+ 1.566e+11Hz -0.0181352 -0.0157743
+ 1.567e+11Hz -0.0181416 -0.0157673
+ 1.568e+11Hz -0.018148 -0.0157603
+ 1.569e+11Hz -0.0181544 -0.0157534
+ 1.57e+11Hz -0.0181608 -0.0157465
+ 1.571e+11Hz -0.0181672 -0.0157397
+ 1.572e+11Hz -0.0181735 -0.0157329
+ 1.573e+11Hz -0.0181798 -0.0157262
+ 1.574e+11Hz -0.0181861 -0.0157196
+ 1.575e+11Hz -0.0181924 -0.0157129
+ 1.576e+11Hz -0.0181986 -0.0157064
+ 1.577e+11Hz -0.0182048 -0.0156999
+ 1.578e+11Hz -0.018211 -0.0156934
+ 1.579e+11Hz -0.0182172 -0.015687
+ 1.58e+11Hz -0.0182234 -0.0156807
+ 1.581e+11Hz -0.0182295 -0.0156744
+ 1.582e+11Hz -0.0182357 -0.0156682
+ 1.583e+11Hz -0.0182418 -0.015662
+ 1.584e+11Hz -0.0182479 -0.0156559
+ 1.585e+11Hz -0.018254 -0.0156498
+ 1.586e+11Hz -0.01826 -0.0156438
+ 1.587e+11Hz -0.0182661 -0.0156379
+ 1.588e+11Hz -0.0182721 -0.015632
+ 1.589e+11Hz -0.0182781 -0.0156262
+ 1.59e+11Hz -0.0182842 -0.0156204
+ 1.591e+11Hz -0.0182901 -0.0156147
+ 1.592e+11Hz -0.0182961 -0.0156091
+ 1.593e+11Hz -0.0183021 -0.0156035
+ 1.594e+11Hz -0.0183081 -0.015598
+ 1.595e+11Hz -0.018314 -0.0155925
+ 1.596e+11Hz -0.01832 -0.0155871
+ 1.597e+11Hz -0.0183259 -0.0155818
+ 1.598e+11Hz -0.0183318 -0.0155765
+ 1.599e+11Hz -0.0183378 -0.0155713
+ 1.6e+11Hz -0.0183437 -0.0155662
+ 1.601e+11Hz -0.0183496 -0.0155611
+ 1.602e+11Hz -0.0183555 -0.0155561
+ 1.603e+11Hz -0.0183614 -0.0155512
+ 1.604e+11Hz -0.0183673 -0.0155463
+ 1.605e+11Hz -0.0183732 -0.0155415
+ 1.606e+11Hz -0.0183791 -0.0155368
+ 1.607e+11Hz -0.018385 -0.0155321
+ 1.608e+11Hz -0.0183909 -0.0155275
+ 1.609e+11Hz -0.0183967 -0.0155229
+ 1.61e+11Hz -0.0184026 -0.0155185
+ 1.611e+11Hz -0.0184085 -0.0155141
+ 1.612e+11Hz -0.0184144 -0.0155098
+ 1.613e+11Hz -0.0184204 -0.0155055
+ 1.614e+11Hz -0.0184263 -0.0155013
+ 1.615e+11Hz -0.0184322 -0.0154972
+ 1.616e+11Hz -0.0184381 -0.0154932
+ 1.617e+11Hz -0.0184441 -0.0154892
+ 1.618e+11Hz -0.01845 -0.0154853
+ 1.619e+11Hz -0.018456 -0.0154814
+ 1.62e+11Hz -0.0184619 -0.0154777
+ 1.621e+11Hz -0.0184679 -0.015474
+ 1.622e+11Hz -0.0184739 -0.0154704
+ 1.623e+11Hz -0.0184799 -0.0154668
+ 1.624e+11Hz -0.0184859 -0.0154634
+ 1.625e+11Hz -0.018492 -0.01546
+ 1.626e+11Hz -0.018498 -0.0154567
+ 1.627e+11Hz -0.0185041 -0.0154534
+ 1.628e+11Hz -0.0185102 -0.0154502
+ 1.629e+11Hz -0.0185164 -0.0154471
+ 1.63e+11Hz -0.0185225 -0.0154441
+ 1.631e+11Hz -0.0185287 -0.0154411
+ 1.632e+11Hz -0.0185349 -0.0154383
+ 1.633e+11Hz -0.0185411 -0.0154354
+ 1.634e+11Hz -0.0185473 -0.0154327
+ 1.635e+11Hz -0.0185536 -0.01543
+ 1.636e+11Hz -0.0185599 -0.0154275
+ 1.637e+11Hz -0.0185663 -0.0154249
+ 1.638e+11Hz -0.0185726 -0.0154225
+ 1.639e+11Hz -0.018579 -0.0154201
+ 1.64e+11Hz -0.0185855 -0.0154178
+ 1.641e+11Hz -0.018592 -0.0154156
+ 1.642e+11Hz -0.0185985 -0.0154135
+ 1.643e+11Hz -0.018605 -0.0154114
+ 1.644e+11Hz -0.0186116 -0.0154094
+ 1.645e+11Hz -0.0186183 -0.0154075
+ 1.646e+11Hz -0.0186249 -0.0154056
+ 1.647e+11Hz -0.0186316 -0.0154038
+ 1.648e+11Hz -0.0186384 -0.0154021
+ 1.649e+11Hz -0.0186452 -0.0154005
+ 1.65e+11Hz -0.0186521 -0.0153989
+ 1.651e+11Hz -0.018659 -0.0153974
+ 1.652e+11Hz -0.0186659 -0.0153959
+ 1.653e+11Hz -0.0186729 -0.0153946
+ 1.654e+11Hz -0.01868 -0.0153933
+ 1.655e+11Hz -0.0186871 -0.0153921
+ 1.656e+11Hz -0.0186943 -0.0153909
+ 1.657e+11Hz -0.0187015 -0.0153898
+ 1.658e+11Hz -0.0187088 -0.0153888
+ 1.659e+11Hz -0.0187161 -0.0153878
+ 1.66e+11Hz -0.0187235 -0.015387
+ 1.661e+11Hz -0.018731 -0.0153861
+ 1.662e+11Hz -0.0187385 -0.0153854
+ 1.663e+11Hz -0.0187461 -0.0153847
+ 1.664e+11Hz -0.0187538 -0.0153841
+ 1.665e+11Hz -0.0187615 -0.0153835
+ 1.666e+11Hz -0.0187693 -0.015383
+ 1.667e+11Hz -0.0187771 -0.0153826
+ 1.668e+11Hz -0.0187851 -0.0153822
+ 1.669e+11Hz -0.0187931 -0.0153819
+ 1.67e+11Hz -0.0188011 -0.0153816
+ 1.671e+11Hz -0.0188093 -0.0153814
+ 1.672e+11Hz -0.0188175 -0.0153813
+ 1.673e+11Hz -0.0188258 -0.0153812
+ 1.674e+11Hz -0.0188342 -0.0153812
+ 1.675e+11Hz -0.0188426 -0.0153812
+ 1.676e+11Hz -0.0188512 -0.0153813
+ 1.677e+11Hz -0.0188598 -0.0153814
+ 1.678e+11Hz -0.0188685 -0.0153816
+ 1.679e+11Hz -0.0188773 -0.0153818
+ 1.68e+11Hz -0.0188861 -0.0153821
+ 1.681e+11Hz -0.0188951 -0.0153825
+ 1.682e+11Hz -0.0189041 -0.0153828
+ 1.683e+11Hz -0.0189132 -0.0153833
+ 1.684e+11Hz -0.0189225 -0.0153837
+ 1.685e+11Hz -0.0189318 -0.0153843
+ 1.686e+11Hz -0.0189412 -0.0153848
+ 1.687e+11Hz -0.0189506 -0.0153854
+ 1.688e+11Hz -0.0189602 -0.0153861
+ 1.689e+11Hz -0.0189699 -0.0153868
+ 1.69e+11Hz -0.0189797 -0.0153875
+ 1.691e+11Hz -0.0189895 -0.0153883
+ 1.692e+11Hz -0.0189995 -0.0153891
+ 1.693e+11Hz -0.0190095 -0.0153899
+ 1.694e+11Hz -0.0190197 -0.0153908
+ 1.695e+11Hz -0.01903 -0.0153917
+ 1.696e+11Hz -0.0190403 -0.0153926
+ 1.697e+11Hz -0.0190508 -0.0153936
+ 1.698e+11Hz -0.0190613 -0.0153946
+ 1.699e+11Hz -0.019072 -0.0153956
+ 1.7e+11Hz -0.0190828 -0.0153966
+ 1.701e+11Hz -0.0190936 -0.0153977
+ 1.702e+11Hz -0.0191046 -0.0153988
+ 1.703e+11Hz -0.0191157 -0.0153999
+ 1.704e+11Hz -0.0191269 -0.015401
+ 1.705e+11Hz -0.0191382 -0.0154022
+ 1.706e+11Hz -0.0191496 -0.0154034
+ 1.707e+11Hz -0.0191611 -0.0154045
+ 1.708e+11Hz -0.0191727 -0.0154057
+ 1.709e+11Hz -0.0191844 -0.0154069
+ 1.71e+11Hz -0.0191963 -0.0154081
+ 1.711e+11Hz -0.0192082 -0.0154094
+ 1.712e+11Hz -0.0192203 -0.0154106
+ 1.713e+11Hz -0.0192325 -0.0154118
+ 1.714e+11Hz -0.0192447 -0.0154131
+ 1.715e+11Hz -0.0192571 -0.0154143
+ 1.716e+11Hz -0.0192696 -0.0154155
+ 1.717e+11Hz -0.0192823 -0.0154168
+ 1.718e+11Hz -0.019295 -0.015418
+ 1.719e+11Hz -0.0193079 -0.0154192
+ 1.72e+11Hz -0.0193208 -0.0154205
+ 1.721e+11Hz -0.0193339 -0.0154217
+ 1.722e+11Hz -0.0193471 -0.0154229
+ 1.723e+11Hz -0.0193604 -0.0154241
+ 1.724e+11Hz -0.0193738 -0.0154252
+ 1.725e+11Hz -0.0193874 -0.0154264
+ 1.726e+11Hz -0.019401 -0.0154276
+ 1.727e+11Hz -0.0194148 -0.0154287
+ 1.728e+11Hz -0.0194287 -0.0154298
+ 1.729e+11Hz -0.0194427 -0.0154309
+ 1.73e+11Hz -0.0194568 -0.0154319
+ 1.731e+11Hz -0.019471 -0.015433
+ 1.732e+11Hz -0.0194854 -0.015434
+ 1.733e+11Hz -0.0194999 -0.015435
+ 1.734e+11Hz -0.0195144 -0.0154359
+ 1.735e+11Hz -0.0195291 -0.0154368
+ 1.736e+11Hz -0.0195439 -0.0154377
+ 1.737e+11Hz -0.0195589 -0.0154386
+ 1.738e+11Hz -0.0195739 -0.0154394
+ 1.739e+11Hz -0.019589 -0.0154402
+ 1.74e+11Hz -0.0196043 -0.0154409
+ 1.741e+11Hz -0.0196197 -0.0154416
+ 1.742e+11Hz -0.0196352 -0.0154422
+ 1.743e+11Hz -0.0196508 -0.0154428
+ 1.744e+11Hz -0.0196665 -0.0154434
+ 1.745e+11Hz -0.0196823 -0.0154439
+ 1.746e+11Hz -0.0196983 -0.0154443
+ 1.747e+11Hz -0.0197143 -0.0154447
+ 1.748e+11Hz -0.0197305 -0.015445
+ 1.749e+11Hz -0.0197468 -0.0154453
+ 1.75e+11Hz -0.0197632 -0.0154455
+ 1.751e+11Hz -0.0197797 -0.0154457
+ 1.752e+11Hz -0.0197963 -0.0154458
+ 1.753e+11Hz -0.019813 -0.0154459
+ 1.754e+11Hz -0.0198298 -0.0154458
+ 1.755e+11Hz -0.0198467 -0.0154457
+ 1.756e+11Hz -0.0198637 -0.0154456
+ 1.757e+11Hz -0.0198809 -0.0154453
+ 1.758e+11Hz -0.0198981 -0.015445
+ 1.759e+11Hz -0.0199154 -0.0154447
+ 1.76e+11Hz -0.0199329 -0.0154442
+ 1.761e+11Hz -0.0199504 -0.0154437
+ 1.762e+11Hz -0.0199681 -0.0154431
+ 1.763e+11Hz -0.0199858 -0.0154424
+ 1.764e+11Hz -0.0200037 -0.0154416
+ 1.765e+11Hz -0.0200216 -0.0154408
+ 1.766e+11Hz -0.0200397 -0.0154399
+ 1.767e+11Hz -0.0200578 -0.0154389
+ 1.768e+11Hz -0.020076 -0.0154378
+ 1.769e+11Hz -0.0200943 -0.0154366
+ 1.77e+11Hz -0.0201128 -0.0154353
+ 1.771e+11Hz -0.0201313 -0.0154339
+ 1.772e+11Hz -0.0201499 -0.0154325
+ 1.773e+11Hz -0.0201685 -0.0154309
+ 1.774e+11Hz -0.0201873 -0.0154293
+ 1.775e+11Hz -0.0202062 -0.0154275
+ 1.776e+11Hz -0.0202251 -0.0154257
+ 1.777e+11Hz -0.0202442 -0.0154237
+ 1.778e+11Hz -0.0202633 -0.0154217
+ 1.779e+11Hz -0.0202825 -0.0154196
+ 1.78e+11Hz -0.0203018 -0.0154173
+ 1.781e+11Hz -0.0203211 -0.015415
+ 1.782e+11Hz -0.0203406 -0.0154125
+ 1.783e+11Hz -0.0203601 -0.01541
+ 1.784e+11Hz -0.0203797 -0.0154073
+ 1.785e+11Hz -0.0203993 -0.0154045
+ 1.786e+11Hz -0.0204191 -0.0154016
+ 1.787e+11Hz -0.0204389 -0.0153986
+ 1.788e+11Hz -0.0204588 -0.0153955
+ 1.789e+11Hz -0.0204787 -0.0153923
+ 1.79e+11Hz -0.0204987 -0.015389
+ 1.791e+11Hz -0.0205188 -0.0153855
+ 1.792e+11Hz -0.0205389 -0.015382
+ 1.793e+11Hz -0.0205592 -0.0153783
+ 1.794e+11Hz -0.0205794 -0.0153745
+ 1.795e+11Hz -0.0205997 -0.0153706
+ 1.796e+11Hz -0.0206201 -0.0153666
+ 1.797e+11Hz -0.0206406 -0.0153624
+ 1.798e+11Hz -0.0206611 -0.0153581
+ 1.799e+11Hz -0.0206816 -0.0153538
+ 1.8e+11Hz -0.0207022 -0.0153492
+ 1.801e+11Hz -0.0207229 -0.0153446
+ 1.802e+11Hz -0.0207436 -0.0153399
+ 1.803e+11Hz -0.0207643 -0.015335
+ 1.804e+11Hz -0.0207851 -0.01533
+ 1.805e+11Hz -0.020806 -0.0153248
+ 1.806e+11Hz -0.0208269 -0.0153196
+ 1.807e+11Hz -0.0208478 -0.0153142
+ 1.808e+11Hz -0.0208688 -0.0153087
+ 1.809e+11Hz -0.0208898 -0.015303
+ 1.81e+11Hz -0.0209108 -0.0152973
+ 1.811e+11Hz -0.0209319 -0.0152914
+ 1.812e+11Hz -0.020953 -0.0152854
+ 1.813e+11Hz -0.0209741 -0.0152792
+ 1.814e+11Hz -0.0209953 -0.0152729
+ 1.815e+11Hz -0.0210165 -0.0152665
+ 1.816e+11Hz -0.0210377 -0.01526
+ 1.817e+11Hz -0.0210589 -0.0152533
+ 1.818e+11Hz -0.0210802 -0.0152465
+ 1.819e+11Hz -0.0211015 -0.0152396
+ 1.82e+11Hz -0.0211228 -0.0152325
+ 1.821e+11Hz -0.0211441 -0.0152253
+ 1.822e+11Hz -0.0211655 -0.015218
+ 1.823e+11Hz -0.0211868 -0.0152105
+ 1.824e+11Hz -0.0212082 -0.0152029
+ 1.825e+11Hz -0.0212296 -0.0151952
+ 1.826e+11Hz -0.021251 -0.0151874
+ 1.827e+11Hz -0.0212724 -0.0151794
+ 1.828e+11Hz -0.0212938 -0.0151713
+ 1.829e+11Hz -0.0213152 -0.015163
+ 1.83e+11Hz -0.0213367 -0.0151546
+ 1.831e+11Hz -0.0213581 -0.0151461
+ 1.832e+11Hz -0.0213795 -0.0151375
+ 1.833e+11Hz -0.0214009 -0.0151287
+ 1.834e+11Hz -0.0214223 -0.0151198
+ 1.835e+11Hz -0.0214438 -0.0151107
+ 1.836e+11Hz -0.0214652 -0.0151016
+ 1.837e+11Hz -0.0214866 -0.0150923
+ 1.838e+11Hz -0.021508 -0.0150828
+ 1.839e+11Hz -0.0215293 -0.0150733
+ 1.84e+11Hz -0.0215507 -0.0150636
+ 1.841e+11Hz -0.0215721 -0.0150538
+ 1.842e+11Hz -0.0215934 -0.0150438
+ 1.843e+11Hz -0.0216147 -0.0150337
+ 1.844e+11Hz -0.021636 -0.0150235
+ 1.845e+11Hz -0.0216573 -0.0150132
+ 1.846e+11Hz -0.0216786 -0.0150027
+ 1.847e+11Hz -0.0216998 -0.0149921
+ 1.848e+11Hz -0.021721 -0.0149814
+ 1.849e+11Hz -0.0217422 -0.0149705
+ 1.85e+11Hz -0.0217634 -0.0149595
+ 1.851e+11Hz -0.0217845 -0.0149484
+ 1.852e+11Hz -0.0218057 -0.0149372
+ 1.853e+11Hz -0.0218267 -0.0149258
+ 1.854e+11Hz -0.0218478 -0.0149144
+ 1.855e+11Hz -0.0218688 -0.0149028
+ 1.856e+11Hz -0.0218898 -0.014891
+ 1.857e+11Hz -0.0219107 -0.0148792
+ 1.858e+11Hz -0.0219316 -0.0148672
+ 1.859e+11Hz -0.0219525 -0.0148551
+ 1.86e+11Hz -0.0219733 -0.0148429
+ 1.861e+11Hz -0.0219941 -0.0148306
+ 1.862e+11Hz -0.0220148 -0.0148181
+ 1.863e+11Hz -0.0220355 -0.0148055
+ 1.864e+11Hz -0.0220561 -0.0147928
+ 1.865e+11Hz -0.0220767 -0.01478
+ 1.866e+11Hz -0.0220973 -0.0147671
+ 1.867e+11Hz -0.0221178 -0.014754
+ 1.868e+11Hz -0.0221382 -0.0147409
+ 1.869e+11Hz -0.0221586 -0.0147276
+ 1.87e+11Hz -0.022179 -0.0147142
+ 1.871e+11Hz -0.0221993 -0.0147007
+ 1.872e+11Hz -0.0222195 -0.0146871
+ 1.873e+11Hz -0.0222397 -0.0146734
+ 1.874e+11Hz -0.0222598 -0.0146595
+ 1.875e+11Hz -0.0222799 -0.0146456
+ 1.876e+11Hz -0.0222999 -0.0146315
+ 1.877e+11Hz -0.0223198 -0.0146174
+ 1.878e+11Hz -0.0223397 -0.0146031
+ 1.879e+11Hz -0.0223595 -0.0145887
+ 1.88e+11Hz -0.0223793 -0.0145742
+ 1.881e+11Hz -0.022399 -0.0145597
+ 1.882e+11Hz -0.0224186 -0.014545
+ 1.883e+11Hz -0.0224381 -0.0145302
+ 1.884e+11Hz -0.0224576 -0.0145153
+ 1.885e+11Hz -0.022477 -0.0145003
+ 1.886e+11Hz -0.0224964 -0.0144852
+ 1.887e+11Hz -0.0225157 -0.01447
+ 1.888e+11Hz -0.0225349 -0.0144547
+ 1.889e+11Hz -0.022554 -0.0144393
+ 1.89e+11Hz -0.0225731 -0.0144238
+ 1.891e+11Hz -0.0225921 -0.0144082
+ 1.892e+11Hz -0.022611 -0.0143926
+ 1.893e+11Hz -0.0226298 -0.0143768
+ 1.894e+11Hz -0.0226486 -0.0143609
+ 1.895e+11Hz -0.0226673 -0.014345
+ 1.896e+11Hz -0.0226859 -0.0143289
+ 1.897e+11Hz -0.0227044 -0.0143128
+ 1.898e+11Hz -0.0227228 -0.0142966
+ 1.899e+11Hz -0.0227412 -0.0142803
+ 1.9e+11Hz -0.0227595 -0.0142639
+ 1.901e+11Hz -0.0227777 -0.0142474
+ 1.902e+11Hz -0.0227958 -0.0142308
+ 1.903e+11Hz -0.0228138 -0.0142142
+ 1.904e+11Hz -0.0228318 -0.0141975
+ 1.905e+11Hz -0.0228496 -0.0141807
+ 1.906e+11Hz -0.0228674 -0.0141638
+ 1.907e+11Hz -0.0228851 -0.0141468
+ 1.908e+11Hz -0.0229027 -0.0141298
+ 1.909e+11Hz -0.0229203 -0.0141127
+ 1.91e+11Hz -0.0229377 -0.0140955
+ 1.911e+11Hz -0.022955 -0.0140782
+ 1.912e+11Hz -0.0229723 -0.0140609
+ 1.913e+11Hz -0.0229894 -0.0140434
+ 1.914e+11Hz -0.0230065 -0.014026
+ 1.915e+11Hz -0.0230235 -0.0140084
+ 1.916e+11Hz -0.0230404 -0.0139908
+ 1.917e+11Hz -0.0230572 -0.0139731
+ 1.918e+11Hz -0.0230739 -0.0139553
+ 1.919e+11Hz -0.0230905 -0.0139375
+ 1.92e+11Hz -0.0231071 -0.0139196
+ 1.921e+11Hz -0.0231235 -0.0139017
+ 1.922e+11Hz -0.0231398 -0.0138837
+ 1.923e+11Hz -0.0231561 -0.0138656
+ 1.924e+11Hz -0.0231722 -0.0138475
+ 1.925e+11Hz -0.0231883 -0.0138293
+ 1.926e+11Hz -0.0232042 -0.013811
+ 1.927e+11Hz -0.0232201 -0.0137927
+ 1.928e+11Hz -0.0232359 -0.0137744
+ 1.929e+11Hz -0.0232516 -0.013756
+ 1.93e+11Hz -0.0232671 -0.0137375
+ 1.931e+11Hz -0.0232826 -0.013719
+ 1.932e+11Hz -0.023298 -0.0137004
+ 1.933e+11Hz -0.0233133 -0.0136818
+ 1.934e+11Hz -0.0233285 -0.0136631
+ 1.935e+11Hz -0.0233435 -0.0136444
+ 1.936e+11Hz -0.0233585 -0.0136257
+ 1.937e+11Hz -0.0233734 -0.0136069
+ 1.938e+11Hz -0.0233882 -0.013588
+ 1.939e+11Hz -0.0234029 -0.0135691
+ 1.94e+11Hz -0.0234175 -0.0135502
+ 1.941e+11Hz -0.023432 -0.0135312
+ 1.942e+11Hz -0.0234464 -0.0135122
+ 1.943e+11Hz -0.0234607 -0.0134932
+ 1.944e+11Hz -0.0234749 -0.0134741
+ 1.945e+11Hz -0.023489 -0.013455
+ 1.946e+11Hz -0.023503 -0.0134358
+ 1.947e+11Hz -0.0235169 -0.0134167
+ 1.948e+11Hz -0.0235307 -0.0133974
+ 1.949e+11Hz -0.0235444 -0.0133782
+ 1.95e+11Hz -0.023558 -0.0133589
+ 1.951e+11Hz -0.0235714 -0.0133396
+ 1.952e+11Hz -0.0235848 -0.0133203
+ 1.953e+11Hz -0.0235981 -0.0133009
+ 1.954e+11Hz -0.0236113 -0.0132815
+ 1.955e+11Hz -0.0236244 -0.0132621
+ 1.956e+11Hz -0.0236374 -0.0132427
+ 1.957e+11Hz -0.0236503 -0.0132232
+ 1.958e+11Hz -0.0236631 -0.0132038
+ 1.959e+11Hz -0.0236758 -0.0131843
+ 1.96e+11Hz -0.0236884 -0.0131648
+ 1.961e+11Hz -0.0237009 -0.0131453
+ 1.962e+11Hz -0.0237132 -0.0131257
+ 1.963e+11Hz -0.0237255 -0.0131062
+ 1.964e+11Hz -0.0237377 -0.0130866
+ 1.965e+11Hz -0.0237498 -0.013067
+ 1.966e+11Hz -0.0237618 -0.0130474
+ 1.967e+11Hz -0.0237737 -0.0130278
+ 1.968e+11Hz -0.0237855 -0.0130082
+ 1.969e+11Hz -0.0237972 -0.0129886
+ 1.97e+11Hz -0.0238088 -0.012969
+ 1.971e+11Hz -0.0238202 -0.0129494
+ 1.972e+11Hz -0.0238316 -0.0129297
+ 1.973e+11Hz -0.0238429 -0.0129101
+ 1.974e+11Hz -0.0238541 -0.0128905
+ 1.975e+11Hz -0.0238652 -0.0128709
+ 1.976e+11Hz -0.0238762 -0.0128512
+ 1.977e+11Hz -0.0238871 -0.0128316
+ 1.978e+11Hz -0.0238979 -0.012812
+ 1.979e+11Hz -0.0239087 -0.0127924
+ 1.98e+11Hz -0.0239193 -0.0127728
+ 1.981e+11Hz -0.0239298 -0.0127532
+ 1.982e+11Hz -0.0239402 -0.0127336
+ 1.983e+11Hz -0.0239505 -0.012714
+ 1.984e+11Hz -0.0239608 -0.0126944
+ 1.985e+11Hz -0.0239709 -0.0126749
+ 1.986e+11Hz -0.023981 -0.0126553
+ 1.987e+11Hz -0.0239909 -0.0126358
+ 1.988e+11Hz -0.0240008 -0.0126163
+ 1.989e+11Hz -0.0240105 -0.0125968
+ 1.99e+11Hz -0.0240202 -0.0125773
+ 1.991e+11Hz -0.0240298 -0.0125579
+ 1.992e+11Hz -0.0240393 -0.0125385
+ 1.993e+11Hz -0.0240487 -0.012519
+ 1.994e+11Hz -0.024058 -0.0124997
+ 1.995e+11Hz -0.0240672 -0.0124803
+ 1.996e+11Hz -0.0240764 -0.0124609
+ 1.997e+11Hz -0.0240854 -0.0124416
+ 1.998e+11Hz -0.0240944 -0.0124224
+ 1.999e+11Hz -0.0241033 -0.0124031
+ 2e+11Hz -0.0241121 -0.0123839
+ 2.001e+11Hz -0.0241208 -0.0123647
+ 2.002e+11Hz -0.0241294 -0.0123455
+ 2.003e+11Hz -0.0241379 -0.0123264
+ 2.004e+11Hz -0.0241464 -0.0123073
+ 2.005e+11Hz -0.0241548 -0.0122883
+ 2.006e+11Hz -0.0241631 -0.0122693
+ 2.007e+11Hz -0.0241713 -0.0122503
+ 2.008e+11Hz -0.0241794 -0.0122313
+ 2.009e+11Hz -0.0241875 -0.0122124
+ 2.01e+11Hz -0.0241955 -0.0121936
+ 2.011e+11Hz -0.0242034 -0.0121748
+ 2.012e+11Hz -0.0242112 -0.012156
+ 2.013e+11Hz -0.024219 -0.0121373
+ 2.014e+11Hz -0.0242267 -0.0121186
+ 2.015e+11Hz -0.0242343 -0.0121
+ 2.016e+11Hz -0.0242418 -0.0120814
+ 2.017e+11Hz -0.0242493 -0.0120629
+ 2.018e+11Hz -0.0242567 -0.0120444
+ 2.019e+11Hz -0.024264 -0.012026
+ 2.02e+11Hz -0.0242713 -0.0120076
+ 2.021e+11Hz -0.0242785 -0.0119893
+ 2.022e+11Hz -0.0242856 -0.011971
+ 2.023e+11Hz -0.0242927 -0.0119528
+ 2.024e+11Hz -0.0242997 -0.0119347
+ 2.025e+11Hz -0.0243067 -0.0119166
+ 2.026e+11Hz -0.0243136 -0.0118985
+ 2.027e+11Hz -0.0243204 -0.0118805
+ 2.028e+11Hz -0.0243272 -0.0118626
+ 2.029e+11Hz -0.0243339 -0.0118448
+ 2.03e+11Hz -0.0243406 -0.011827
+ 2.031e+11Hz -0.0243472 -0.0118093
+ 2.032e+11Hz -0.0243538 -0.0117916
+ 2.033e+11Hz -0.0243603 -0.011774
+ 2.034e+11Hz -0.0243668 -0.0117564
+ 2.035e+11Hz -0.0243732 -0.011739
+ 2.036e+11Hz -0.0243796 -0.0117216
+ 2.037e+11Hz -0.0243859 -0.0117042
+ 2.038e+11Hz -0.0243922 -0.011687
+ 2.039e+11Hz -0.0243984 -0.0116698
+ 2.04e+11Hz -0.0244046 -0.0116526
+ 2.041e+11Hz -0.0244108 -0.0116356
+ 2.042e+11Hz -0.024417 -0.0116186
+ 2.043e+11Hz -0.0244231 -0.0116017
+ 2.044e+11Hz -0.0244291 -0.0115848
+ 2.045e+11Hz -0.0244352 -0.0115681
+ 2.046e+11Hz -0.0244412 -0.0115514
+ 2.047e+11Hz -0.0244472 -0.0115348
+ 2.048e+11Hz -0.0244531 -0.0115182
+ 2.049e+11Hz -0.0244591 -0.0115017
+ 2.05e+11Hz -0.024465 -0.0114853
+ 2.051e+11Hz -0.0244709 -0.011469
+ 2.052e+11Hz -0.0244767 -0.0114528
+ 2.053e+11Hz -0.0244826 -0.0114366
+ 2.054e+11Hz -0.0244884 -0.0114205
+ 2.055e+11Hz -0.0244943 -0.0114045
+ 2.056e+11Hz -0.0245001 -0.0113886
+ 2.057e+11Hz -0.0245059 -0.0113727
+ 2.058e+11Hz -0.0245117 -0.0113569
+ 2.059e+11Hz -0.0245175 -0.0113412
+ 2.06e+11Hz -0.0245233 -0.0113256
+ 2.061e+11Hz -0.0245291 -0.0113101
+ 2.062e+11Hz -0.0245349 -0.0112946
+ 2.063e+11Hz -0.0245407 -0.0112792
+ 2.064e+11Hz -0.0245465 -0.0112639
+ 2.065e+11Hz -0.0245523 -0.0112487
+ 2.066e+11Hz -0.0245581 -0.0112335
+ 2.067e+11Hz -0.0245639 -0.0112184
+ 2.068e+11Hz -0.0245698 -0.0112034
+ 2.069e+11Hz -0.0245756 -0.0111885
+ 2.07e+11Hz -0.0245815 -0.0111737
+ 2.071e+11Hz -0.0245874 -0.0111589
+ 2.072e+11Hz -0.0245933 -0.0111442
+ 2.073e+11Hz -0.0245993 -0.0111296
+ 2.074e+11Hz -0.0246052 -0.0111151
+ 2.075e+11Hz -0.0246112 -0.0111006
+ 2.076e+11Hz -0.0246172 -0.0110862
+ 2.077e+11Hz -0.0246233 -0.0110719
+ 2.078e+11Hz -0.0246294 -0.0110577
+ 2.079e+11Hz -0.0246355 -0.0110435
+ 2.08e+11Hz -0.0246417 -0.0110294
+ 2.081e+11Hz -0.0246479 -0.0110154
+ 2.082e+11Hz -0.0246541 -0.0110014
+ 2.083e+11Hz -0.0246604 -0.0109876
+ 2.084e+11Hz -0.0246667 -0.0109738
+ 2.085e+11Hz -0.0246731 -0.01096
+ 2.086e+11Hz -0.0246795 -0.0109464
+ 2.087e+11Hz -0.024686 -0.0109328
+ 2.088e+11Hz -0.0246926 -0.0109192
+ 2.089e+11Hz -0.0246992 -0.0109058
+ 2.09e+11Hz -0.0247058 -0.0108923
+ 2.091e+11Hz -0.0247125 -0.010879
+ 2.092e+11Hz -0.0247193 -0.0108657
+ 2.093e+11Hz -0.0247262 -0.0108525
+ 2.094e+11Hz -0.0247331 -0.0108393
+ 2.095e+11Hz -0.0247401 -0.0108262
+ 2.096e+11Hz -0.0247471 -0.0108132
+ 2.097e+11Hz -0.0247543 -0.0108002
+ 2.098e+11Hz -0.0247615 -0.0107873
+ 2.099e+11Hz -0.0247688 -0.0107744
+ 2.1e+11Hz -0.0247761 -0.0107615
+ 2.101e+11Hz -0.0247836 -0.0107488
+ 2.102e+11Hz -0.0247911 -0.010736
+ 2.103e+11Hz -0.0247988 -0.0107233
+ 2.104e+11Hz -0.0248065 -0.0107107
+ 2.105e+11Hz -0.0248143 -0.0106981
+ 2.106e+11Hz -0.0248222 -0.0106855
+ 2.107e+11Hz -0.0248301 -0.010673
+ 2.108e+11Hz -0.0248382 -0.0106605
+ 2.109e+11Hz -0.0248464 -0.010648
+ 2.11e+11Hz -0.0248547 -0.0106356
+ 2.111e+11Hz -0.0248631 -0.0106232
+ 2.112e+11Hz -0.0248715 -0.0106109
+ 2.113e+11Hz -0.0248801 -0.0105985
+ 2.114e+11Hz -0.0248888 -0.0105862
+ 2.115e+11Hz -0.0248976 -0.0105739
+ 2.116e+11Hz -0.0249065 -0.0105616
+ 2.117e+11Hz -0.0249155 -0.0105494
+ 2.118e+11Hz -0.0249247 -0.0105372
+ 2.119e+11Hz -0.0249339 -0.0105249
+ 2.12e+11Hz -0.0249433 -0.0105127
+ 2.121e+11Hz -0.0249527 -0.0105005
+ 2.122e+11Hz -0.0249623 -0.0104883
+ 2.123e+11Hz -0.024972 -0.0104761
+ 2.124e+11Hz -0.0249819 -0.0104639
+ 2.125e+11Hz -0.0249918 -0.0104517
+ 2.126e+11Hz -0.0250019 -0.0104395
+ 2.127e+11Hz -0.0250121 -0.0104273
+ 2.128e+11Hz -0.0250225 -0.010415
+ 2.129e+11Hz -0.0250329 -0.0104028
+ 2.13e+11Hz -0.0250435 -0.0103905
+ 2.131e+11Hz -0.0250542 -0.0103783
+ 2.132e+11Hz -0.0250651 -0.010366
+ 2.133e+11Hz -0.025076 -0.0103536
+ 2.134e+11Hz -0.0250871 -0.0103413
+ 2.135e+11Hz -0.0250984 -0.0103289
+ 2.136e+11Hz -0.0251098 -0.0103165
+ 2.137e+11Hz -0.0251213 -0.010304
+ 2.138e+11Hz -0.0251329 -0.0102915
+ 2.139e+11Hz -0.0251447 -0.010279
+ 2.14e+11Hz -0.0251566 -0.0102664
+ 2.141e+11Hz -0.0251687 -0.0102538
+ 2.142e+11Hz -0.0251808 -0.0102411
+ 2.143e+11Hz -0.0251932 -0.0102283
+ 2.144e+11Hz -0.0252056 -0.0102155
+ 2.145e+11Hz -0.0252182 -0.0102026
+ 2.146e+11Hz -0.025231 -0.0101897
+ 2.147e+11Hz -0.0252438 -0.0101767
+ 2.148e+11Hz -0.0252569 -0.0101636
+ 2.149e+11Hz -0.02527 -0.0101504
+ 2.15e+11Hz -0.0252833 -0.0101372
+ 2.151e+11Hz -0.0252967 -0.0101239
+ 2.152e+11Hz -0.0253103 -0.0101105
+ 2.153e+11Hz -0.025324 -0.010097
+ 2.154e+11Hz -0.0253378 -0.0100834
+ 2.155e+11Hz -0.0253518 -0.0100697
+ 2.156e+11Hz -0.0253659 -0.0100559
+ 2.157e+11Hz -0.0253802 -0.010042
+ 2.158e+11Hz -0.0253946 -0.010028
+ 2.159e+11Hz -0.0254091 -0.0100139
+ 2.16e+11Hz -0.0254238 -0.00999965
+ 2.161e+11Hz -0.0254385 -0.0099853
+ 2.162e+11Hz -0.0254535 -0.00997083
+ 2.163e+11Hz -0.0254685 -0.00995624
+ 2.164e+11Hz -0.0254837 -0.00994151
+ 2.165e+11Hz -0.025499 -0.00992666
+ 2.166e+11Hz -0.0255145 -0.00991166
+ 2.167e+11Hz -0.02553 -0.00989653
+ 2.168e+11Hz -0.0255457 -0.00988125
+ 2.169e+11Hz -0.0255615 -0.00986583
+ 2.17e+11Hz -0.0255775 -0.00985026
+ 2.171e+11Hz -0.0255935 -0.00983453
+ 2.172e+11Hz -0.0256097 -0.00981864
+ 2.173e+11Hz -0.025626 -0.0098026
+ 2.174e+11Hz -0.0256424 -0.00978639
+ 2.175e+11Hz -0.025659 -0.00977001
+ 2.176e+11Hz -0.0256756 -0.00975347
+ 2.177e+11Hz -0.0256924 -0.00973675
+ 2.178e+11Hz -0.0257093 -0.00971985
+ 2.179e+11Hz -0.0257262 -0.00970276
+ 2.18e+11Hz -0.0257433 -0.0096855
+ 2.181e+11Hz -0.0257605 -0.00966805
+ 2.182e+11Hz -0.0257778 -0.0096504
+ 2.183e+11Hz -0.0257952 -0.00963256
+ 2.184e+11Hz -0.0258126 -0.00961452
+ 2.185e+11Hz -0.0258302 -0.00959629
+ 2.186e+11Hz -0.0258479 -0.00957785
+ 2.187e+11Hz -0.0258656 -0.0095592
+ 2.188e+11Hz -0.0258834 -0.00954034
+ 2.189e+11Hz -0.0259014 -0.00952126
+ 2.19e+11Hz -0.0259194 -0.00950197
+ 2.191e+11Hz -0.0259374 -0.00948247
+ 2.192e+11Hz -0.0259556 -0.00946273
+ 2.193e+11Hz -0.0259738 -0.00944278
+ 2.194e+11Hz -0.0259921 -0.00942259
+ 2.195e+11Hz -0.0260104 -0.00940218
+ 2.196e+11Hz -0.0260288 -0.00938153
+ 2.197e+11Hz -0.0260473 -0.00936064
+ 2.198e+11Hz -0.0260658 -0.00933951
+ 2.199e+11Hz -0.0260844 -0.00931815
+ 2.2e+11Hz -0.026103 -0.00929654
+ 2.201e+11Hz -0.0261217 -0.00927468
+ 2.202e+11Hz -0.0261404 -0.00925257
+ 2.203e+11Hz -0.0261591 -0.00923021
+ 2.204e+11Hz -0.0261779 -0.00920759
+ 2.205e+11Hz -0.0261967 -0.00918472
+ 2.206e+11Hz -0.0262156 -0.00916159
+ 2.207e+11Hz -0.0262344 -0.0091382
+ 2.208e+11Hz -0.0262533 -0.00911455
+ 2.209e+11Hz -0.0262722 -0.00909063
+ 2.21e+11Hz -0.0262911 -0.00906644
+ 2.211e+11Hz -0.0263099 -0.00904199
+ 2.212e+11Hz -0.0263288 -0.00901726
+ 2.213e+11Hz -0.0263477 -0.00899226
+ 2.214e+11Hz -0.0263666 -0.00896699
+ 2.215e+11Hz -0.0263855 -0.00894144
+ 2.216e+11Hz -0.0264044 -0.00891561
+ 2.217e+11Hz -0.0264232 -0.00888951
+ 2.218e+11Hz -0.026442 -0.00886312
+ 2.219e+11Hz -0.0264608 -0.00883645
+ 2.22e+11Hz -0.0264796 -0.0088095
+ 2.221e+11Hz -0.0264983 -0.00878227
+ 2.222e+11Hz -0.0265169 -0.00875475
+ 2.223e+11Hz -0.0265356 -0.00872694
+ 2.224e+11Hz -0.0265541 -0.00869884
+ 2.225e+11Hz -0.0265727 -0.00867046
+ 2.226e+11Hz -0.0265911 -0.00864179
+ 2.227e+11Hz -0.0266095 -0.00861283
+ 2.228e+11Hz -0.0266278 -0.00858358
+ 2.229e+11Hz -0.026646 -0.00855404
+ 2.23e+11Hz -0.0266642 -0.0085242
+ 2.231e+11Hz -0.0266823 -0.00849408
+ 2.232e+11Hz -0.0267003 -0.00846366
+ 2.233e+11Hz -0.0267181 -0.00843296
+ 2.234e+11Hz -0.0267359 -0.00840196
+ 2.235e+11Hz -0.0267536 -0.00837066
+ 2.236e+11Hz -0.0267712 -0.00833908
+ 2.237e+11Hz -0.0267886 -0.0083072
+ 2.238e+11Hz -0.026806 -0.00827504
+ 2.239e+11Hz -0.0268232 -0.00824258
+ 2.24e+11Hz -0.0268402 -0.00820983
+ 2.241e+11Hz -0.0268572 -0.00817679
+ 2.242e+11Hz -0.026874 -0.00814346
+ 2.243e+11Hz -0.0268906 -0.00810984
+ 2.244e+11Hz -0.0269071 -0.00807593
+ 2.245e+11Hz -0.0269235 -0.00804174
+ 2.246e+11Hz -0.0269397 -0.00800726
+ 2.247e+11Hz -0.0269557 -0.0079725
+ 2.248e+11Hz -0.0269716 -0.00793745
+ 2.249e+11Hz -0.0269872 -0.00790212
+ 2.25e+11Hz -0.0270027 -0.00786651
+ 2.251e+11Hz -0.027018 -0.00783062
+ 2.252e+11Hz -0.0270332 -0.00779445
+ 2.253e+11Hz -0.0270481 -0.007758
+ 2.254e+11Hz -0.0270628 -0.00772128
+ 2.255e+11Hz -0.0270773 -0.00768429
+ 2.256e+11Hz -0.0270917 -0.00764702
+ 2.257e+11Hz -0.0271058 -0.00760949
+ 2.258e+11Hz -0.0271196 -0.00757169
+ 2.259e+11Hz -0.0271333 -0.00753363
+ 2.26e+11Hz -0.0271467 -0.0074953
+ 2.261e+11Hz -0.0271599 -0.00745671
+ 2.262e+11Hz -0.0271729 -0.00741787
+ 2.263e+11Hz -0.0271856 -0.00737877
+ 2.264e+11Hz -0.0271981 -0.00733942
+ 2.265e+11Hz -0.0272103 -0.00729982
+ 2.266e+11Hz -0.0272222 -0.00725997
+ 2.267e+11Hz -0.0272339 -0.00721988
+ 2.268e+11Hz -0.0272453 -0.00717955
+ 2.269e+11Hz -0.0272565 -0.00713898
+ 2.27e+11Hz -0.0272674 -0.00709817
+ 2.271e+11Hz -0.027278 -0.00705714
+ 2.272e+11Hz -0.0272883 -0.00701587
+ 2.273e+11Hz -0.0272984 -0.00697438
+ 2.274e+11Hz -0.0273081 -0.00693267
+ 2.275e+11Hz -0.0273176 -0.00689075
+ 2.276e+11Hz -0.0273267 -0.00684861
+ 2.277e+11Hz -0.0273356 -0.00680626
+ 2.278e+11Hz -0.0273441 -0.0067637
+ 2.279e+11Hz -0.0273523 -0.00672094
+ 2.28e+11Hz -0.0273602 -0.00667798
+ 2.281e+11Hz -0.0273678 -0.00663483
+ 2.282e+11Hz -0.0273751 -0.00659148
+ 2.283e+11Hz -0.0273821 -0.00654795
+ 2.284e+11Hz -0.0273887 -0.00650424
+ 2.285e+11Hz -0.027395 -0.00646035
+ 2.286e+11Hz -0.0274009 -0.00641629
+ 2.287e+11Hz -0.0274065 -0.00637206
+ 2.288e+11Hz -0.0274118 -0.00632767
+ 2.289e+11Hz -0.0274167 -0.00628311
+ 2.29e+11Hz -0.0274213 -0.0062384
+ 2.291e+11Hz -0.0274255 -0.00619354
+ 2.292e+11Hz -0.0274294 -0.00614853
+ 2.293e+11Hz -0.0274329 -0.00610338
+ 2.294e+11Hz -0.0274361 -0.0060581
+ 2.295e+11Hz -0.0274388 -0.00601268
+ 2.296e+11Hz -0.0274413 -0.00596714
+ 2.297e+11Hz -0.0274433 -0.00592148
+ 2.298e+11Hz -0.027445 -0.0058757
+ 2.299e+11Hz -0.0274463 -0.00582981
+ 2.3e+11Hz -0.0274472 -0.00578382
+ 2.301e+11Hz -0.0274478 -0.00573772
+ 2.302e+11Hz -0.027448 -0.00569153
+ 2.303e+11Hz -0.0274478 -0.00564524
+ 2.304e+11Hz -0.0274472 -0.00559888
+ 2.305e+11Hz -0.0274462 -0.00555243
+ 2.306e+11Hz -0.0274449 -0.00550591
+ 2.307e+11Hz -0.0274431 -0.00545932
+ 2.308e+11Hz -0.027441 -0.00541266
+ 2.309e+11Hz -0.0274384 -0.00536595
+ 2.31e+11Hz -0.0274355 -0.00531919
+ 2.311e+11Hz -0.0274322 -0.00527237
+ 2.312e+11Hz -0.0274285 -0.00522552
+ 2.313e+11Hz -0.0274244 -0.00517863
+ 2.314e+11Hz -0.0274199 -0.00513171
+ 2.315e+11Hz -0.027415 -0.00508477
+ 2.316e+11Hz -0.0274097 -0.00503781
+ 2.317e+11Hz -0.027404 -0.00499083
+ 2.318e+11Hz -0.0273979 -0.00494384
+ 2.319e+11Hz -0.0273914 -0.00489686
+ 2.32e+11Hz -0.0273845 -0.00484988
+ 2.321e+11Hz -0.0273773 -0.0048029
+ 2.322e+11Hz -0.0273696 -0.00475594
+ 2.323e+11Hz -0.0273615 -0.004709
+ 2.324e+11Hz -0.027353 -0.00466209
+ 2.325e+11Hz -0.0273441 -0.00461521
+ 2.326e+11Hz -0.0273348 -0.00456836
+ 2.327e+11Hz -0.0273251 -0.00452156
+ 2.328e+11Hz -0.027315 -0.00447481
+ 2.329e+11Hz -0.0273045 -0.00442811
+ 2.33e+11Hz -0.0272936 -0.00438147
+ 2.331e+11Hz -0.0272824 -0.0043349
+ 2.332e+11Hz -0.0272707 -0.0042884
+ 2.333e+11Hz -0.0272586 -0.00424197
+ 2.334e+11Hz -0.0272461 -0.00419563
+ 2.335e+11Hz -0.0272333 -0.00414937
+ 2.336e+11Hz -0.02722 -0.00410321
+ 2.337e+11Hz -0.0272064 -0.00405715
+ 2.338e+11Hz -0.0271923 -0.00401119
+ 2.339e+11Hz -0.0271779 -0.00396534
+ 2.34e+11Hz -0.0271631 -0.0039196
+ 2.341e+11Hz -0.0271479 -0.00387399
+ 2.342e+11Hz -0.0271324 -0.0038285
+ 2.343e+11Hz -0.0271164 -0.00378314
+ 2.344e+11Hz -0.0271001 -0.00373791
+ 2.345e+11Hz -0.0270834 -0.00369283
+ 2.346e+11Hz -0.0270663 -0.00364789
+ 2.347e+11Hz -0.0270489 -0.00360311
+ 2.348e+11Hz -0.027031 -0.00355848
+ 2.349e+11Hz -0.0270129 -0.00351401
+ 2.35e+11Hz -0.0269943 -0.00346971
+ 2.351e+11Hz -0.0269754 -0.00342559
+ 2.352e+11Hz -0.0269561 -0.00338163
+ 2.353e+11Hz -0.0269365 -0.00333786
+ 2.354e+11Hz -0.0269165 -0.00329428
+ 2.355e+11Hz -0.0268962 -0.00325088
+ 2.356e+11Hz -0.0268755 -0.00320768
+ 2.357e+11Hz -0.0268545 -0.00316468
+ 2.358e+11Hz -0.0268331 -0.00312188
+ 2.359e+11Hz -0.0268114 -0.0030793
+ 2.36e+11Hz -0.0267894 -0.00303692
+ 2.361e+11Hz -0.026767 -0.00299476
+ 2.362e+11Hz -0.0267443 -0.00295283
+ 2.363e+11Hz -0.0267213 -0.00291112
+ 2.364e+11Hz -0.026698 -0.00286964
+ 2.365e+11Hz -0.0266743 -0.00282839
+ 2.366e+11Hz -0.0266503 -0.00278739
+ 2.367e+11Hz -0.0266261 -0.00274662
+ 2.368e+11Hz -0.0266015 -0.0027061
+ 2.369e+11Hz -0.0265766 -0.00266583
+ 2.37e+11Hz -0.0265514 -0.00262581
+ 2.371e+11Hz -0.0265259 -0.00258605
+ 2.372e+11Hz -0.0265002 -0.00254655
+ 2.373e+11Hz -0.0264741 -0.00250732
+ 2.374e+11Hz -0.0264478 -0.00246835
+ 2.375e+11Hz -0.0264212 -0.00242965
+ 2.376e+11Hz -0.0263943 -0.00239123
+ 2.377e+11Hz -0.0263671 -0.00235308
+ 2.378e+11Hz -0.0263397 -0.00231521
+ 2.379e+11Hz -0.026312 -0.00227762
+ 2.38e+11Hz -0.0262841 -0.00224033
+ 2.381e+11Hz -0.0262559 -0.00220331
+ 2.382e+11Hz -0.0262275 -0.00216659
+ 2.383e+11Hz -0.0261988 -0.00213017
+ 2.384e+11Hz -0.0261699 -0.00209404
+ 2.385e+11Hz -0.0261408 -0.00205821
+ 2.386e+11Hz -0.0261114 -0.00202268
+ 2.387e+11Hz -0.0260818 -0.00198746
+ 2.388e+11Hz -0.026052 -0.00195254
+ 2.389e+11Hz -0.0260219 -0.00191792
+ 2.39e+11Hz -0.0259917 -0.00188362
+ 2.391e+11Hz -0.0259613 -0.00184963
+ 2.392e+11Hz -0.0259306 -0.00181595
+ 2.393e+11Hz -0.0258998 -0.00178259
+ 2.394e+11Hz -0.0258687 -0.00174955
+ 2.395e+11Hz -0.0258375 -0.00171682
+ 2.396e+11Hz -0.0258061 -0.00168442
+ 2.397e+11Hz -0.0257746 -0.00165234
+ 2.398e+11Hz -0.0257428 -0.00162058
+ 2.399e+11Hz -0.0257109 -0.00158914
+ 2.4e+11Hz -0.0256788 -0.00155803
+ 2.401e+11Hz -0.0256466 -0.00152724
+ 2.402e+11Hz -0.0256142 -0.00149679
+ 2.403e+11Hz -0.0255817 -0.00146666
+ 2.404e+11Hz -0.025549 -0.00143686
+ 2.405e+11Hz -0.0255162 -0.00140739
+ 2.406e+11Hz -0.0254833 -0.00137825
+ 2.407e+11Hz -0.0254502 -0.00134944
+ 2.408e+11Hz -0.025417 -0.00132096
+ 2.409e+11Hz -0.0253837 -0.00129281
+ 2.41e+11Hz -0.0253503 -0.001265
+ 2.411e+11Hz -0.0253168 -0.00123752
+ 2.412e+11Hz -0.0252831 -0.00121037
+ 2.413e+11Hz -0.0252494 -0.00118355
+ 2.414e+11Hz -0.0252156 -0.00115707
+ 2.415e+11Hz -0.0251817 -0.00113092
+ 2.416e+11Hz -0.0251477 -0.0011051
+ 2.417e+11Hz -0.0251136 -0.00107961
+ 2.418e+11Hz -0.0250794 -0.00105445
+ 2.419e+11Hz -0.0250452 -0.00102962
+ 2.42e+11Hz -0.0250109 -0.00100513
+ 2.421e+11Hz -0.0249766 -0.000980965
+ 2.422e+11Hz -0.0249422 -0.000957129
+ 2.423e+11Hz -0.0249077 -0.000933622
+ 2.424e+11Hz -0.0248732 -0.000910443
+ 2.425e+11Hz -0.0248386 -0.00088759
+ 2.426e+11Hz -0.024804 -0.000865064
+ 2.427e+11Hz -0.0247694 -0.000842863
+ 2.428e+11Hz -0.0247347 -0.000820986
+ 2.429e+11Hz -0.0247001 -0.000799432
+ 2.43e+11Hz -0.0246653 -0.000778199
+ 2.431e+11Hz -0.0246306 -0.000757287
+ 2.432e+11Hz -0.0245959 -0.000736694
+ 2.433e+11Hz -0.0245611 -0.000716418
+ 2.434e+11Hz -0.0245264 -0.000696459
+ 2.435e+11Hz -0.0244916 -0.000676815
+ 2.436e+11Hz -0.0244568 -0.000657484
+ 2.437e+11Hz -0.0244221 -0.000638464
+ 2.438e+11Hz -0.0243873 -0.000619755
+ 2.439e+11Hz -0.0243526 -0.000601353
+ 2.44e+11Hz -0.0243179 -0.000583258
+ 2.441e+11Hz -0.0242832 -0.000565468
+ 2.442e+11Hz -0.0242485 -0.000547981
+ 2.443e+11Hz -0.0242139 -0.000530794
+ 2.444e+11Hz -0.0241793 -0.000513906
+ 2.445e+11Hz -0.0241447 -0.000497316
+ 2.446e+11Hz -0.0241101 -0.00048102
+ 2.447e+11Hz -0.0240756 -0.000465017
+ 2.448e+11Hz -0.0240412 -0.000449304
+ 2.449e+11Hz -0.0240068 -0.00043388
+ 2.45e+11Hz -0.0239724 -0.000418742
+ 2.451e+11Hz -0.0239381 -0.000403888
+ 2.452e+11Hz -0.0239039 -0.000389316
+ 2.453e+11Hz -0.0238697 -0.000375023
+ 2.454e+11Hz -0.0238356 -0.000361008
+ 2.455e+11Hz -0.0238015 -0.000347267
+ 2.456e+11Hz -0.0237676 -0.000333798
+ 2.457e+11Hz -0.0237337 -0.0003206
+ 2.458e+11Hz -0.0236998 -0.000307669
+ 2.459e+11Hz -0.0236661 -0.000295002
+ 2.46e+11Hz -0.0236324 -0.000282599
+ 2.461e+11Hz -0.0235988 -0.000270455
+ 2.462e+11Hz -0.0235653 -0.000258569
+ 2.463e+11Hz -0.0235319 -0.000246937
+ 2.464e+11Hz -0.0234985 -0.000235558
+ 2.465e+11Hz -0.0234653 -0.000224429
+ 2.466e+11Hz -0.0234321 -0.000213547
+ 2.467e+11Hz -0.0233991 -0.000202909
+ 2.468e+11Hz -0.0233662 -0.000192513
+ 2.469e+11Hz -0.0233333 -0.000182357
+ 2.47e+11Hz -0.0233006 -0.000172437
+ 2.471e+11Hz -0.0232679 -0.000162751
+ 2.472e+11Hz -0.0232354 -0.000153296
+ 2.473e+11Hz -0.023203 -0.00014407
+ 2.474e+11Hz -0.0231706 -0.00013507
+ 2.475e+11Hz -0.0231384 -0.000126293
+ 2.476e+11Hz -0.0231063 -0.000117737
+ 2.477e+11Hz -0.0230744 -0.000109399
+ 2.478e+11Hz -0.0230425 -0.000101277
+ 2.479e+11Hz -0.0230108 -9.33669e-05
+ 2.48e+11Hz -0.0229792 -8.5667e-05
+ 2.481e+11Hz -0.0229477 -7.81745e-05
+ 2.482e+11Hz -0.0229163 -7.08868e-05
+ 2.483e+11Hz -0.022885 -6.38012e-05
+ 2.484e+11Hz -0.0228539 -5.6915e-05
+ 2.485e+11Hz -0.0228229 -5.02257e-05
+ 2.486e+11Hz -0.0227921 -4.37307e-05
+ 2.487e+11Hz -0.0227613 -3.74273e-05
+ 2.488e+11Hz -0.0227307 -3.13131e-05
+ 2.489e+11Hz -0.0227002 -2.53853e-05
+ 2.49e+11Hz -0.0226699 -1.96415e-05
+ 2.491e+11Hz -0.0226397 -1.4079e-05
+ 2.492e+11Hz -0.0226096 -8.69551e-06
+ 2.493e+11Hz -0.0225796 -3.48836e-06
+ 2.494e+11Hz -0.0225498 1.5449e-06
+ 2.495e+11Hz -0.0225202 6.40676e-06
+ 2.496e+11Hz -0.0224906 1.10997e-05
+ 2.497e+11Hz -0.0224612 1.5626e-05
+ 2.498e+11Hz -0.022432 1.99883e-05
+ 2.499e+11Hz -0.0224029 2.41889e-05
+ 2.5e+11Hz -0.0223739 2.82301e-05
+ 2.501e+11Hz -0.022345 3.21144e-05
+ 2.502e+11Hz -0.0223163 3.5844e-05
+ 2.503e+11Hz -0.0222878 3.94213e-05
+ 2.504e+11Hz -0.0222594 4.28485e-05
+ 2.505e+11Hz -0.0222311 4.61279e-05
+ 2.506e+11Hz -0.022203 4.92618e-05
+ 2.507e+11Hz -0.022175 5.22523e-05
+ 2.508e+11Hz -0.0221471 5.51017e-05
+ 2.509e+11Hz -0.0221194 5.78121e-05
+ 2.51e+11Hz -0.0220919 6.03856e-05
+ 2.511e+11Hz -0.0220645 6.28245e-05
+ 2.512e+11Hz -0.0220372 6.51306e-05
+ 2.513e+11Hz -0.0220101 6.73063e-05
+ 2.514e+11Hz -0.0219831 6.93533e-05
+ 2.515e+11Hz -0.0219563 7.12739e-05
+ 2.516e+11Hz -0.0219296 7.307e-05
+ 2.517e+11Hz -0.0219031 7.47435e-05
+ 2.518e+11Hz -0.0218767 7.62963e-05
+ 2.519e+11Hz -0.0218505 7.77305e-05
+ 2.52e+11Hz -0.0218244 7.90478e-05
+ 2.521e+11Hz -0.0217984 8.02503e-05
+ 2.522e+11Hz -0.0217726 8.13396e-05
+ 2.523e+11Hz -0.021747 8.23176e-05
+ 2.524e+11Hz -0.0217215 8.31861e-05
+ 2.525e+11Hz -0.0216961 8.39469e-05
+ 2.526e+11Hz -0.0216709 8.46017e-05
+ 2.527e+11Hz -0.0216458 8.51522e-05
+ 2.528e+11Hz -0.0216209 8.56002e-05
+ 2.529e+11Hz -0.0215961 8.59473e-05
+ 2.53e+11Hz -0.0215715 8.61952e-05
+ 2.531e+11Hz -0.021547 8.63456e-05
+ 2.532e+11Hz -0.0215227 8.63999e-05
+ 2.533e+11Hz -0.0214985 8.63598e-05
+ 2.534e+11Hz -0.0214745 8.6227e-05
+ 2.535e+11Hz -0.0214506 8.60029e-05
+ 2.536e+11Hz -0.0214269 8.56891e-05
+ 2.537e+11Hz -0.0214033 8.52871e-05
+ 2.538e+11Hz -0.0213798 8.47985e-05
+ 2.539e+11Hz -0.0213565 8.42246e-05
+ 2.54e+11Hz -0.0213334 8.3567e-05
+ 2.541e+11Hz -0.0213104 8.28271e-05
+ 2.542e+11Hz -0.0212875 8.20064e-05
+ 2.543e+11Hz -0.0212648 8.11063e-05
+ 2.544e+11Hz -0.0212423 8.01282e-05
+ 2.545e+11Hz -0.0212199 7.90735e-05
+ 2.546e+11Hz -0.0211976 7.79437e-05
+ 2.547e+11Hz -0.0211755 7.674e-05
+ 2.548e+11Hz -0.0211536 7.54639e-05
+ 2.549e+11Hz -0.0211318 7.41168e-05
+ 2.55e+11Hz -0.0211101 7.26999e-05
+ 2.551e+11Hz -0.0210886 7.12146e-05
+ 2.552e+11Hz -0.0210673 6.96624e-05
+ 2.553e+11Hz -0.0210461 6.80445e-05
+ 2.554e+11Hz -0.021025 6.63622e-05
+ 2.555e+11Hz -0.0210041 6.4617e-05
+ 2.556e+11Hz -0.0209833 6.28101e-05
+ 2.557e+11Hz -0.0209627 6.09428e-05
+ 2.558e+11Hz -0.0209423 5.90166e-05
+ 2.559e+11Hz -0.020922 5.70326e-05
+ 2.56e+11Hz -0.0209018 5.49924e-05
+ 2.561e+11Hz -0.0208818 5.28972e-05
+ 2.562e+11Hz -0.020862 5.07483e-05
+ 2.563e+11Hz -0.0208423 4.85471e-05
+ 2.564e+11Hz -0.0208228 4.62949e-05
+ 2.565e+11Hz -0.0208034 4.39932e-05
+ 2.566e+11Hz -0.0207841 4.16432e-05
+ 2.567e+11Hz -0.0207651 3.92464e-05
+ 2.568e+11Hz -0.0207461 3.68041e-05
+ 2.569e+11Hz -0.0207274 3.43178e-05
+ 2.57e+11Hz -0.0207088 3.17889e-05
+ 2.571e+11Hz -0.0206903 2.92187e-05
+ 2.572e+11Hz -0.020672 2.66087e-05
+ 2.573e+11Hz -0.0206538 2.39604e-05
+ 2.574e+11Hz -0.0206359 2.12753e-05
+ 2.575e+11Hz -0.020618 1.85547e-05
+ 2.576e+11Hz -0.0206004 1.58003e-05
+ 2.577e+11Hz -0.0205828 1.30135e-05
+ 2.578e+11Hz -0.0205655 1.0196e-05
+ 2.579e+11Hz -0.0205483 7.34912e-06
+ 2.58e+11Hz -0.0205312 4.47462e-06
+ 2.581e+11Hz -0.0205144 1.57405e-06
+ 2.582e+11Hz -0.0204976 -1.35096e-06
+ 2.583e+11Hz -0.0204811 -4.29876e-06
+ 2.584e+11Hz -0.0204647 -7.26767e-06
+ 2.585e+11Hz -0.0204485 -1.0256e-05
+ 2.586e+11Hz -0.0204324 -1.3262e-05
+ 2.587e+11Hz -0.0204165 -1.6284e-05
+ 2.588e+11Hz -0.0204007 -1.93201e-05
+ 2.589e+11Hz -0.0203852 -2.23686e-05
+ 2.59e+11Hz -0.0203697 -2.54275e-05
+ 2.591e+11Hz -0.0203545 -2.84952e-05
+ 2.592e+11Hz -0.0203394 -3.15696e-05
+ 2.593e+11Hz -0.0203245 -3.46488e-05
+ 2.594e+11Hz -0.0203097 -3.77309e-05
+ 2.595e+11Hz -0.0202951 -4.08139e-05
+ 2.596e+11Hz -0.0202807 -4.38958e-05
+ 2.597e+11Hz -0.0202665 -4.69745e-05
+ 2.598e+11Hz -0.0202524 -5.00479e-05
+ 2.599e+11Hz -0.0202385 -5.3114e-05
+ 2.6e+11Hz -0.0202247 -5.61705e-05
+ 2.601e+11Hz -0.0202112 -5.92153e-05
+ 2.602e+11Hz -0.0201977 -6.22462e-05
+ 2.603e+11Hz -0.0201845 -6.5261e-05
+ 2.604e+11Hz -0.0201714 -6.82573e-05
+ 2.605e+11Hz -0.0201585 -7.12328e-05
+ 2.606e+11Hz -0.0201458 -7.41852e-05
+ 2.607e+11Hz -0.0201333 -7.71121e-05
+ 2.608e+11Hz -0.0201209 -8.00111e-05
+ 2.609e+11Hz -0.0201087 -8.28796e-05
+ 2.61e+11Hz -0.0200966 -8.57153e-05
+ 2.611e+11Hz -0.0200848 -8.85157e-05
+ 2.612e+11Hz -0.0200731 -9.1278e-05
+ 2.613e+11Hz -0.0200616 -9.39998e-05
+ 2.614e+11Hz -0.0200502 -9.66785e-05
+ 2.615e+11Hz -0.020039 -9.93113e-05
+ 2.616e+11Hz -0.020028 -0.000101896
+ 2.617e+11Hz -0.0200172 -0.000104429
+ 2.618e+11Hz -0.0200065 -0.000106908
+ 2.619e+11Hz -0.019996 -0.00010933
+ 2.62e+11Hz -0.0199857 -0.000111693
+ 2.621e+11Hz -0.0199756 -0.000113993
+ 2.622e+11Hz -0.0199656 -0.000116228
+ 2.623e+11Hz -0.0199558 -0.000118394
+ 2.624e+11Hz -0.0199462 -0.00012049
+ 2.625e+11Hz -0.0199367 -0.000122511
+ 2.626e+11Hz -0.0199274 -0.000124455
+ 2.627e+11Hz -0.0199183 -0.000126319
+ 2.628e+11Hz -0.0199094 -0.0001281
+ 2.629e+11Hz -0.0199006 -0.000129794
+ 2.63e+11Hz -0.019892 -0.000131399
+ 2.631e+11Hz -0.0198835 -0.000132912
+ 2.632e+11Hz -0.0198753 -0.000134329
+ 2.633e+11Hz -0.0198672 -0.000135647
+ 2.634e+11Hz -0.0198592 -0.000136863
+ 2.635e+11Hz -0.0198514 -0.000137973
+ 2.636e+11Hz -0.0198438 -0.000138976
+ 2.637e+11Hz -0.0198364 -0.000139866
+ 2.638e+11Hz -0.0198291 -0.000140642
+ 2.639e+11Hz -0.0198219 -0.0001413
+ 2.64e+11Hz -0.0198149 -0.000141836
+ 2.641e+11Hz -0.0198081 -0.000142247
+ 2.642e+11Hz -0.0198015 -0.00014253
+ 2.643e+11Hz -0.019795 -0.000142682
+ 2.644e+11Hz -0.0197886 -0.000142699
+ 2.645e+11Hz -0.0197824 -0.000142578
+ 2.646e+11Hz -0.0197764 -0.000142315
+ 2.647e+11Hz -0.0197705 -0.000141908
+ 2.648e+11Hz -0.0197647 -0.000141353
+ 2.649e+11Hz -0.0197591 -0.000140646
+ 2.65e+11Hz -0.0197536 -0.000139785
+ 2.651e+11Hz -0.0197483 -0.000138766
+ 2.652e+11Hz -0.0197431 -0.000137585
+ 2.653e+11Hz -0.0197381 -0.00013624
+ 2.654e+11Hz -0.0197332 -0.000134726
+ 2.655e+11Hz -0.0197284 -0.000133042
+ 2.656e+11Hz -0.0197237 -0.000131182
+ 2.657e+11Hz -0.0197192 -0.000129145
+ 2.658e+11Hz -0.0197148 -0.000126927
+ 2.659e+11Hz -0.0197105 -0.000124524
+ 2.66e+11Hz -0.0197064 -0.000121934
+ 2.661e+11Hz -0.0197023 -0.000119153
+ 2.662e+11Hz -0.0196984 -0.000116178
+ 2.663e+11Hz -0.0196946 -0.000113006
+ 2.664e+11Hz -0.0196909 -0.000109633
+ 2.665e+11Hz -0.0196873 -0.000106058
+ 2.666e+11Hz -0.0196838 -0.000102276
+ 2.667e+11Hz -0.0196804 -9.82843e-05
+ 2.668e+11Hz -0.0196771 -9.40805e-05
+ 2.669e+11Hz -0.0196739 -8.96614e-05
+ 2.67e+11Hz -0.0196708 -8.5024e-05
+ 2.671e+11Hz -0.0196678 -8.01655e-05
+ 2.672e+11Hz -0.0196648 -7.5083e-05
+ 2.673e+11Hz -0.019662 -6.97738e-05
+ 2.674e+11Hz -0.0196592 -6.42351e-05
+ 2.675e+11Hz -0.0196564 -5.84643e-05
+ 2.676e+11Hz -0.0196538 -5.24586e-05
+ 2.677e+11Hz -0.0196512 -4.62156e-05
+ 2.678e+11Hz -0.0196486 -3.97327e-05
+ 2.679e+11Hz -0.0196462 -3.30074e-05
+ 2.68e+11Hz -0.0196437 -2.60373e-05
+ 2.681e+11Hz -0.0196413 -1.88202e-05
+ 2.682e+11Hz -0.019639 -1.13536e-05
+ 2.683e+11Hz -0.0196367 -3.63541e-06
+ 2.684e+11Hz -0.0196344 4.33653e-06
+ 2.685e+11Hz -0.0196322 1.25643e-05
+ 2.686e+11Hz -0.01963 2.10499e-05
+ 2.687e+11Hz -0.0196278 2.97953e-05
+ 2.688e+11Hz -0.0196256 3.88023e-05
+ 2.689e+11Hz -0.0196234 4.80727e-05
+ 2.69e+11Hz -0.0196212 5.76082e-05
+ 2.691e+11Hz -0.0196191 6.74105e-05
+ 2.692e+11Hz -0.0196169 7.74809e-05
+ 2.693e+11Hz -0.0196147 8.78211e-05
+ 2.694e+11Hz -0.0196125 9.84323e-05
+ 2.695e+11Hz -0.0196103 0.000109316
+ 2.696e+11Hz -0.019608 0.000120473
+ 2.697e+11Hz -0.0196058 0.000131905
+ 2.698e+11Hz -0.0196035 0.000143612
+ 2.699e+11Hz -0.0196011 0.000155596
+ 2.7e+11Hz -0.0195987 0.000167857
+ 2.701e+11Hz -0.0195962 0.000180396
+ 2.702e+11Hz -0.0195937 0.000193214
+ 2.703e+11Hz -0.0195912 0.00020631
+ 2.704e+11Hz -0.0195885 0.000219687
+ 2.705e+11Hz -0.0195858 0.000233343
+ 2.706e+11Hz -0.019583 0.000247279
+ 2.707e+11Hz -0.0195801 0.000261495
+ 2.708e+11Hz -0.0195771 0.000275991
+ 2.709e+11Hz -0.0195741 0.000290768
+ 2.71e+11Hz -0.0195709 0.000305823
+ 2.711e+11Hz -0.0195676 0.000321159
+ 2.712e+11Hz -0.0195642 0.000336773
+ 2.713e+11Hz -0.0195607 0.000352665
+ 2.714e+11Hz -0.019557 0.000368835
+ 2.715e+11Hz -0.0195532 0.000385281
+ 2.716e+11Hz -0.0195493 0.000402004
+ 2.717e+11Hz -0.0195453 0.000419001
+ 2.718e+11Hz -0.019541 0.000436272
+ 2.719e+11Hz -0.0195367 0.000453815
+ 2.72e+11Hz -0.0195321 0.000471629
+ 2.721e+11Hz -0.0195274 0.000489712
+ 2.722e+11Hz -0.0195226 0.000508063
+ 2.723e+11Hz -0.0195175 0.00052668
+ 2.724e+11Hz -0.0195123 0.000545561
+ 2.725e+11Hz -0.0195069 0.000564704
+ 2.726e+11Hz -0.0195012 0.000584106
+ 2.727e+11Hz -0.0194954 0.000603767
+ 2.728e+11Hz -0.0194894 0.000623682
+ 2.729e+11Hz -0.0194831 0.000643851
+ 2.73e+11Hz -0.0194766 0.000664269
+ 2.731e+11Hz -0.0194699 0.000684935
+ 2.732e+11Hz -0.019463 0.000705845
+ 2.733e+11Hz -0.0194558 0.000726996
+ 2.734e+11Hz -0.0194484 0.000748386
+ 2.735e+11Hz -0.0194408 0.000770011
+ 2.736e+11Hz -0.0194329 0.000791868
+ 2.737e+11Hz -0.0194247 0.000813953
+ 2.738e+11Hz -0.0194162 0.000836262
+ 2.739e+11Hz -0.0194075 0.000858792
+ 2.74e+11Hz -0.0193985 0.000881539
+ 2.741e+11Hz -0.0193893 0.000904499
+ 2.742e+11Hz -0.0193797 0.000927668
+ 2.743e+11Hz -0.0193699 0.000951042
+ 2.744e+11Hz -0.0193597 0.000974616
+ 2.745e+11Hz -0.0193493 0.000998386
+ 2.746e+11Hz -0.0193385 0.00102235
+ 2.747e+11Hz -0.0193275 0.0010465
+ 2.748e+11Hz -0.0193161 0.00107083
+ 2.749e+11Hz -0.0193044 0.00109533
+ 2.75e+11Hz -0.0192923 0.00112001
+ 2.751e+11Hz -0.01928 0.00114486
+ 2.752e+11Hz -0.0192673 0.00116986
+ 2.753e+11Hz -0.0192542 0.00119503
+ 2.754e+11Hz -0.0192409 0.00122034
+ 2.755e+11Hz -0.0192271 0.0012458
+ 2.756e+11Hz -0.019213 0.0012714
+ 2.757e+11Hz -0.0191986 0.00129713
+ 2.758e+11Hz -0.0191838 0.00132299
+ 2.759e+11Hz -0.0191686 0.00134898
+ 2.76e+11Hz -0.0191531 0.00137508
+ 2.761e+11Hz -0.0191372 0.00140129
+ 2.762e+11Hz -0.0191209 0.0014276
+ 2.763e+11Hz -0.0191042 0.00145401
+ 2.764e+11Hz -0.0190872 0.00148051
+ 2.765e+11Hz -0.0190698 0.0015071
+ 2.766e+11Hz -0.0190519 0.00153376
+ 2.767e+11Hz -0.0190337 0.0015605
+ 2.768e+11Hz -0.0190151 0.0015873
+ 2.769e+11Hz -0.0189961 0.00161415
+ 2.77e+11Hz -0.0189767 0.00164106
+ 2.771e+11Hz -0.0189569 0.00166802
+ 2.772e+11Hz -0.0189367 0.001695
+ 2.773e+11Hz -0.0189161 0.00172202
+ 2.774e+11Hz -0.018895 0.00174907
+ 2.775e+11Hz -0.0188736 0.00177613
+ 2.776e+11Hz -0.0188518 0.00180319
+ 2.777e+11Hz -0.0188295 0.00183026
+ 2.778e+11Hz -0.0188068 0.00185732
+ 2.779e+11Hz -0.0187837 0.00188437
+ 2.78e+11Hz -0.0187602 0.0019114
+ 2.781e+11Hz -0.0187363 0.0019384
+ 2.782e+11Hz -0.0187119 0.00196536
+ 2.783e+11Hz -0.0186871 0.00199228
+ 2.784e+11Hz -0.0186619 0.00201915
+ 2.785e+11Hz -0.0186363 0.00204596
+ 2.786e+11Hz -0.0186103 0.0020727
+ 2.787e+11Hz -0.0185838 0.00209937
+ 2.788e+11Hz -0.0185569 0.00212596
+ 2.789e+11Hz -0.0185296 0.00215246
+ 2.79e+11Hz -0.0185019 0.00217886
+ 2.791e+11Hz -0.0184737 0.00220516
+ 2.792e+11Hz -0.0184451 0.00223134
+ 2.793e+11Hz -0.0184161 0.00225741
+ 2.794e+11Hz -0.0183867 0.00228334
+ 2.795e+11Hz -0.0183569 0.00230914
+ 2.796e+11Hz -0.0183266 0.0023348
+ 2.797e+11Hz -0.018296 0.00236031
+ 2.798e+11Hz -0.0182649 0.00238565
+ 2.799e+11Hz -0.0182334 0.00241084
+ 2.8e+11Hz -0.0182015 0.00243584
+ 2.801e+11Hz -0.0181691 0.00246067
+ 2.802e+11Hz -0.0181364 0.0024853
+ 2.803e+11Hz -0.0181033 0.00250974
+ 2.804e+11Hz -0.0180698 0.00253398
+ 2.805e+11Hz -0.0180358 0.002558
+ 2.806e+11Hz -0.0180015 0.00258181
+ 2.807e+11Hz -0.0179668 0.00260538
+ 2.808e+11Hz -0.0179317 0.00262873
+ 2.809e+11Hz -0.0178962 0.00265183
+ 2.81e+11Hz -0.0178603 0.00267468
+ 2.811e+11Hz -0.017824 0.00269728
+ 2.812e+11Hz -0.0177874 0.00271962
+ 2.813e+11Hz -0.0177504 0.00274168
+ 2.814e+11Hz -0.017713 0.00276347
+ 2.815e+11Hz -0.0176752 0.00278497
+ 2.816e+11Hz -0.0176371 0.00280619
+ 2.817e+11Hz -0.0175986 0.0028271
+ 2.818e+11Hz -0.0175598 0.00284772
+ 2.819e+11Hz -0.0175207 0.00286802
+ 2.82e+11Hz -0.0174811 0.002888
+ 2.821e+11Hz -0.0174413 0.00290766
+ 2.822e+11Hz -0.0174011 0.00292699
+ 2.823e+11Hz -0.0173606 0.00294599
+ 2.824e+11Hz -0.0173198 0.00296464
+ 2.825e+11Hz -0.0172786 0.00298294
+ 2.826e+11Hz -0.0172372 0.00300089
+ 2.827e+11Hz -0.0171954 0.00301848
+ 2.828e+11Hz -0.0171533 0.0030357
+ 2.829e+11Hz -0.017111 0.00305255
+ 2.83e+11Hz -0.0170683 0.00306903
+ 2.831e+11Hz -0.0170254 0.00308512
+ 2.832e+11Hz -0.0169822 0.00310083
+ 2.833e+11Hz -0.0169388 0.00311614
+ 2.834e+11Hz -0.016895 0.00313105
+ 2.835e+11Hz -0.016851 0.00314556
+ 2.836e+11Hz -0.0168068 0.00315967
+ 2.837e+11Hz -0.0167623 0.00317336
+ 2.838e+11Hz -0.0167176 0.00318664
+ 2.839e+11Hz -0.0166727 0.0031995
+ 2.84e+11Hz -0.0166275 0.00321193
+ 2.841e+11Hz -0.0165821 0.00322393
+ 2.842e+11Hz -0.0165366 0.0032355
+ 2.843e+11Hz -0.0164908 0.00324664
+ 2.844e+11Hz -0.0164448 0.00325733
+ 2.845e+11Hz -0.0163986 0.00326758
+ 2.846e+11Hz -0.0163523 0.00327739
+ 2.847e+11Hz -0.0163058 0.00328674
+ 2.848e+11Hz -0.0162591 0.00329564
+ 2.849e+11Hz -0.0162123 0.00330409
+ 2.85e+11Hz -0.0161653 0.00331208
+ 2.851e+11Hz -0.0161182 0.00331961
+ 2.852e+11Hz -0.016071 0.00332667
+ 2.853e+11Hz -0.0160236 0.00333327
+ 2.854e+11Hz -0.0159762 0.0033394
+ 2.855e+11Hz -0.0159286 0.00334506
+ 2.856e+11Hz -0.0158809 0.00335025
+ 2.857e+11Hz -0.0158331 0.00335497
+ 2.858e+11Hz -0.0157853 0.00335922
+ 2.859e+11Hz -0.0157373 0.00336299
+ 2.86e+11Hz -0.0156893 0.00336628
+ 2.861e+11Hz -0.0156413 0.0033691
+ 2.862e+11Hz -0.0155932 0.00337144
+ 2.863e+11Hz -0.015545 0.0033733
+ 2.864e+11Hz -0.0154969 0.00337469
+ 2.865e+11Hz -0.0154487 0.00337559
+ 2.866e+11Hz -0.0154004 0.00337602
+ 2.867e+11Hz -0.0153522 0.00337596
+ 2.868e+11Hz -0.015304 0.00337543
+ 2.869e+11Hz -0.0152558 0.00337442
+ 2.87e+11Hz -0.0152075 0.00337293
+ 2.871e+11Hz -0.0151594 0.00337097
+ 2.872e+11Hz -0.0151112 0.00336853
+ 2.873e+11Hz -0.0150631 0.00336562
+ 2.874e+11Hz -0.015015 0.00336223
+ 2.875e+11Hz -0.014967 0.00335837
+ 2.876e+11Hz -0.014919 0.00335404
+ 2.877e+11Hz -0.0148712 0.00334925
+ 2.878e+11Hz -0.0148234 0.00334398
+ 2.879e+11Hz -0.0147756 0.00333825
+ 2.88e+11Hz -0.014728 0.00333206
+ 2.881e+11Hz -0.0146805 0.00332541
+ 2.882e+11Hz -0.0146331 0.0033183
+ 2.883e+11Hz -0.0145858 0.00331074
+ 2.884e+11Hz -0.0145386 0.00330273
+ 2.885e+11Hz -0.0144916 0.00329427
+ 2.886e+11Hz -0.0144447 0.00328536
+ 2.887e+11Hz -0.014398 0.003276
+ 2.888e+11Hz -0.0143514 0.00326621
+ 2.889e+11Hz -0.0143049 0.00325599
+ 2.89e+11Hz -0.0142587 0.00324533
+ 2.891e+11Hz -0.0142126 0.00323425
+ 2.892e+11Hz -0.0141666 0.00322274
+ 2.893e+11Hz -0.0141209 0.00321081
+ 2.894e+11Hz -0.0140754 0.00319846
+ 2.895e+11Hz -0.0140301 0.0031857
+ 2.896e+11Hz -0.0139849 0.00317254
+ 2.897e+11Hz -0.01394 0.00315898
+ 2.898e+11Hz -0.0138954 0.00314501
+ 2.899e+11Hz -0.0138509 0.00313066
+ 2.9e+11Hz -0.0138067 0.00311591
+ 2.901e+11Hz -0.0137627 0.00310079
+ 2.902e+11Hz -0.0137189 0.00308528
+ 2.903e+11Hz -0.0136754 0.0030694
+ 2.904e+11Hz -0.0136322 0.00305316
+ 2.905e+11Hz -0.0135892 0.00303656
+ 2.906e+11Hz -0.0135465 0.00301959
+ 2.907e+11Hz -0.0135041 0.00300228
+ 2.908e+11Hz -0.0134619 0.00298463
+ 2.909e+11Hz -0.01342 0.00296663
+ 2.91e+11Hz -0.0133784 0.0029483
+ 2.911e+11Hz -0.0133371 0.00292965
+ 2.912e+11Hz -0.013296 0.00291067
+ 2.913e+11Hz -0.0132553 0.00289138
+ 2.914e+11Hz -0.0132149 0.00287178
+ 2.915e+11Hz -0.0131748 0.00285188
+ 2.916e+11Hz -0.013135 0.00283168
+ 2.917e+11Hz -0.0130955 0.0028112
+ 2.918e+11Hz -0.0130563 0.00279043
+ 2.919e+11Hz -0.0130175 0.00276938
+ 2.92e+11Hz -0.0129789 0.00274806
+ 2.921e+11Hz -0.0129407 0.00272648
+ 2.922e+11Hz -0.0129029 0.00270464
+ 2.923e+11Hz -0.0128653 0.00268255
+ 2.924e+11Hz -0.0128281 0.00266022
+ 2.925e+11Hz -0.0127913 0.00263765
+ 2.926e+11Hz -0.0127547 0.00261485
+ 2.927e+11Hz -0.0127186 0.00259183
+ 2.928e+11Hz -0.0126827 0.00256859
+ 2.929e+11Hz -0.0126472 0.00254514
+ 2.93e+11Hz -0.0126121 0.00252149
+ 2.931e+11Hz -0.0125773 0.00249764
+ 2.932e+11Hz -0.0125429 0.0024736
+ 2.933e+11Hz -0.0125088 0.00244938
+ 2.934e+11Hz -0.012475 0.00242498
+ 2.935e+11Hz -0.0124417 0.00240041
+ 2.936e+11Hz -0.0124087 0.00237569
+ 2.937e+11Hz -0.012376 0.0023508
+ 2.938e+11Hz -0.0123437 0.00232577
+ 2.939e+11Hz -0.0123117 0.00230059
+ 2.94e+11Hz -0.0122801 0.00227528
+ 2.941e+11Hz -0.0122489 0.00224984
+ 2.942e+11Hz -0.012218 0.00222428
+ 2.943e+11Hz -0.0121875 0.00219861
+ 2.944e+11Hz -0.0121574 0.00217282
+ 2.945e+11Hz -0.0121276 0.00214693
+ 2.946e+11Hz -0.0120981 0.00212095
+ 2.947e+11Hz -0.012069 0.00209488
+ 2.948e+11Hz -0.0120403 0.00206872
+ 2.949e+11Hz -0.0120119 0.00204249
+ 2.95e+11Hz -0.0119839 0.00201619
+ 2.951e+11Hz -0.0119562 0.00198983
+ 2.952e+11Hz -0.0119289 0.0019634
+ 2.953e+11Hz -0.0119019 0.00193693
+ 2.954e+11Hz -0.0118753 0.00191041
+ 2.955e+11Hz -0.011849 0.00188385
+ 2.956e+11Hz -0.0118231 0.00185725
+ 2.957e+11Hz -0.0117975 0.00183063
+ 2.958e+11Hz -0.0117722 0.00180398
+ 2.959e+11Hz -0.0117473 0.00177732
+ 2.96e+11Hz -0.0117228 0.00175065
+ 2.961e+11Hz -0.0116985 0.00172397
+ 2.962e+11Hz -0.0116746 0.0016973
+ 2.963e+11Hz -0.011651 0.00167063
+ 2.964e+11Hz -0.0116278 0.00164396
+ 2.965e+11Hz -0.0116048 0.00161732
+ 2.966e+11Hz -0.0115822 0.00159069
+ 2.967e+11Hz -0.0115599 0.00156409
+ 2.968e+11Hz -0.0115379 0.00153752
+ 2.969e+11Hz -0.0115163 0.00151099
+ 2.97e+11Hz -0.0114949 0.0014845
+ 2.971e+11Hz -0.0114738 0.00145805
+ 2.972e+11Hz -0.0114531 0.00143165
+ 2.973e+11Hz -0.0114326 0.0014053
+ 2.974e+11Hz -0.0114124 0.00137901
+ 2.975e+11Hz -0.0113926 0.00135278
+ 2.976e+11Hz -0.011373 0.00132662
+ 2.977e+11Hz -0.0113537 0.00130052
+ 2.978e+11Hz -0.0113347 0.0012745
+ 2.979e+11Hz -0.0113159 0.00124856
+ 2.98e+11Hz -0.0112974 0.00122269
+ 2.981e+11Hz -0.0112792 0.00119691
+ 2.982e+11Hz -0.0112613 0.00117122
+ 2.983e+11Hz -0.0112436 0.00114562
+ 2.984e+11Hz -0.0112262 0.00112011
+ 2.985e+11Hz -0.011209 0.0010947
+ 2.986e+11Hz -0.0111921 0.00106938
+ 2.987e+11Hz -0.0111754 0.00104417
+ 2.988e+11Hz -0.011159 0.00101906
+ 2.989e+11Hz -0.0111428 0.000994064
+ 2.99e+11Hz -0.0111268 0.000969174
+ 2.991e+11Hz -0.0111111 0.000944394
+ 2.992e+11Hz -0.0110956 0.000919729
+ 2.993e+11Hz -0.0110803 0.000895179
+ 2.994e+11Hz -0.0110652 0.000870747
+ 2.995e+11Hz -0.0110503 0.000846435
+ 2.996e+11Hz -0.0110357 0.000822244
+ 2.997e+11Hz -0.0110212 0.000798175
+ 2.998e+11Hz -0.0110069 0.000774231
+ 2.999e+11Hz -0.0109929 0.000750413
+ 3e+11Hz -0.010979 0.000726721
+ ]

.ENDS
.SUBCKT Sub_SPfile_X1 1 2 3
R1N 1 10 -50
R1P 10 11 100
R2N 2 20 -50
R2P 20 21 100

A11 %vd(10 3) %vd(11, 12) xfer1
.model xfer1 xfer R_I=true table=[
+ 0Hz 0.0101636 0
+ 1e+08Hz 0.0101645 2.67428e-05
+ 2e+08Hz 0.0101671 5.34374e-05
+ 3e+08Hz 0.0101713 8.00355e-05
+ 4e+08Hz 0.0101773 0.000106489
+ 5e+08Hz 0.010185 0.00013275
+ 6e+08Hz 0.0101944 0.000158771
+ 7e+08Hz 0.0102055 0.000184505
+ 8e+08Hz 0.0102183 0.000209903
+ 9e+08Hz 0.0102327 0.00023492
+ 1e+09Hz 0.0102488 0.000259509
+ 1.1e+09Hz 0.0102665 0.000283624
+ 1.2e+09Hz 0.0102859 0.00030722
+ 1.3e+09Hz 0.0103069 0.000330251
+ 1.4e+09Hz 0.0103294 0.000352674
+ 1.5e+09Hz 0.0103536 0.000374444
+ 1.6e+09Hz 0.0103793 0.000395519
+ 1.7e+09Hz 0.0104065 0.000415857
+ 1.8e+09Hz 0.0104352 0.000435416
+ 1.9e+09Hz 0.0104654 0.000454156
+ 2e+09Hz 0.0104971 0.000472036
+ 2.1e+09Hz 0.0105302 0.000489017
+ 2.2e+09Hz 0.0105647 0.000505063
+ 2.3e+09Hz 0.0106006 0.000520135
+ 2.4e+09Hz 0.0106378 0.000534198
+ 2.5e+09Hz 0.0106763 0.000547216
+ 2.6e+09Hz 0.0107161 0.000559156
+ 2.7e+09Hz 0.0107572 0.000569984
+ 2.8e+09Hz 0.0107995 0.00057967
+ 2.9e+09Hz 0.010843 0.000588182
+ 3e+09Hz 0.0108876 0.00059549
+ 3.1e+09Hz 0.0109333 0.000601568
+ 3.2e+09Hz 0.0109801 0.000606386
+ 3.3e+09Hz 0.0110279 0.00060992
+ 3.4e+09Hz 0.0110768 0.000612145
+ 3.5e+09Hz 0.0111265 0.000613037
+ 3.6e+09Hz 0.0111773 0.000612574
+ 3.7e+09Hz 0.0112288 0.000610735
+ 3.8e+09Hz 0.0112813 0.000607501
+ 3.9e+09Hz 0.0113345 0.000602854
+ 4e+09Hz 0.0113885 0.000596776
+ 4.1e+09Hz 0.0114432 0.000589251
+ 4.2e+09Hz 0.0114986 0.000580266
+ 4.3e+09Hz 0.0115546 0.000569807
+ 4.4e+09Hz 0.0116112 0.000557862
+ 4.5e+09Hz 0.0116684 0.000544421
+ 4.6e+09Hz 0.0117261 0.000529474
+ 4.7e+09Hz 0.0117842 0.000513014
+ 4.8e+09Hz 0.0118428 0.000495034
+ 4.9e+09Hz 0.0119017 0.000475529
+ 5e+09Hz 0.011961 0.000454494
+ 5.1e+09Hz 0.0120206 0.000431927
+ 5.2e+09Hz 0.0120805 0.000407826
+ 5.3e+09Hz 0.0121405 0.000382191
+ 5.4e+09Hz 0.0122008 0.000355023
+ 5.5e+09Hz 0.0122611 0.000326323
+ 5.6e+09Hz 0.0123216 0.000296095
+ 5.7e+09Hz 0.0123821 0.000264344
+ 5.8e+09Hz 0.0124426 0.000231075
+ 5.9e+09Hz 0.0125031 0.000196294
+ 6e+09Hz 0.0125636 0.00016001
+ 6.1e+09Hz 0.0126239 0.000122231
+ 6.2e+09Hz 0.0126841 8.2968e-05
+ 6.3e+09Hz 0.0127441 4.22309e-05
+ 6.4e+09Hz 0.0128039 3.21247e-08
+ 6.5e+09Hz 0.0128635 -4.36153e-05
+ 6.6e+09Hz 0.0129227 -8.86976e-05
+ 6.7e+09Hz 0.0129816 -0.0001352
+ 6.8e+09Hz 0.0130402 -0.000183106
+ 6.9e+09Hz 0.0130984 -0.000232399
+ 7e+09Hz 0.0131561 -0.000283062
+ 7.1e+09Hz 0.0132134 -0.000335077
+ 7.2e+09Hz 0.0132702 -0.000388424
+ 7.3e+09Hz 0.0133265 -0.000443084
+ 7.4e+09Hz 0.0133822 -0.000499035
+ 7.5e+09Hz 0.0134374 -0.000556257
+ 7.6e+09Hz 0.0134919 -0.000614727
+ 7.7e+09Hz 0.0135458 -0.000674422
+ 7.8e+09Hz 0.0135991 -0.00073532
+ 7.9e+09Hz 0.0136516 -0.000797397
+ 8e+09Hz 0.0137035 -0.000860627
+ 8.1e+09Hz 0.0137546 -0.000924987
+ 8.2e+09Hz 0.0138049 -0.00099045
+ 8.3e+09Hz 0.0138545 -0.00105699
+ 8.4e+09Hz 0.0139033 -0.00112458
+ 8.5e+09Hz 0.0139512 -0.0011932
+ 8.6e+09Hz 0.0139983 -0.00126281
+ 8.7e+09Hz 0.0140446 -0.0013334
+ 8.8e+09Hz 0.0140899 -0.00140493
+ 8.9e+09Hz 0.0141344 -0.00147737
+ 9e+09Hz 0.0141779 -0.00155069
+ 9.1e+09Hz 0.0142206 -0.00162488
+ 9.2e+09Hz 0.0142622 -0.00169989
+ 9.3e+09Hz 0.014303 -0.00177571
+ 9.4e+09Hz 0.0143427 -0.00185229
+ 9.5e+09Hz 0.0143815 -0.00192962
+ 9.6e+09Hz 0.0144193 -0.00200766
+ 9.7e+09Hz 0.0144561 -0.00208638
+ 9.8e+09Hz 0.014492 -0.00216576
+ 9.9e+09Hz 0.0145267 -0.00224576
+ 1e+10Hz 0.0145605 -0.00232636
+ 1.01e+10Hz 0.0145933 -0.00240753
+ 1.02e+10Hz 0.014625 -0.00248923
+ 1.03e+10Hz 0.0146557 -0.00257145
+ 1.04e+10Hz 0.0146854 -0.00265414
+ 1.05e+10Hz 0.014714 -0.00273729
+ 1.06e+10Hz 0.0147416 -0.00282086
+ 1.07e+10Hz 0.0147681 -0.00290483
+ 1.08e+10Hz 0.0147936 -0.00298917
+ 1.09e+10Hz 0.0148181 -0.00307384
+ 1.1e+10Hz 0.0148415 -0.00315883
+ 1.11e+10Hz 0.014864 -0.00324411
+ 1.12e+10Hz 0.0148853 -0.00332965
+ 1.13e+10Hz 0.0149057 -0.00341542
+ 1.14e+10Hz 0.014925 -0.00350139
+ 1.15e+10Hz 0.0149433 -0.00358755
+ 1.16e+10Hz 0.0149607 -0.00367387
+ 1.17e+10Hz 0.014977 -0.00376032
+ 1.18e+10Hz 0.0149923 -0.00384688
+ 1.19e+10Hz 0.0150066 -0.00393352
+ 1.2e+10Hz 0.01502 -0.00402022
+ 1.21e+10Hz 0.0150324 -0.00410697
+ 1.22e+10Hz 0.0150438 -0.00419372
+ 1.23e+10Hz 0.0150543 -0.00428048
+ 1.24e+10Hz 0.0150639 -0.0043672
+ 1.25e+10Hz 0.0150726 -0.00445389
+ 1.26e+10Hz 0.0150803 -0.0045405
+ 1.27e+10Hz 0.0150871 -0.00462703
+ 1.28e+10Hz 0.0150931 -0.00471345
+ 1.29e+10Hz 0.0150982 -0.00479975
+ 1.3e+10Hz 0.0151024 -0.00488591
+ 1.31e+10Hz 0.0151058 -0.00497191
+ 1.32e+10Hz 0.0151084 -0.00505774
+ 1.33e+10Hz 0.0151101 -0.00514338
+ 1.34e+10Hz 0.0151111 -0.00522881
+ 1.35e+10Hz 0.0151113 -0.00531402
+ 1.36e+10Hz 0.0151107 -0.00539901
+ 1.37e+10Hz 0.0151093 -0.00548374
+ 1.38e+10Hz 0.0151073 -0.00556822
+ 1.39e+10Hz 0.0151045 -0.00565243
+ 1.4e+10Hz 0.015101 -0.00573636
+ 1.41e+10Hz 0.0150969 -0.00581999
+ 1.42e+10Hz 0.015092 -0.00590333
+ 1.43e+10Hz 0.0150866 -0.00598636
+ 1.44e+10Hz 0.0150805 -0.00606906
+ 1.45e+10Hz 0.0150738 -0.00615145
+ 1.46e+10Hz 0.0150665 -0.00623349
+ 1.47e+10Hz 0.0150586 -0.0063152
+ 1.48e+10Hz 0.0150501 -0.00639657
+ 1.49e+10Hz 0.0150412 -0.00647758
+ 1.5e+10Hz 0.0150317 -0.00655824
+ 1.51e+10Hz 0.0150216 -0.00663855
+ 1.52e+10Hz 0.0150111 -0.00671849
+ 1.53e+10Hz 0.0150002 -0.00679806
+ 1.54e+10Hz 0.0149887 -0.00687727
+ 1.55e+10Hz 0.0149769 -0.00695612
+ 1.56e+10Hz 0.0149646 -0.00703459
+ 1.57e+10Hz 0.0149519 -0.0071127
+ 1.58e+10Hz 0.0149388 -0.00719044
+ 1.59e+10Hz 0.0149253 -0.00726782
+ 1.6e+10Hz 0.0149115 -0.00734483
+ 1.61e+10Hz 0.0148973 -0.00742147
+ 1.62e+10Hz 0.0148828 -0.00749776
+ 1.63e+10Hz 0.014868 -0.00757369
+ 1.64e+10Hz 0.0148529 -0.00764926
+ 1.65e+10Hz 0.0148375 -0.00772449
+ 1.66e+10Hz 0.0148218 -0.00779937
+ 1.67e+10Hz 0.0148058 -0.00787391
+ 1.68e+10Hz 0.0147897 -0.00794812
+ 1.69e+10Hz 0.0147733 -0.00802199
+ 1.7e+10Hz 0.0147566 -0.00809555
+ 1.71e+10Hz 0.0147398 -0.00816879
+ 1.72e+10Hz 0.0147227 -0.00824172
+ 1.73e+10Hz 0.0147055 -0.00831435
+ 1.74e+10Hz 0.0146881 -0.00838668
+ 1.75e+10Hz 0.0146705 -0.00845873
+ 1.76e+10Hz 0.0146528 -0.00853049
+ 1.77e+10Hz 0.0146349 -0.00860199
+ 1.78e+10Hz 0.0146169 -0.00867323
+ 1.79e+10Hz 0.0145987 -0.00874421
+ 1.8e+10Hz 0.0145804 -0.00881495
+ 1.81e+10Hz 0.014562 -0.00888546
+ 1.82e+10Hz 0.0145435 -0.00895574
+ 1.83e+10Hz 0.0145249 -0.0090258
+ 1.84e+10Hz 0.0145062 -0.00909566
+ 1.85e+10Hz 0.0144874 -0.00916532
+ 1.86e+10Hz 0.0144685 -0.0092348
+ 1.87e+10Hz 0.0144495 -0.0093041
+ 1.88e+10Hz 0.0144305 -0.00937323
+ 1.89e+10Hz 0.0144113 -0.0094422
+ 1.9e+10Hz 0.0143921 -0.00951103
+ 1.91e+10Hz 0.0143728 -0.00957972
+ 1.92e+10Hz 0.0143535 -0.00964828
+ 1.93e+10Hz 0.014334 -0.00971672
+ 1.94e+10Hz 0.0143145 -0.00978506
+ 1.95e+10Hz 0.014295 -0.00985329
+ 1.96e+10Hz 0.0142753 -0.00992144
+ 1.97e+10Hz 0.0142556 -0.00998951
+ 1.98e+10Hz 0.0142358 -0.0100575
+ 1.99e+10Hz 0.014216 -0.0101254
+ 2e+10Hz 0.014196 -0.0101933
+ 2.01e+10Hz 0.014176 -0.0102612
+ 2.02e+10Hz 0.014156 -0.010329
+ 2.03e+10Hz 0.0141358 -0.0103967
+ 2.04e+10Hz 0.0141155 -0.0104645
+ 2.05e+10Hz 0.0140952 -0.0105322
+ 2.06e+10Hz 0.0140748 -0.0106
+ 2.07e+10Hz 0.0140543 -0.0106677
+ 2.08e+10Hz 0.0140336 -0.0107354
+ 2.09e+10Hz 0.0140129 -0.0108032
+ 2.1e+10Hz 0.013992 -0.010871
+ 2.11e+10Hz 0.0139711 -0.0109388
+ 2.12e+10Hz 0.01395 -0.0110067
+ 2.13e+10Hz 0.0139288 -0.0110746
+ 2.14e+10Hz 0.0139074 -0.0111425
+ 2.15e+10Hz 0.0138859 -0.0112105
+ 2.16e+10Hz 0.0138643 -0.0112785
+ 2.17e+10Hz 0.0138425 -0.0113466
+ 2.18e+10Hz 0.0138205 -0.0114148
+ 2.19e+10Hz 0.0137984 -0.011483
+ 2.2e+10Hz 0.0137761 -0.0115513
+ 2.21e+10Hz 0.0137536 -0.0116197
+ 2.22e+10Hz 0.0137309 -0.0116881
+ 2.23e+10Hz 0.0137081 -0.0117566
+ 2.24e+10Hz 0.013685 -0.0118252
+ 2.25e+10Hz 0.0136617 -0.0118939
+ 2.26e+10Hz 0.0136382 -0.0119626
+ 2.27e+10Hz 0.0136144 -0.0120314
+ 2.28e+10Hz 0.0135904 -0.0121003
+ 2.29e+10Hz 0.0135662 -0.0121693
+ 2.3e+10Hz 0.0135417 -0.0122384
+ 2.31e+10Hz 0.013517 -0.0123075
+ 2.32e+10Hz 0.0134919 -0.0123767
+ 2.33e+10Hz 0.0134667 -0.012446
+ 2.34e+10Hz 0.0134411 -0.0125153
+ 2.35e+10Hz 0.0134152 -0.0125848
+ 2.36e+10Hz 0.013389 -0.0126542
+ 2.37e+10Hz 0.0133626 -0.0127238
+ 2.38e+10Hz 0.0133358 -0.0127934
+ 2.39e+10Hz 0.0133087 -0.0128631
+ 2.4e+10Hz 0.0132813 -0.0129328
+ 2.41e+10Hz 0.0132535 -0.0130025
+ 2.42e+10Hz 0.0132254 -0.0130723
+ 2.43e+10Hz 0.013197 -0.0131422
+ 2.44e+10Hz 0.0131682 -0.013212
+ 2.45e+10Hz 0.013139 -0.0132819
+ 2.46e+10Hz 0.0131095 -0.0133519
+ 2.47e+10Hz 0.0130796 -0.0134218
+ 2.48e+10Hz 0.0130494 -0.0134917
+ 2.49e+10Hz 0.0130187 -0.0135617
+ 2.5e+10Hz 0.0129877 -0.0136316
+ 2.51e+10Hz 0.0129563 -0.0137015
+ 2.52e+10Hz 0.0129245 -0.0137714
+ 2.53e+10Hz 0.0128923 -0.0138413
+ 2.54e+10Hz 0.0128597 -0.0139112
+ 2.55e+10Hz 0.0128267 -0.013981
+ 2.56e+10Hz 0.0127933 -0.0140508
+ 2.57e+10Hz 0.0127595 -0.0141205
+ 2.58e+10Hz 0.0127253 -0.0141901
+ 2.59e+10Hz 0.0126907 -0.0142597
+ 2.6e+10Hz 0.0126556 -0.0143292
+ 2.61e+10Hz 0.0126202 -0.0143986
+ 2.62e+10Hz 0.0125843 -0.0144679
+ 2.63e+10Hz 0.012548 -0.0145371
+ 2.64e+10Hz 0.0125113 -0.0146062
+ 2.65e+10Hz 0.0124742 -0.0146751
+ 2.66e+10Hz 0.0124366 -0.014744
+ 2.67e+10Hz 0.0123986 -0.0148127
+ 2.68e+10Hz 0.0123602 -0.0148812
+ 2.69e+10Hz 0.0123214 -0.0149496
+ 2.7e+10Hz 0.0122822 -0.0150178
+ 2.71e+10Hz 0.0122426 -0.0150859
+ 2.72e+10Hz 0.0122025 -0.0151538
+ 2.73e+10Hz 0.0121621 -0.0152215
+ 2.74e+10Hz 0.0121212 -0.015289
+ 2.75e+10Hz 0.0120799 -0.0153563
+ 2.76e+10Hz 0.0120383 -0.0154234
+ 2.77e+10Hz 0.0119962 -0.0154902
+ 2.78e+10Hz 0.0119537 -0.0155569
+ 2.79e+10Hz 0.0119109 -0.0156233
+ 2.8e+10Hz 0.0118676 -0.0156894
+ 2.81e+10Hz 0.011824 -0.0157553
+ 2.82e+10Hz 0.01178 -0.015821
+ 2.83e+10Hz 0.0117356 -0.0158864
+ 2.84e+10Hz 0.0116909 -0.0159515
+ 2.85e+10Hz 0.0116457 -0.0160163
+ 2.86e+10Hz 0.0116003 -0.0160809
+ 2.87e+10Hz 0.0115545 -0.0161451
+ 2.88e+10Hz 0.0115083 -0.0162091
+ 2.89e+10Hz 0.0114618 -0.0162728
+ 2.9e+10Hz 0.0114149 -0.0163361
+ 2.91e+10Hz 0.0113677 -0.0163992
+ 2.92e+10Hz 0.0113203 -0.0164619
+ 2.93e+10Hz 0.0112724 -0.0165243
+ 2.94e+10Hz 0.0112243 -0.0165864
+ 2.95e+10Hz 0.0111759 -0.0166481
+ 2.96e+10Hz 0.0111272 -0.0167095
+ 2.97e+10Hz 0.0110782 -0.0167706
+ 2.98e+10Hz 0.0110289 -0.0168313
+ 2.99e+10Hz 0.0109794 -0.0168917
+ 3e+10Hz 0.0109296 -0.0169518
+ 3.01e+10Hz 0.0108795 -0.0170115
+ 3.02e+10Hz 0.0108292 -0.0170708
+ 3.03e+10Hz 0.0107786 -0.0171298
+ 3.04e+10Hz 0.0107279 -0.0171884
+ 3.05e+10Hz 0.0106768 -0.0172466
+ 3.06e+10Hz 0.0106256 -0.0173045
+ 3.07e+10Hz 0.0105742 -0.017362
+ 3.08e+10Hz 0.0105225 -0.0174192
+ 3.09e+10Hz 0.0104707 -0.017476
+ 3.1e+10Hz 0.0104187 -0.0175324
+ 3.11e+10Hz 0.0103665 -0.0175885
+ 3.12e+10Hz 0.0103141 -0.0176442
+ 3.13e+10Hz 0.0102616 -0.0176996
+ 3.14e+10Hz 0.0102089 -0.0177545
+ 3.15e+10Hz 0.0101561 -0.0178092
+ 3.16e+10Hz 0.0101031 -0.0178634
+ 3.17e+10Hz 0.01005 -0.0179173
+ 3.18e+10Hz 0.00999675 -0.0179709
+ 3.19e+10Hz 0.00994339 -0.018024
+ 3.2e+10Hz 0.00988993 -0.0180769
+ 3.21e+10Hz 0.00983636 -0.0181294
+ 3.22e+10Hz 0.0097827 -0.0181815
+ 3.23e+10Hz 0.00972894 -0.0182333
+ 3.24e+10Hz 0.0096751 -0.0182847
+ 3.25e+10Hz 0.00962118 -0.0183358
+ 3.26e+10Hz 0.00956719 -0.0183866
+ 3.27e+10Hz 0.00951313 -0.0184371
+ 3.28e+10Hz 0.00945901 -0.0184872
+ 3.29e+10Hz 0.00940483 -0.018537
+ 3.3e+10Hz 0.00935061 -0.0185864
+ 3.31e+10Hz 0.00929633 -0.0186356
+ 3.32e+10Hz 0.00924202 -0.0186844
+ 3.33e+10Hz 0.00918768 -0.018733
+ 3.34e+10Hz 0.0091333 -0.0187812
+ 3.35e+10Hz 0.0090789 -0.0188292
+ 3.36e+10Hz 0.00902447 -0.0188768
+ 3.37e+10Hz 0.00897003 -0.0189242
+ 3.38e+10Hz 0.00891557 -0.0189713
+ 3.39e+10Hz 0.0088611 -0.0190181
+ 3.4e+10Hz 0.00880662 -0.0190646
+ 3.41e+10Hz 0.00875213 -0.0191109
+ 3.42e+10Hz 0.00869764 -0.019157
+ 3.43e+10Hz 0.00864315 -0.0192027
+ 3.44e+10Hz 0.00858867 -0.0192483
+ 3.45e+10Hz 0.00853418 -0.0192935
+ 3.46e+10Hz 0.0084797 -0.0193386
+ 3.47e+10Hz 0.00842523 -0.0193834
+ 3.48e+10Hz 0.00837076 -0.019428
+ 3.49e+10Hz 0.0083163 -0.0194724
+ 3.5e+10Hz 0.00826185 -0.0195166
+ 3.51e+10Hz 0.00820741 -0.0195605
+ 3.52e+10Hz 0.00815299 -0.0196043
+ 3.53e+10Hz 0.00809856 -0.0196478
+ 3.54e+10Hz 0.00804415 -0.0196912
+ 3.55e+10Hz 0.00798975 -0.0197344
+ 3.56e+10Hz 0.00793536 -0.0197774
+ 3.57e+10Hz 0.00788097 -0.0198202
+ 3.58e+10Hz 0.00782659 -0.0198629
+ 3.59e+10Hz 0.00777222 -0.0199054
+ 3.6e+10Hz 0.00771784 -0.0199477
+ 3.61e+10Hz 0.00766347 -0.0199899
+ 3.62e+10Hz 0.0076091 -0.0200319
+ 3.63e+10Hz 0.00755472 -0.0200738
+ 3.64e+10Hz 0.00750034 -0.0201156
+ 3.65e+10Hz 0.00744595 -0.0201572
+ 3.66e+10Hz 0.00739156 -0.0201987
+ 3.67e+10Hz 0.00733714 -0.02024
+ 3.68e+10Hz 0.00728271 -0.0202812
+ 3.69e+10Hz 0.00722827 -0.0203223
+ 3.7e+10Hz 0.00717379 -0.0203633
+ 3.71e+10Hz 0.0071193 -0.0204042
+ 3.72e+10Hz 0.00706477 -0.020445
+ 3.73e+10Hz 0.00701021 -0.0204856
+ 3.74e+10Hz 0.00695561 -0.0205262
+ 3.75e+10Hz 0.00690097 -0.0205666
+ 3.76e+10Hz 0.00684628 -0.020607
+ 3.77e+10Hz 0.00679155 -0.0206472
+ 3.78e+10Hz 0.00673676 -0.0206874
+ 3.79e+10Hz 0.00668191 -0.0207274
+ 3.8e+10Hz 0.006627 -0.0207674
+ 3.81e+10Hz 0.00657203 -0.0208073
+ 3.82e+10Hz 0.00651698 -0.020847
+ 3.83e+10Hz 0.00646186 -0.0208867
+ 3.84e+10Hz 0.00640666 -0.0209263
+ 3.85e+10Hz 0.00635137 -0.0209658
+ 3.86e+10Hz 0.00629599 -0.0210052
+ 3.87e+10Hz 0.00624053 -0.0210446
+ 3.88e+10Hz 0.00618496 -0.0210838
+ 3.89e+10Hz 0.00612929 -0.021123
+ 3.9e+10Hz 0.00607351 -0.021162
+ 3.91e+10Hz 0.00601763 -0.021201
+ 3.92e+10Hz 0.00596162 -0.0212399
+ 3.93e+10Hz 0.0059055 -0.0212787
+ 3.94e+10Hz 0.00584925 -0.0213173
+ 3.95e+10Hz 0.00579288 -0.0213559
+ 3.96e+10Hz 0.00573637 -0.0213944
+ 3.97e+10Hz 0.00567972 -0.0214328
+ 3.98e+10Hz 0.00562294 -0.0214711
+ 3.99e+10Hz 0.00556601 -0.0215093
+ 4e+10Hz 0.00550893 -0.0215474
+ 4.01e+10Hz 0.0054517 -0.0215853
+ 4.02e+10Hz 0.00539432 -0.0216232
+ 4.03e+10Hz 0.00533677 -0.0216609
+ 4.04e+10Hz 0.00527907 -0.0216985
+ 4.05e+10Hz 0.0052212 -0.021736
+ 4.06e+10Hz 0.00516316 -0.0217734
+ 4.07e+10Hz 0.00510495 -0.0218106
+ 4.08e+10Hz 0.00504656 -0.0218477
+ 4.09e+10Hz 0.004988 -0.0218846
+ 4.1e+10Hz 0.00492926 -0.0219214
+ 4.11e+10Hz 0.00487034 -0.0219581
+ 4.12e+10Hz 0.00481124 -0.0219946
+ 4.13e+10Hz 0.00475195 -0.022031
+ 4.14e+10Hz 0.00469248 -0.0220671
+ 4.15e+10Hz 0.00463282 -0.0221032
+ 4.16e+10Hz 0.00457296 -0.022139
+ 4.17e+10Hz 0.00451292 -0.0221747
+ 4.18e+10Hz 0.00445269 -0.0222102
+ 4.19e+10Hz 0.00439226 -0.0222455
+ 4.2e+10Hz 0.00433164 -0.0222806
+ 4.21e+10Hz 0.00427083 -0.0223155
+ 4.22e+10Hz 0.00420982 -0.0223503
+ 4.23e+10Hz 0.00414862 -0.0223848
+ 4.24e+10Hz 0.00408723 -0.0224191
+ 4.25e+10Hz 0.00402565 -0.0224532
+ 4.26e+10Hz 0.00396387 -0.0224871
+ 4.27e+10Hz 0.0039019 -0.0225207
+ 4.28e+10Hz 0.00383974 -0.0225541
+ 4.29e+10Hz 0.00377739 -0.0225873
+ 4.3e+10Hz 0.00371485 -0.0226202
+ 4.31e+10Hz 0.00365212 -0.0226529
+ 4.32e+10Hz 0.00358921 -0.0226853
+ 4.33e+10Hz 0.00352612 -0.0227175
+ 4.34e+10Hz 0.00346285 -0.0227494
+ 4.35e+10Hz 0.0033994 -0.0227811
+ 4.36e+10Hz 0.00333577 -0.0228124
+ 4.37e+10Hz 0.00327197 -0.0228435
+ 4.38e+10Hz 0.003208 -0.0228743
+ 4.39e+10Hz 0.00314386 -0.0229049
+ 4.4e+10Hz 0.00307955 -0.0229351
+ 4.41e+10Hz 0.00301509 -0.022965
+ 4.42e+10Hz 0.00295047 -0.0229947
+ 4.43e+10Hz 0.00288569 -0.023024
+ 4.44e+10Hz 0.00282077 -0.0230531
+ 4.45e+10Hz 0.0027557 -0.0230818
+ 4.46e+10Hz 0.00269049 -0.0231102
+ 4.47e+10Hz 0.00262514 -0.0231383
+ 4.48e+10Hz 0.00255965 -0.023166
+ 4.49e+10Hz 0.00249404 -0.0231935
+ 4.5e+10Hz 0.00242831 -0.0232206
+ 4.51e+10Hz 0.00236245 -0.0232473
+ 4.52e+10Hz 0.00229648 -0.0232738
+ 4.53e+10Hz 0.0022304 -0.0232999
+ 4.54e+10Hz 0.00216422 -0.0233256
+ 4.55e+10Hz 0.00209794 -0.0233511
+ 4.56e+10Hz 0.00203156 -0.0233761
+ 4.57e+10Hz 0.0019651 -0.0234008
+ 4.58e+10Hz 0.00189855 -0.0234252
+ 4.59e+10Hz 0.00183192 -0.0234492
+ 4.6e+10Hz 0.00176522 -0.0234729
+ 4.61e+10Hz 0.00169846 -0.0234962
+ 4.62e+10Hz 0.00163163 -0.0235191
+ 4.63e+10Hz 0.00156475 -0.0235417
+ 4.64e+10Hz 0.00149781 -0.023564
+ 4.65e+10Hz 0.00143084 -0.0235858
+ 4.66e+10Hz 0.00136382 -0.0236074
+ 4.67e+10Hz 0.00129677 -0.0236285
+ 4.68e+10Hz 0.00122969 -0.0236493
+ 4.69e+10Hz 0.0011626 -0.0236697
+ 4.7e+10Hz 0.00109548 -0.0236898
+ 4.71e+10Hz 0.00102836 -0.0237095
+ 4.72e+10Hz 0.000961229 -0.0237289
+ 4.73e+10Hz 0.000894101 -0.0237479
+ 4.74e+10Hz 0.00082698 -0.0237665
+ 4.75e+10Hz 0.000759871 -0.0237848
+ 4.76e+10Hz 0.000692779 -0.0238027
+ 4.77e+10Hz 0.00062571 -0.0238202
+ 4.78e+10Hz 0.00055867 -0.0238375
+ 4.79e+10Hz 0.000491664 -0.0238543
+ 4.8e+10Hz 0.000424696 -0.0238708
+ 4.81e+10Hz 0.000357773 -0.023887
+ 4.82e+10Hz 0.000290899 -0.0239028
+ 4.83e+10Hz 0.000224078 -0.0239183
+ 4.84e+10Hz 0.000157317 -0.0239334
+ 4.85e+10Hz 9.06197e-05 -0.0239482
+ 4.86e+10Hz 2.39906e-05 -0.0239626
+ 4.87e+10Hz -4.25655e-05 -0.0239768
+ 4.88e+10Hz -0.000109044 -0.0239906
+ 4.89e+10Hz -0.000175441 -0.024004
+ 4.9e+10Hz -0.000241752 -0.0240172
+ 4.91e+10Hz -0.000307973 -0.02403
+ 4.92e+10Hz -0.0003741 -0.0240425
+ 4.93e+10Hz -0.00044013 -0.0240547
+ 4.94e+10Hz -0.000506057 -0.0240666
+ 4.95e+10Hz -0.00057188 -0.0240781
+ 4.96e+10Hz -0.000637595 -0.0240894
+ 4.97e+10Hz -0.000703198 -0.0241004
+ 4.98e+10Hz -0.000768686 -0.024111
+ 4.99e+10Hz -0.000834056 -0.0241214
+ 5e+10Hz -0.000899306 -0.0241315
+ 5.01e+10Hz -0.000964432 -0.0241413
+ 5.02e+10Hz -0.00102943 -0.0241509
+ 5.03e+10Hz -0.00109431 -0.0241601
+ 5.04e+10Hz -0.00115905 -0.0241691
+ 5.05e+10Hz -0.00122366 -0.0241779
+ 5.06e+10Hz -0.00128814 -0.0241863
+ 5.07e+10Hz -0.00135248 -0.0241945
+ 5.08e+10Hz -0.00141668 -0.0242025
+ 5.09e+10Hz -0.00148074 -0.0242102
+ 5.1e+10Hz -0.00154467 -0.0242176
+ 5.11e+10Hz -0.00160845 -0.0242248
+ 5.12e+10Hz -0.00167209 -0.0242318
+ 5.13e+10Hz -0.00173559 -0.0242386
+ 5.14e+10Hz -0.00179894 -0.0242451
+ 5.15e+10Hz -0.00186215 -0.0242514
+ 5.16e+10Hz -0.00192521 -0.0242575
+ 5.17e+10Hz -0.00198813 -0.0242633
+ 5.18e+10Hz -0.00205091 -0.024269
+ 5.19e+10Hz -0.00211354 -0.0242744
+ 5.2e+10Hz -0.00217602 -0.0242796
+ 5.21e+10Hz -0.00223836 -0.0242847
+ 5.22e+10Hz -0.00230056 -0.0242895
+ 5.23e+10Hz -0.00236261 -0.0242941
+ 5.24e+10Hz -0.00242452 -0.0242986
+ 5.25e+10Hz -0.00248628 -0.0243029
+ 5.26e+10Hz -0.00254791 -0.024307
+ 5.27e+10Hz -0.00260939 -0.0243109
+ 5.28e+10Hz -0.00267074 -0.0243146
+ 5.29e+10Hz -0.00273195 -0.0243182
+ 5.3e+10Hz -0.00279302 -0.0243216
+ 5.31e+10Hz -0.00285395 -0.0243248
+ 5.32e+10Hz -0.00291476 -0.0243278
+ 5.33e+10Hz -0.00297543 -0.0243307
+ 5.34e+10Hz -0.00303596 -0.0243335
+ 5.35e+10Hz -0.00309637 -0.0243361
+ 5.36e+10Hz -0.00315665 -0.0243385
+ 5.37e+10Hz -0.00321681 -0.0243408
+ 5.38e+10Hz -0.00327684 -0.0243429
+ 5.39e+10Hz -0.00333675 -0.0243449
+ 5.4e+10Hz -0.00339654 -0.0243468
+ 5.41e+10Hz -0.00345621 -0.0243485
+ 5.42e+10Hz -0.00351577 -0.02435
+ 5.43e+10Hz -0.00357521 -0.0243514
+ 5.44e+10Hz -0.00363454 -0.0243527
+ 5.45e+10Hz -0.00369376 -0.0243539
+ 5.46e+10Hz -0.00375287 -0.0243549
+ 5.47e+10Hz -0.00381188 -0.0243558
+ 5.48e+10Hz -0.00387078 -0.0243565
+ 5.49e+10Hz -0.00392958 -0.0243571
+ 5.5e+10Hz -0.00398828 -0.0243576
+ 5.51e+10Hz -0.00404688 -0.0243579
+ 5.52e+10Hz -0.00410539 -0.0243581
+ 5.53e+10Hz -0.0041638 -0.0243582
+ 5.54e+10Hz -0.00422212 -0.0243582
+ 5.55e+10Hz -0.00428036 -0.024358
+ 5.56e+10Hz -0.0043385 -0.0243577
+ 5.57e+10Hz -0.00439656 -0.0243572
+ 5.58e+10Hz -0.00445453 -0.0243567
+ 5.59e+10Hz -0.00451242 -0.024356
+ 5.6e+10Hz -0.00457023 -0.0243551
+ 5.61e+10Hz -0.00462796 -0.0243542
+ 5.62e+10Hz -0.00468561 -0.0243531
+ 5.63e+10Hz -0.00474318 -0.0243518
+ 5.64e+10Hz -0.00480068 -0.0243505
+ 5.65e+10Hz -0.0048581 -0.024349
+ 5.66e+10Hz -0.00491546 -0.0243473
+ 5.67e+10Hz -0.00497274 -0.0243455
+ 5.68e+10Hz -0.00502994 -0.0243436
+ 5.69e+10Hz -0.00508708 -0.0243416
+ 5.7e+10Hz -0.00514415 -0.0243394
+ 5.71e+10Hz -0.00520116 -0.024337
+ 5.72e+10Hz -0.00525809 -0.0243345
+ 5.73e+10Hz -0.00531496 -0.0243319
+ 5.74e+10Hz -0.00537176 -0.0243291
+ 5.75e+10Hz -0.00542849 -0.0243262
+ 5.76e+10Hz -0.00548516 -0.0243231
+ 5.77e+10Hz -0.00554176 -0.0243199
+ 5.78e+10Hz -0.00559829 -0.0243165
+ 5.79e+10Hz -0.00565476 -0.024313
+ 5.8e+10Hz -0.00571116 -0.0243093
+ 5.81e+10Hz -0.00576749 -0.0243055
+ 5.82e+10Hz -0.00582376 -0.0243014
+ 5.83e+10Hz -0.00587996 -0.0242973
+ 5.84e+10Hz -0.00593608 -0.0242929
+ 5.85e+10Hz -0.00599214 -0.0242885
+ 5.86e+10Hz -0.00604813 -0.0242838
+ 5.87e+10Hz -0.00610405 -0.024279
+ 5.88e+10Hz -0.00615989 -0.024274
+ 5.89e+10Hz -0.00621566 -0.0242688
+ 5.9e+10Hz -0.00627136 -0.0242635
+ 5.91e+10Hz -0.00632697 -0.0242579
+ 5.92e+10Hz -0.00638251 -0.0242523
+ 5.93e+10Hz -0.00643797 -0.0242464
+ 5.94e+10Hz -0.00649334 -0.0242403
+ 5.95e+10Hz -0.00654863 -0.0242341
+ 5.96e+10Hz -0.00660384 -0.0242277
+ 5.97e+10Hz -0.00665896 -0.0242211
+ 5.98e+10Hz -0.00671398 -0.0242144
+ 5.99e+10Hz -0.00676891 -0.0242074
+ 6e+10Hz -0.00682375 -0.0242003
+ 6.01e+10Hz -0.00687849 -0.024193
+ 6.02e+10Hz -0.00693313 -0.0241855
+ 6.03e+10Hz -0.00698767 -0.0241778
+ 6.04e+10Hz -0.0070421 -0.0241699
+ 6.05e+10Hz -0.00709643 -0.0241618
+ 6.06e+10Hz -0.00715064 -0.0241536
+ 6.07e+10Hz -0.00720474 -0.0241451
+ 6.08e+10Hz -0.00725872 -0.0241365
+ 6.09e+10Hz -0.00731258 -0.0241277
+ 6.1e+10Hz -0.00736632 -0.0241186
+ 6.11e+10Hz -0.00741993 -0.0241095
+ 6.12e+10Hz -0.00747341 -0.0241001
+ 6.13e+10Hz -0.00752677 -0.0240905
+ 6.14e+10Hz -0.00757998 -0.0240807
+ 6.15e+10Hz -0.00763306 -0.0240708
+ 6.16e+10Hz -0.00768599 -0.0240607
+ 6.17e+10Hz -0.00773878 -0.0240503
+ 6.18e+10Hz -0.00779142 -0.0240398
+ 6.19e+10Hz -0.00784391 -0.0240292
+ 6.2e+10Hz -0.00789624 -0.0240183
+ 6.21e+10Hz -0.00794842 -0.0240073
+ 6.22e+10Hz -0.00800043 -0.023996
+ 6.23e+10Hz -0.00805228 -0.0239846
+ 6.24e+10Hz -0.00810396 -0.0239731
+ 6.25e+10Hz -0.00815547 -0.0239613
+ 6.26e+10Hz -0.0082068 -0.0239494
+ 6.27e+10Hz -0.00825796 -0.0239373
+ 6.28e+10Hz -0.00830893 -0.0239251
+ 6.29e+10Hz -0.00835972 -0.0239127
+ 6.3e+10Hz -0.00841033 -0.0239001
+ 6.31e+10Hz -0.00846074 -0.0238874
+ 6.32e+10Hz -0.00851096 -0.0238745
+ 6.33e+10Hz -0.00856098 -0.0238614
+ 6.34e+10Hz -0.00861081 -0.0238482
+ 6.35e+10Hz -0.00866044 -0.0238349
+ 6.36e+10Hz -0.00870986 -0.0238214
+ 6.37e+10Hz -0.00875907 -0.0238078
+ 6.38e+10Hz -0.00880808 -0.023794
+ 6.39e+10Hz -0.00885687 -0.0237801
+ 6.4e+10Hz -0.00890545 -0.0237661
+ 6.41e+10Hz -0.00895382 -0.0237519
+ 6.42e+10Hz -0.00900197 -0.0237377
+ 6.43e+10Hz -0.00904989 -0.0237233
+ 6.44e+10Hz -0.0090976 -0.0237088
+ 6.45e+10Hz -0.00914508 -0.0236941
+ 6.46e+10Hz -0.00919234 -0.0236794
+ 6.47e+10Hz -0.00923937 -0.0236646
+ 6.48e+10Hz -0.00928617 -0.0236497
+ 6.49e+10Hz -0.00933274 -0.0236346
+ 6.5e+10Hz -0.00937908 -0.0236195
+ 6.51e+10Hz -0.00942519 -0.0236043
+ 6.52e+10Hz -0.00947106 -0.0235891
+ 6.53e+10Hz -0.00951671 -0.0235737
+ 6.54e+10Hz -0.00956211 -0.0235583
+ 6.55e+10Hz -0.00960729 -0.0235428
+ 6.56e+10Hz -0.00965222 -0.0235272
+ 6.57e+10Hz -0.00969693 -0.0235116
+ 6.58e+10Hz -0.00974139 -0.023496
+ 6.59e+10Hz -0.00978562 -0.0234802
+ 6.6e+10Hz -0.00982962 -0.0234645
+ 6.61e+10Hz -0.00987338 -0.0234487
+ 6.62e+10Hz -0.0099169 -0.0234329
+ 6.63e+10Hz -0.00996019 -0.023417
+ 6.64e+10Hz -0.0100032 -0.0234011
+ 6.65e+10Hz -0.0100461 -0.0233852
+ 6.66e+10Hz -0.0100887 -0.0233693
+ 6.67e+10Hz -0.010131 -0.0233534
+ 6.68e+10Hz -0.0101732 -0.0233374
+ 6.69e+10Hz -0.0102151 -0.0233215
+ 6.7e+10Hz -0.0102567 -0.0233056
+ 6.71e+10Hz -0.0102982 -0.0232896
+ 6.72e+10Hz -0.0103394 -0.0232737
+ 6.73e+10Hz -0.0103804 -0.0232578
+ 6.74e+10Hz -0.0104212 -0.0232419
+ 6.75e+10Hz -0.0104618 -0.0232261
+ 6.76e+10Hz -0.0105021 -0.0232103
+ 6.77e+10Hz -0.0105423 -0.0231945
+ 6.78e+10Hz -0.0105822 -0.0231787
+ 6.79e+10Hz -0.0106219 -0.023163
+ 6.8e+10Hz -0.0106614 -0.0231473
+ 6.81e+10Hz -0.0107007 -0.0231317
+ 6.82e+10Hz -0.0107399 -0.0231161
+ 6.83e+10Hz -0.0107788 -0.0231006
+ 6.84e+10Hz -0.0108175 -0.0230852
+ 6.85e+10Hz -0.010856 -0.0230698
+ 6.86e+10Hz -0.0108944 -0.0230544
+ 6.87e+10Hz -0.0109326 -0.0230392
+ 6.88e+10Hz -0.0109705 -0.023024
+ 6.89e+10Hz -0.0110084 -0.0230089
+ 6.9e+10Hz -0.011046 -0.0229939
+ 6.91e+10Hz -0.0110835 -0.0229789
+ 6.92e+10Hz -0.0111208 -0.0229641
+ 6.93e+10Hz -0.0111579 -0.0229493
+ 6.94e+10Hz -0.0111949 -0.0229346
+ 6.95e+10Hz -0.0112317 -0.02292
+ 6.96e+10Hz -0.0112684 -0.0229055
+ 6.97e+10Hz -0.0113049 -0.0228911
+ 6.98e+10Hz -0.0113413 -0.0228768
+ 6.99e+10Hz -0.0113776 -0.0228626
+ 7e+10Hz -0.0114137 -0.0228485
+ 7.01e+10Hz -0.0114497 -0.0228345
+ 7.02e+10Hz -0.0114856 -0.0228206
+ 7.03e+10Hz -0.0115213 -0.0228068
+ 7.04e+10Hz -0.0115569 -0.0227931
+ 7.05e+10Hz -0.0115925 -0.0227796
+ 7.06e+10Hz -0.0116279 -0.0227661
+ 7.07e+10Hz -0.0116632 -0.0227527
+ 7.08e+10Hz -0.0116984 -0.0227395
+ 7.09e+10Hz -0.0117335 -0.0227263
+ 7.1e+10Hz -0.0117685 -0.0227133
+ 7.11e+10Hz -0.0118034 -0.0227004
+ 7.12e+10Hz -0.0118383 -0.0226876
+ 7.13e+10Hz -0.011873 -0.0226749
+ 7.14e+10Hz -0.0119077 -0.0226623
+ 7.15e+10Hz -0.0119423 -0.0226498
+ 7.16e+10Hz -0.0119769 -0.0226375
+ 7.17e+10Hz -0.0120113 -0.0226252
+ 7.18e+10Hz -0.0120458 -0.0226131
+ 7.19e+10Hz -0.0120801 -0.0226011
+ 7.2e+10Hz -0.0121144 -0.0225891
+ 7.21e+10Hz -0.0121487 -0.0225773
+ 7.22e+10Hz -0.0121829 -0.0225656
+ 7.23e+10Hz -0.0122171 -0.022554
+ 7.24e+10Hz -0.0122512 -0.0225425
+ 7.25e+10Hz -0.0122853 -0.0225312
+ 7.26e+10Hz -0.0123194 -0.0225199
+ 7.27e+10Hz -0.0123534 -0.0225087
+ 7.28e+10Hz -0.0123875 -0.0224976
+ 7.29e+10Hz -0.0124215 -0.0224866
+ 7.3e+10Hz -0.0124554 -0.0224757
+ 7.31e+10Hz -0.0124894 -0.0224649
+ 7.32e+10Hz -0.0125233 -0.0224542
+ 7.33e+10Hz -0.0125572 -0.0224436
+ 7.34e+10Hz -0.0125912 -0.0224331
+ 7.35e+10Hz -0.0126251 -0.0224227
+ 7.36e+10Hz -0.012659 -0.0224123
+ 7.37e+10Hz -0.0126929 -0.0224021
+ 7.38e+10Hz -0.0127268 -0.0223919
+ 7.39e+10Hz -0.0127607 -0.0223818
+ 7.4e+10Hz -0.0127946 -0.0223718
+ 7.41e+10Hz -0.0128286 -0.0223618
+ 7.42e+10Hz -0.0128625 -0.022352
+ 7.43e+10Hz -0.0128964 -0.0223422
+ 7.44e+10Hz -0.0129304 -0.0223325
+ 7.45e+10Hz -0.0129643 -0.0223228
+ 7.46e+10Hz -0.0129983 -0.0223132
+ 7.47e+10Hz -0.0130323 -0.0223037
+ 7.48e+10Hz -0.0130663 -0.0222942
+ 7.49e+10Hz -0.0131003 -0.0222848
+ 7.5e+10Hz -0.0131344 -0.0222755
+ 7.51e+10Hz -0.0131684 -0.0222662
+ 7.52e+10Hz -0.0132025 -0.022257
+ 7.53e+10Hz -0.0132366 -0.0222478
+ 7.54e+10Hz -0.0132708 -0.0222387
+ 7.55e+10Hz -0.0133049 -0.0222296
+ 7.56e+10Hz -0.0133391 -0.0222205
+ 7.57e+10Hz -0.0133733 -0.0222116
+ 7.58e+10Hz -0.0134075 -0.0222026
+ 7.59e+10Hz -0.0134417 -0.0221937
+ 7.6e+10Hz -0.013476 -0.0221848
+ 7.61e+10Hz -0.0135103 -0.022176
+ 7.62e+10Hz -0.0135446 -0.0221672
+ 7.63e+10Hz -0.0135789 -0.0221585
+ 7.64e+10Hz -0.0136133 -0.0221498
+ 7.65e+10Hz -0.0136477 -0.0221411
+ 7.66e+10Hz -0.0136821 -0.0221324
+ 7.67e+10Hz -0.0137165 -0.0221238
+ 7.68e+10Hz -0.0137509 -0.0221152
+ 7.69e+10Hz -0.0137854 -0.0221066
+ 7.7e+10Hz -0.0138199 -0.0220981
+ 7.71e+10Hz -0.0138544 -0.0220896
+ 7.72e+10Hz -0.0138889 -0.0220811
+ 7.73e+10Hz -0.0139235 -0.0220727
+ 7.74e+10Hz -0.013958 -0.0220642
+ 7.75e+10Hz -0.0139926 -0.0220558
+ 7.76e+10Hz -0.0140272 -0.0220474
+ 7.77e+10Hz -0.0140618 -0.0220391
+ 7.78e+10Hz -0.0140965 -0.0220307
+ 7.79e+10Hz -0.0141311 -0.0220224
+ 7.8e+10Hz -0.0141658 -0.0220141
+ 7.81e+10Hz -0.0142005 -0.0220059
+ 7.82e+10Hz -0.0142352 -0.0219976
+ 7.83e+10Hz -0.0142699 -0.0219894
+ 7.84e+10Hz -0.0143046 -0.0219812
+ 7.85e+10Hz -0.0143394 -0.0219731
+ 7.86e+10Hz -0.0143741 -0.0219649
+ 7.87e+10Hz -0.0144089 -0.0219568
+ 7.88e+10Hz -0.0144436 -0.0219487
+ 7.89e+10Hz -0.0144784 -0.0219407
+ 7.9e+10Hz -0.0145132 -0.0219326
+ 7.91e+10Hz -0.014548 -0.0219246
+ 7.92e+10Hz -0.0145828 -0.0219167
+ 7.93e+10Hz -0.0146176 -0.0219087
+ 7.94e+10Hz -0.0146525 -0.0219008
+ 7.95e+10Hz -0.0146873 -0.021893
+ 7.96e+10Hz -0.0147221 -0.0218852
+ 7.97e+10Hz -0.014757 -0.0218774
+ 7.98e+10Hz -0.0147919 -0.0218696
+ 7.99e+10Hz -0.0148268 -0.0218619
+ 8e+10Hz -0.0148616 -0.0218542
+ 8.01e+10Hz -0.0148965 -0.0218466
+ 8.02e+10Hz -0.0149315 -0.0218391
+ 8.03e+10Hz -0.0149664 -0.0218315
+ 8.04e+10Hz -0.0150013 -0.0218241
+ 8.05e+10Hz -0.0150363 -0.0218166
+ 8.06e+10Hz -0.0150712 -0.0218093
+ 8.07e+10Hz -0.0151062 -0.021802
+ 8.08e+10Hz -0.0151412 -0.0217947
+ 8.09e+10Hz -0.0151762 -0.0217875
+ 8.1e+10Hz -0.0152113 -0.0217804
+ 8.11e+10Hz -0.0152463 -0.0217733
+ 8.12e+10Hz -0.0152814 -0.0217663
+ 8.13e+10Hz -0.0153165 -0.0217594
+ 8.14e+10Hz -0.0153517 -0.0217526
+ 8.15e+10Hz -0.0153868 -0.0217458
+ 8.16e+10Hz -0.015422 -0.0217391
+ 8.17e+10Hz -0.0154573 -0.0217324
+ 8.18e+10Hz -0.0154926 -0.0217259
+ 8.19e+10Hz -0.0155279 -0.0217194
+ 8.2e+10Hz -0.0155632 -0.0217131
+ 8.21e+10Hz -0.0155986 -0.0217068
+ 8.22e+10Hz -0.0156341 -0.0217006
+ 8.23e+10Hz -0.0156696 -0.0216944
+ 8.24e+10Hz -0.0157051 -0.0216884
+ 8.25e+10Hz -0.0157407 -0.0216825
+ 8.26e+10Hz -0.0157764 -0.0216766
+ 8.27e+10Hz -0.0158121 -0.0216709
+ 8.28e+10Hz -0.0158479 -0.0216653
+ 8.29e+10Hz -0.0158838 -0.0216597
+ 8.3e+10Hz -0.0159198 -0.0216543
+ 8.31e+10Hz -0.0159558 -0.021649
+ 8.32e+10Hz -0.0159919 -0.0216437
+ 8.33e+10Hz -0.0160281 -0.0216386
+ 8.34e+10Hz -0.0160645 -0.0216336
+ 8.35e+10Hz -0.0161009 -0.0216287
+ 8.36e+10Hz -0.0161374 -0.0216239
+ 8.37e+10Hz -0.016174 -0.0216192
+ 8.38e+10Hz -0.0162107 -0.0216147
+ 8.39e+10Hz -0.0162476 -0.0216102
+ 8.4e+10Hz -0.0162846 -0.0216058
+ 8.41e+10Hz -0.0163217 -0.0216016
+ 8.42e+10Hz -0.0163589 -0.0215975
+ 8.43e+10Hz -0.0163963 -0.0215935
+ 8.44e+10Hz -0.0164338 -0.0215895
+ 8.45e+10Hz -0.0164715 -0.0215858
+ 8.46e+10Hz -0.0165093 -0.0215821
+ 8.47e+10Hz -0.0165473 -0.0215785
+ 8.48e+10Hz -0.0165855 -0.021575
+ 8.49e+10Hz -0.0166239 -0.0215717
+ 8.5e+10Hz -0.0166624 -0.0215684
+ 8.51e+10Hz -0.0167011 -0.0215653
+ 8.52e+10Hz -0.01674 -0.0215623
+ 8.53e+10Hz -0.0167791 -0.0215593
+ 8.54e+10Hz -0.0168185 -0.0215565
+ 8.55e+10Hz -0.016858 -0.0215538
+ 8.56e+10Hz -0.0168977 -0.0215511
+ 8.57e+10Hz -0.0169377 -0.0215486
+ 8.58e+10Hz -0.0169779 -0.0215461
+ 8.59e+10Hz -0.0170184 -0.0215438
+ 8.6e+10Hz -0.017059 -0.0215415
+ 8.61e+10Hz -0.0171 -0.0215393
+ 8.62e+10Hz -0.0171412 -0.0215372
+ 8.63e+10Hz -0.0171826 -0.0215352
+ 8.64e+10Hz -0.0172243 -0.0215332
+ 8.65e+10Hz -0.0172663 -0.0215313
+ 8.66e+10Hz -0.0173086 -0.0215295
+ 8.67e+10Hz -0.0173512 -0.0215277
+ 8.68e+10Hz -0.0173941 -0.021526
+ 8.69e+10Hz -0.0174372 -0.0215243
+ 8.7e+10Hz -0.0174807 -0.0215227
+ 8.71e+10Hz -0.0175245 -0.0215211
+ 8.72e+10Hz -0.0175686 -0.0215195
+ 8.73e+10Hz -0.017613 -0.021518
+ 8.74e+10Hz -0.0176577 -0.0215165
+ 8.75e+10Hz -0.0177028 -0.021515
+ 8.76e+10Hz -0.0177483 -0.0215135
+ 8.77e+10Hz -0.017794 -0.021512
+ 8.78e+10Hz -0.0178401 -0.0215105
+ 8.79e+10Hz -0.0178866 -0.021509
+ 8.8e+10Hz -0.0179335 -0.0215075
+ 8.81e+10Hz -0.0179807 -0.021506
+ 8.82e+10Hz -0.0180282 -0.0215044
+ 8.83e+10Hz -0.0180762 -0.0215028
+ 8.84e+10Hz -0.0181245 -0.0215012
+ 8.85e+10Hz -0.0181733 -0.0214994
+ 8.86e+10Hz -0.0182224 -0.0214977
+ 8.87e+10Hz -0.0182719 -0.0214958
+ 8.88e+10Hz -0.0183218 -0.0214939
+ 8.89e+10Hz -0.018372 -0.0214919
+ 8.9e+10Hz -0.0184227 -0.0214898
+ 8.91e+10Hz -0.0184739 -0.0214876
+ 8.92e+10Hz -0.0185254 -0.0214852
+ 8.93e+10Hz -0.0185773 -0.0214828
+ 8.94e+10Hz -0.0186296 -0.0214802
+ 8.95e+10Hz -0.0186824 -0.0214774
+ 8.96e+10Hz -0.0187356 -0.0214745
+ 8.97e+10Hz -0.0187892 -0.0214715
+ 8.98e+10Hz -0.0188432 -0.0214683
+ 8.99e+10Hz -0.0188977 -0.0214648
+ 9e+10Hz -0.0189526 -0.0214612
+ 9.01e+10Hz -0.0190079 -0.0214574
+ 9.02e+10Hz -0.0190636 -0.0214534
+ 9.03e+10Hz -0.0191198 -0.0214492
+ 9.04e+10Hz -0.0191764 -0.0214447
+ 9.05e+10Hz -0.0192334 -0.02144
+ 9.06e+10Hz -0.0192909 -0.021435
+ 9.07e+10Hz -0.0193488 -0.0214298
+ 9.08e+10Hz -0.0194071 -0.0214243
+ 9.09e+10Hz -0.0194659 -0.0214185
+ 9.1e+10Hz -0.0195251 -0.0214124
+ 9.11e+10Hz -0.0195847 -0.0214059
+ 9.12e+10Hz -0.0196447 -0.0213992
+ 9.13e+10Hz -0.0197052 -0.0213922
+ 9.14e+10Hz -0.019766 -0.0213848
+ 9.15e+10Hz -0.0198273 -0.021377
+ 9.16e+10Hz -0.0198891 -0.0213689
+ 9.17e+10Hz -0.0199512 -0.0213604
+ 9.18e+10Hz -0.0200137 -0.0213516
+ 9.19e+10Hz -0.0200767 -0.0213423
+ 9.2e+10Hz -0.02014 -0.0213326
+ 9.21e+10Hz -0.0202038 -0.0213225
+ 9.22e+10Hz -0.0202679 -0.021312
+ 9.23e+10Hz -0.0203325 -0.0213011
+ 9.24e+10Hz -0.0203974 -0.0212897
+ 9.25e+10Hz -0.0204627 -0.0212778
+ 9.26e+10Hz -0.0205284 -0.0212655
+ 9.27e+10Hz -0.0205945 -0.0212527
+ 9.28e+10Hz -0.0206609 -0.0212394
+ 9.29e+10Hz -0.0207277 -0.0212256
+ 9.3e+10Hz -0.0207948 -0.0212113
+ 9.31e+10Hz -0.0208623 -0.0211965
+ 9.32e+10Hz -0.0209301 -0.0211811
+ 9.33e+10Hz -0.0209982 -0.0211653
+ 9.34e+10Hz -0.0210667 -0.0211488
+ 9.35e+10Hz -0.0211355 -0.0211318
+ 9.36e+10Hz -0.0212046 -0.0211143
+ 9.37e+10Hz -0.021274 -0.0210961
+ 9.38e+10Hz -0.0213437 -0.0210774
+ 9.39e+10Hz -0.0214137 -0.0210581
+ 9.4e+10Hz -0.0214839 -0.0210382
+ 9.41e+10Hz -0.0215545 -0.0210176
+ 9.42e+10Hz -0.0216253 -0.0209965
+ 9.43e+10Hz -0.0216963 -0.0209747
+ 9.44e+10Hz -0.0217676 -0.0209523
+ 9.45e+10Hz -0.0218391 -0.0209292
+ 9.46e+10Hz -0.0219108 -0.0209055
+ 9.47e+10Hz -0.0219827 -0.0208811
+ 9.48e+10Hz -0.0220549 -0.0208561
+ 9.49e+10Hz -0.0221272 -0.0208304
+ 9.5e+10Hz -0.0221997 -0.020804
+ 9.51e+10Hz -0.0222724 -0.0207769
+ 9.52e+10Hz -0.0223452 -0.0207491
+ 9.53e+10Hz -0.0224182 -0.0207207
+ 9.54e+10Hz -0.0224913 -0.0206915
+ 9.55e+10Hz -0.0225646 -0.0206616
+ 9.56e+10Hz -0.0226379 -0.020631
+ 9.57e+10Hz -0.0227114 -0.0205997
+ 9.58e+10Hz -0.0227849 -0.0205676
+ 9.59e+10Hz -0.0228585 -0.0205349
+ 9.6e+10Hz -0.0229322 -0.0205014
+ 9.61e+10Hz -0.0230059 -0.0204671
+ 9.62e+10Hz -0.0230797 -0.0204321
+ 9.63e+10Hz -0.0231535 -0.0203964
+ 9.64e+10Hz -0.0232273 -0.0203599
+ 9.65e+10Hz -0.0233011 -0.0203227
+ 9.66e+10Hz -0.0233749 -0.0202847
+ 9.67e+10Hz -0.0234487 -0.020246
+ 9.68e+10Hz -0.0235225 -0.0202065
+ 9.69e+10Hz -0.0235962 -0.0201662
+ 9.7e+10Hz -0.0236698 -0.0201252
+ 9.71e+10Hz -0.0237434 -0.0200834
+ 9.72e+10Hz -0.0238169 -0.0200408
+ 9.73e+10Hz -0.0238903 -0.0199975
+ 9.74e+10Hz -0.0239636 -0.0199534
+ 9.75e+10Hz -0.0240367 -0.0199085
+ 9.76e+10Hz -0.0241097 -0.0198629
+ 9.77e+10Hz -0.0241826 -0.0198165
+ 9.78e+10Hz -0.0242553 -0.0197694
+ 9.79e+10Hz -0.0243278 -0.0197214
+ 9.8e+10Hz -0.0244001 -0.0196728
+ 9.81e+10Hz -0.0244723 -0.0196233
+ 9.82e+10Hz -0.0245442 -0.0195731
+ 9.83e+10Hz -0.0246159 -0.0195221
+ 9.84e+10Hz -0.0246873 -0.0194704
+ 9.85e+10Hz -0.0247585 -0.0194179
+ 9.86e+10Hz -0.0248294 -0.0193647
+ 9.87e+10Hz -0.0249001 -0.0193107
+ 9.88e+10Hz -0.0249704 -0.0192559
+ 9.89e+10Hz -0.0250405 -0.0192005
+ 9.9e+10Hz -0.0251102 -0.0191443
+ 9.91e+10Hz -0.0251796 -0.0190873
+ 9.92e+10Hz -0.0252487 -0.0190296
+ 9.93e+10Hz -0.0253174 -0.0189712
+ 9.94e+10Hz -0.0253858 -0.0189121
+ 9.95e+10Hz -0.0254537 -0.0188522
+ 9.96e+10Hz -0.0255213 -0.0187917
+ 9.97e+10Hz -0.0255885 -0.0187304
+ 9.98e+10Hz -0.0256553 -0.0186684
+ 9.99e+10Hz -0.0257216 -0.0186058
+ 1e+11Hz -0.0257875 -0.0185424
+ 1.001e+11Hz -0.025853 -0.0184784
+ 1.002e+11Hz -0.025918 -0.0184137
+ 1.003e+11Hz -0.0259826 -0.0183483
+ 1.004e+11Hz -0.0260467 -0.0182823
+ 1.005e+11Hz -0.0261102 -0.0182156
+ 1.006e+11Hz -0.0261733 -0.0181483
+ 1.007e+11Hz -0.0262359 -0.0180803
+ 1.008e+11Hz -0.026298 -0.0180117
+ 1.009e+11Hz -0.0263595 -0.0179424
+ 1.01e+11Hz -0.0264205 -0.0178726
+ 1.011e+11Hz -0.026481 -0.0178021
+ 1.012e+11Hz -0.0265408 -0.0177311
+ 1.013e+11Hz -0.0266002 -0.0176594
+ 1.014e+11Hz -0.0266589 -0.0175872
+ 1.015e+11Hz -0.0267171 -0.0175144
+ 1.016e+11Hz -0.0267747 -0.017441
+ 1.017e+11Hz -0.0268317 -0.0173671
+ 1.018e+11Hz -0.026888 -0.0172926
+ 1.019e+11Hz -0.0269438 -0.0172176
+ 1.02e+11Hz -0.0269989 -0.017142
+ 1.021e+11Hz -0.0270534 -0.017066
+ 1.022e+11Hz -0.0271073 -0.0169894
+ 1.023e+11Hz -0.0271605 -0.0169124
+ 1.024e+11Hz -0.0272131 -0.0168348
+ 1.025e+11Hz -0.027265 -0.0167568
+ 1.026e+11Hz -0.0273163 -0.0166783
+ 1.027e+11Hz -0.0273669 -0.0165993
+ 1.028e+11Hz -0.0274168 -0.0165199
+ 1.029e+11Hz -0.027466 -0.0164401
+ 1.03e+11Hz -0.0275145 -0.0163599
+ 1.031e+11Hz -0.0275624 -0.0162792
+ 1.032e+11Hz -0.0276095 -0.0161981
+ 1.033e+11Hz -0.027656 -0.0161166
+ 1.034e+11Hz -0.0277017 -0.0160348
+ 1.035e+11Hz -0.0277467 -0.0159526
+ 1.036e+11Hz -0.027791 -0.01587
+ 1.037e+11Hz -0.0278346 -0.0157871
+ 1.038e+11Hz -0.0278775 -0.0157038
+ 1.039e+11Hz -0.0279196 -0.0156202
+ 1.04e+11Hz -0.027961 -0.0155363
+ 1.041e+11Hz -0.0280017 -0.0154521
+ 1.042e+11Hz -0.0280416 -0.0153676
+ 1.043e+11Hz -0.0280808 -0.0152828
+ 1.044e+11Hz -0.0281193 -0.0151977
+ 1.045e+11Hz -0.028157 -0.0151124
+ 1.046e+11Hz -0.028194 -0.0150268
+ 1.047e+11Hz -0.0282302 -0.014941
+ 1.048e+11Hz -0.0282656 -0.0148549
+ 1.049e+11Hz -0.0283004 -0.0147687
+ 1.05e+11Hz -0.0283343 -0.0146822
+ 1.051e+11Hz -0.0283675 -0.0145955
+ 1.052e+11Hz -0.0284 -0.0145087
+ 1.053e+11Hz -0.0284317 -0.0144217
+ 1.054e+11Hz -0.0284627 -0.0143345
+ 1.055e+11Hz -0.0284929 -0.0142472
+ 1.056e+11Hz -0.0285223 -0.0141597
+ 1.057e+11Hz -0.028551 -0.0140721
+ 1.058e+11Hz -0.028579 -0.0139844
+ 1.059e+11Hz -0.0286061 -0.0138966
+ 1.06e+11Hz -0.0286326 -0.0138086
+ 1.061e+11Hz -0.0286583 -0.0137206
+ 1.062e+11Hz -0.0286832 -0.0136325
+ 1.063e+11Hz -0.0287074 -0.0135444
+ 1.064e+11Hz -0.0287308 -0.0134562
+ 1.065e+11Hz -0.0287535 -0.0133679
+ 1.066e+11Hz -0.0287755 -0.0132797
+ 1.067e+11Hz -0.0287967 -0.0131914
+ 1.068e+11Hz -0.0288172 -0.013103
+ 1.069e+11Hz -0.0288369 -0.0130147
+ 1.07e+11Hz -0.0288559 -0.0129264
+ 1.071e+11Hz -0.0288742 -0.0128381
+ 1.072e+11Hz -0.0288917 -0.0127498
+ 1.073e+11Hz -0.0289086 -0.0126615
+ 1.074e+11Hz -0.0289247 -0.0125733
+ 1.075e+11Hz -0.0289401 -0.0124852
+ 1.076e+11Hz -0.0289547 -0.0123971
+ 1.077e+11Hz -0.0289687 -0.0123091
+ 1.078e+11Hz -0.0289819 -0.0122211
+ 1.079e+11Hz -0.0289945 -0.0121333
+ 1.08e+11Hz -0.0290063 -0.0120456
+ 1.081e+11Hz -0.0290175 -0.0119579
+ 1.082e+11Hz -0.029028 -0.0118704
+ 1.083e+11Hz -0.0290377 -0.011783
+ 1.084e+11Hz -0.0290469 -0.0116957
+ 1.085e+11Hz -0.0290553 -0.0116086
+ 1.086e+11Hz -0.029063 -0.0115216
+ 1.087e+11Hz -0.0290701 -0.0114348
+ 1.088e+11Hz -0.0290765 -0.0113481
+ 1.089e+11Hz -0.0290823 -0.0112616
+ 1.09e+11Hz -0.0290874 -0.0111753
+ 1.091e+11Hz -0.0290919 -0.0110892
+ 1.092e+11Hz -0.0290957 -0.0110033
+ 1.093e+11Hz -0.0290989 -0.0109176
+ 1.094e+11Hz -0.0291015 -0.010832
+ 1.095e+11Hz -0.0291035 -0.0107467
+ 1.096e+11Hz -0.0291048 -0.0106617
+ 1.097e+11Hz -0.0291055 -0.0105768
+ 1.098e+11Hz -0.0291056 -0.0104922
+ 1.099e+11Hz -0.0291051 -0.0104078
+ 1.1e+11Hz -0.0291041 -0.0103237
+ 1.101e+11Hz -0.0291024 -0.0102398
+ 1.102e+11Hz -0.0291002 -0.0101562
+ 1.103e+11Hz -0.0290973 -0.0100729
+ 1.104e+11Hz -0.029094 -0.00998981
+ 1.105e+11Hz -0.02909 -0.00990701
+ 1.106e+11Hz -0.0290855 -0.0098245
+ 1.107e+11Hz -0.0290805 -0.00974227
+ 1.108e+11Hz -0.0290749 -0.00966034
+ 1.109e+11Hz -0.0290688 -0.0095787
+ 1.11e+11Hz -0.0290621 -0.00949737
+ 1.111e+11Hz -0.029055 -0.00941634
+ 1.112e+11Hz -0.0290473 -0.00933562
+ 1.113e+11Hz -0.0290391 -0.00925522
+ 1.114e+11Hz -0.0290304 -0.00917514
+ 1.115e+11Hz -0.0290212 -0.00909538
+ 1.116e+11Hz -0.0290116 -0.00901595
+ 1.117e+11Hz -0.0290014 -0.00893685
+ 1.118e+11Hz -0.0289908 -0.00885809
+ 1.119e+11Hz -0.0289797 -0.00877966
+ 1.12e+11Hz -0.0289682 -0.00870158
+ 1.121e+11Hz -0.0289562 -0.00862384
+ 1.122e+11Hz -0.0289438 -0.00854645
+ 1.123e+11Hz -0.0289309 -0.00846941
+ 1.124e+11Hz -0.0289176 -0.00839272
+ 1.125e+11Hz -0.0289039 -0.00831639
+ 1.126e+11Hz -0.0288898 -0.00824042
+ 1.127e+11Hz -0.0288752 -0.00816481
+ 1.128e+11Hz -0.0288603 -0.00808956
+ 1.129e+11Hz -0.0288449 -0.00801468
+ 1.13e+11Hz -0.0288292 -0.00794016
+ 1.131e+11Hz -0.0288131 -0.00786602
+ 1.132e+11Hz -0.0287967 -0.00779224
+ 1.133e+11Hz -0.0287798 -0.00771884
+ 1.134e+11Hz -0.0287626 -0.00764581
+ 1.135e+11Hz -0.0287451 -0.00757315
+ 1.136e+11Hz -0.0287272 -0.00750087
+ 1.137e+11Hz -0.0287089 -0.00742897
+ 1.138e+11Hz -0.0286904 -0.00735745
+ 1.139e+11Hz -0.0286715 -0.0072863
+ 1.14e+11Hz -0.0286523 -0.00721553
+ 1.141e+11Hz -0.0286328 -0.00714514
+ 1.142e+11Hz -0.028613 -0.00707514
+ 1.143e+11Hz -0.0285929 -0.00700551
+ 1.144e+11Hz -0.0285725 -0.00693626
+ 1.145e+11Hz -0.0285518 -0.0068674
+ 1.146e+11Hz -0.0285308 -0.00679891
+ 1.147e+11Hz -0.0285096 -0.0067308
+ 1.148e+11Hz -0.0284881 -0.00666307
+ 1.149e+11Hz -0.0284663 -0.00659573
+ 1.15e+11Hz -0.0284443 -0.00652876
+ 1.151e+11Hz -0.0284221 -0.00646217
+ 1.152e+11Hz -0.0283996 -0.00639595
+ 1.153e+11Hz -0.0283769 -0.00633012
+ 1.154e+11Hz -0.0283539 -0.00626465
+ 1.155e+11Hz -0.0283307 -0.00619957
+ 1.156e+11Hz -0.0283074 -0.00613485
+ 1.157e+11Hz -0.0282838 -0.00607051
+ 1.158e+11Hz -0.02826 -0.00600654
+ 1.159e+11Hz -0.028236 -0.00594293
+ 1.16e+11Hz -0.0282118 -0.0058797
+ 1.161e+11Hz -0.0281874 -0.00581683
+ 1.162e+11Hz -0.0281629 -0.00575432
+ 1.163e+11Hz -0.0281382 -0.00569218
+ 1.164e+11Hz -0.0281133 -0.0056304
+ 1.165e+11Hz -0.0280882 -0.00556897
+ 1.166e+11Hz -0.028063 -0.00550791
+ 1.167e+11Hz -0.0280376 -0.00544719
+ 1.168e+11Hz -0.0280121 -0.00538683
+ 1.169e+11Hz -0.0279864 -0.00532682
+ 1.17e+11Hz -0.0279606 -0.00526716
+ 1.171e+11Hz -0.0279347 -0.00520784
+ 1.172e+11Hz -0.0279086 -0.00514887
+ 1.173e+11Hz -0.0278824 -0.00509024
+ 1.174e+11Hz -0.0278561 -0.00503194
+ 1.175e+11Hz -0.0278297 -0.00497398
+ 1.176e+11Hz -0.0278031 -0.00491635
+ 1.177e+11Hz -0.0277765 -0.00485906
+ 1.178e+11Hz -0.0277497 -0.00480208
+ 1.179e+11Hz -0.0277229 -0.00474544
+ 1.18e+11Hz -0.0276959 -0.00468911
+ 1.181e+11Hz -0.0276689 -0.00463311
+ 1.182e+11Hz -0.0276417 -0.00457742
+ 1.183e+11Hz -0.0276145 -0.00452204
+ 1.184e+11Hz -0.0275872 -0.00446697
+ 1.185e+11Hz -0.0275599 -0.00441221
+ 1.186e+11Hz -0.0275324 -0.00435776
+ 1.187e+11Hz -0.0275049 -0.0043036
+ 1.188e+11Hz -0.0274773 -0.00424974
+ 1.189e+11Hz -0.0274497 -0.00419618
+ 1.19e+11Hz -0.027422 -0.00414291
+ 1.191e+11Hz -0.0273942 -0.00408992
+ 1.192e+11Hz -0.0273664 -0.00403722
+ 1.193e+11Hz -0.0273385 -0.00398481
+ 1.194e+11Hz -0.0273106 -0.00393267
+ 1.195e+11Hz -0.0272826 -0.0038808
+ 1.196e+11Hz -0.0272546 -0.00382921
+ 1.197e+11Hz -0.0272265 -0.00377789
+ 1.198e+11Hz -0.0271984 -0.00372684
+ 1.199e+11Hz -0.0271703 -0.00367604
+ 1.2e+11Hz -0.0271421 -0.00362551
+ 1.201e+11Hz -0.0271139 -0.00357523
+ 1.202e+11Hz -0.0270856 -0.00352521
+ 1.203e+11Hz -0.0270574 -0.00347544
+ 1.204e+11Hz -0.0270291 -0.00342591
+ 1.205e+11Hz -0.0270007 -0.00337663
+ 1.206e+11Hz -0.0269724 -0.00332759
+ 1.207e+11Hz -0.026944 -0.00327878
+ 1.208e+11Hz -0.0269156 -0.00323021
+ 1.209e+11Hz -0.0268872 -0.00318187
+ 1.21e+11Hz -0.0268588 -0.00313376
+ 1.211e+11Hz -0.0268303 -0.00308588
+ 1.212e+11Hz -0.0268019 -0.00303821
+ 1.213e+11Hz -0.0267734 -0.00299077
+ 1.214e+11Hz -0.0267449 -0.00294354
+ 1.215e+11Hz -0.0267164 -0.00289653
+ 1.216e+11Hz -0.0266879 -0.00284973
+ 1.217e+11Hz -0.0266593 -0.00280313
+ 1.218e+11Hz -0.0266308 -0.00275674
+ 1.219e+11Hz -0.0266022 -0.00271055
+ 1.22e+11Hz -0.0265737 -0.00266456
+ 1.221e+11Hz -0.0265451 -0.00261877
+ 1.222e+11Hz -0.0265166 -0.00257317
+ 1.223e+11Hz -0.026488 -0.00252776
+ 1.224e+11Hz -0.0264594 -0.00248255
+ 1.225e+11Hz -0.0264308 -0.00243751
+ 1.226e+11Hz -0.0264022 -0.00239267
+ 1.227e+11Hz -0.0263736 -0.002348
+ 1.228e+11Hz -0.026345 -0.00230351
+ 1.229e+11Hz -0.0263164 -0.0022592
+ 1.23e+11Hz -0.0262878 -0.00221506
+ 1.231e+11Hz -0.0262592 -0.00217109
+ 1.232e+11Hz -0.0262306 -0.0021273
+ 1.233e+11Hz -0.026202 -0.00208367
+ 1.234e+11Hz -0.0261734 -0.0020402
+ 1.235e+11Hz -0.0261447 -0.0019969
+ 1.236e+11Hz -0.0261161 -0.00195375
+ 1.237e+11Hz -0.0260875 -0.00191077
+ 1.238e+11Hz -0.0260589 -0.00186794
+ 1.239e+11Hz -0.0260303 -0.00182527
+ 1.24e+11Hz -0.0260016 -0.00178275
+ 1.241e+11Hz -0.025973 -0.00174038
+ 1.242e+11Hz -0.0259444 -0.00169816
+ 1.243e+11Hz -0.0259157 -0.00165609
+ 1.244e+11Hz -0.0258871 -0.00161416
+ 1.245e+11Hz -0.0258585 -0.00157237
+ 1.246e+11Hz -0.0258299 -0.00153073
+ 1.247e+11Hz -0.0258012 -0.00148922
+ 1.248e+11Hz -0.0257726 -0.00144785
+ 1.249e+11Hz -0.025744 -0.00140662
+ 1.25e+11Hz -0.0257153 -0.00136553
+ 1.251e+11Hz -0.0256867 -0.00132457
+ 1.252e+11Hz -0.0256581 -0.00128374
+ 1.253e+11Hz -0.0256295 -0.00124304
+ 1.254e+11Hz -0.0256008 -0.00120246
+ 1.255e+11Hz -0.0255722 -0.00116202
+ 1.256e+11Hz -0.0255436 -0.0011217
+ 1.257e+11Hz -0.0255149 -0.0010815
+ 1.258e+11Hz -0.0254863 -0.00104143
+ 1.259e+11Hz -0.0254577 -0.00100148
+ 1.26e+11Hz -0.025429 -0.00096165
+ 1.261e+11Hz -0.0254004 -0.000921938
+ 1.262e+11Hz -0.0253718 -0.000882342
+ 1.263e+11Hz -0.0253432 -0.000842863
+ 1.264e+11Hz -0.0253145 -0.000803498
+ 1.265e+11Hz -0.0252859 -0.000764246
+ 1.266e+11Hz -0.0252573 -0.000725106
+ 1.267e+11Hz -0.0252287 -0.000686076
+ 1.268e+11Hz -0.0252001 -0.000647155
+ 1.269e+11Hz -0.0251715 -0.000608342
+ 1.27e+11Hz -0.0251429 -0.000569636
+ 1.271e+11Hz -0.0251143 -0.000531035
+ 1.272e+11Hz -0.0250857 -0.000492537
+ 1.273e+11Hz -0.0250571 -0.000454142
+ 1.274e+11Hz -0.0250285 -0.000415847
+ 1.275e+11Hz -0.0249999 -0.000377653
+ 1.276e+11Hz -0.0249713 -0.000339556
+ 1.277e+11Hz -0.0249427 -0.000301556
+ 1.278e+11Hz -0.0249142 -0.000263652
+ 1.279e+11Hz -0.0248856 -0.000225841
+ 1.28e+11Hz -0.024857 -0.000188123
+ 1.281e+11Hz -0.0248285 -0.000150496
+ 1.282e+11Hz -0.0248 -0.000112958
+ 1.283e+11Hz -0.0247714 -7.55082e-05
+ 1.284e+11Hz -0.0247429 -3.81444e-05
+ 1.285e+11Hz -0.0247144 -8.65244e-07
+ 1.286e+11Hz -0.0246859 3.63309e-05
+ 1.287e+11Hz -0.0246574 7.34458e-05
+ 1.288e+11Hz -0.0246289 0.000110481
+ 1.289e+11Hz -0.0246005 0.000147438
+ 1.29e+11Hz -0.024572 0.00018432
+ 1.291e+11Hz -0.0245436 0.000221127
+ 1.292e+11Hz -0.0245152 0.000257862
+ 1.293e+11Hz -0.0244868 0.000294526
+ 1.294e+11Hz -0.0244584 0.000331122
+ 1.295e+11Hz -0.02443 0.000367652
+ 1.296e+11Hz -0.0244016 0.000404117
+ 1.297e+11Hz -0.0243733 0.00044052
+ 1.298e+11Hz -0.024345 0.000476862
+ 1.299e+11Hz -0.0243166 0.000513147
+ 1.3e+11Hz -0.0242884 0.000549376
+ 1.301e+11Hz -0.0242601 0.000585552
+ 1.302e+11Hz -0.0242318 0.000621676
+ 1.303e+11Hz -0.0242036 0.000657752
+ 1.304e+11Hz -0.0241754 0.000693782
+ 1.305e+11Hz -0.0241472 0.000729768
+ 1.306e+11Hz -0.024119 0.000765713
+ 1.307e+11Hz -0.0240909 0.000801619
+ 1.308e+11Hz -0.0240627 0.000837489
+ 1.309e+11Hz -0.0240346 0.000873326
+ 1.31e+11Hz -0.0240065 0.000909133
+ 1.311e+11Hz -0.0239785 0.000944912
+ 1.312e+11Hz -0.0239504 0.000980667
+ 1.313e+11Hz -0.0239224 0.0010164
+ 1.314e+11Hz -0.0238944 0.00105211
+ 1.315e+11Hz -0.0238664 0.00108781
+ 1.316e+11Hz -0.0238384 0.0011235
+ 1.317e+11Hz -0.0238105 0.00115917
+ 1.318e+11Hz -0.0237826 0.00119484
+ 1.319e+11Hz -0.0237547 0.00123051
+ 1.32e+11Hz -0.0237268 0.00126617
+ 1.321e+11Hz -0.0236989 0.00130184
+ 1.322e+11Hz -0.0236711 0.00133752
+ 1.323e+11Hz -0.0236432 0.00137321
+ 1.324e+11Hz -0.0236154 0.00140891
+ 1.325e+11Hz -0.0235876 0.00144462
+ 1.326e+11Hz -0.0235599 0.00148036
+ 1.327e+11Hz -0.0235321 0.00151612
+ 1.328e+11Hz -0.0235043 0.00155191
+ 1.329e+11Hz -0.0234766 0.00158773
+ 1.33e+11Hz -0.0234489 0.00162358
+ 1.331e+11Hz -0.0234211 0.00165947
+ 1.332e+11Hz -0.0233934 0.00169541
+ 1.333e+11Hz -0.0233657 0.00173139
+ 1.334e+11Hz -0.023338 0.00176742
+ 1.335e+11Hz -0.0233103 0.0018035
+ 1.336e+11Hz -0.0232826 0.00183964
+ 1.337e+11Hz -0.0232549 0.00187584
+ 1.338e+11Hz -0.0232272 0.0019121
+ 1.339e+11Hz -0.0231995 0.00194843
+ 1.34e+11Hz -0.0231717 0.00198484
+ 1.341e+11Hz -0.023144 0.00202131
+ 1.342e+11Hz -0.0231163 0.00205787
+ 1.343e+11Hz -0.0230885 0.00209451
+ 1.344e+11Hz -0.0230607 0.00213124
+ 1.345e+11Hz -0.0230329 0.00216805
+ 1.346e+11Hz -0.0230051 0.00220496
+ 1.347e+11Hz -0.0229772 0.00224197
+ 1.348e+11Hz -0.0229493 0.00227908
+ 1.349e+11Hz -0.0229214 0.00231629
+ 1.35e+11Hz -0.0228934 0.00235361
+ 1.351e+11Hz -0.0228654 0.00239104
+ 1.352e+11Hz -0.0228373 0.00242858
+ 1.353e+11Hz -0.0228092 0.00246625
+ 1.354e+11Hz -0.022781 0.00250403
+ 1.355e+11Hz -0.0227528 0.00254194
+ 1.356e+11Hz -0.0227245 0.00257997
+ 1.357e+11Hz -0.0226961 0.00261814
+ 1.358e+11Hz -0.0226677 0.00265644
+ 1.359e+11Hz -0.0226392 0.00269488
+ 1.36e+11Hz -0.0226106 0.00273345
+ 1.361e+11Hz -0.0225819 0.00277217
+ 1.362e+11Hz -0.0225531 0.00281103
+ 1.363e+11Hz -0.0225242 0.00285004
+ 1.364e+11Hz -0.0224952 0.0028892
+ 1.365e+11Hz -0.0224662 0.00292851
+ 1.366e+11Hz -0.0224369 0.00296798
+ 1.367e+11Hz -0.0224076 0.0030076
+ 1.368e+11Hz -0.0223782 0.00304738
+ 1.369e+11Hz -0.0223486 0.00308732
+ 1.37e+11Hz -0.0223188 0.00312742
+ 1.371e+11Hz -0.0222889 0.00316769
+ 1.372e+11Hz -0.0222589 0.00320812
+ 1.373e+11Hz -0.0222287 0.00324872
+ 1.374e+11Hz -0.0221984 0.00328949
+ 1.375e+11Hz -0.0221679 0.00333042
+ 1.376e+11Hz -0.0221372 0.00337153
+ 1.377e+11Hz -0.0221063 0.0034128
+ 1.378e+11Hz -0.0220752 0.00345425
+ 1.379e+11Hz -0.0220439 0.00349587
+ 1.38e+11Hz -0.0220124 0.00353766
+ 1.381e+11Hz -0.0219807 0.00357963
+ 1.382e+11Hz -0.0219488 0.00362176
+ 1.383e+11Hz -0.0219167 0.00366407
+ 1.384e+11Hz -0.0218843 0.00370655
+ 1.385e+11Hz -0.0218517 0.0037492
+ 1.386e+11Hz -0.0218188 0.00379202
+ 1.387e+11Hz -0.0217857 0.00383501
+ 1.388e+11Hz -0.0217523 0.00387816
+ 1.389e+11Hz -0.0217187 0.00392149
+ 1.39e+11Hz -0.0216847 0.00396498
+ 1.391e+11Hz -0.0216505 0.00400863
+ 1.392e+11Hz -0.021616 0.00405245
+ 1.393e+11Hz -0.0215812 0.00409642
+ 1.394e+11Hz -0.021546 0.00414055
+ 1.395e+11Hz -0.0215106 0.00418484
+ 1.396e+11Hz -0.0214748 0.00422928
+ 1.397e+11Hz -0.0214387 0.00427387
+ 1.398e+11Hz -0.0214023 0.0043186
+ 1.399e+11Hz -0.0213655 0.00436348
+ 1.4e+11Hz -0.0213284 0.0044085
+ 1.401e+11Hz -0.0212909 0.00445365
+ 1.402e+11Hz -0.021253 0.00449893
+ 1.403e+11Hz -0.0212147 0.00454434
+ 1.404e+11Hz -0.0211761 0.00458988
+ 1.405e+11Hz -0.0211371 0.00463553
+ 1.406e+11Hz -0.0210976 0.0046813
+ 1.407e+11Hz -0.0210578 0.00472717
+ 1.408e+11Hz -0.0210175 0.00477315
+ 1.409e+11Hz -0.0209769 0.00481923
+ 1.41e+11Hz -0.0209358 0.0048654
+ 1.411e+11Hz -0.0208942 0.00491165
+ 1.412e+11Hz -0.0208523 0.00495799
+ 1.413e+11Hz -0.0208098 0.0050044
+ 1.414e+11Hz -0.0207669 0.00505088
+ 1.415e+11Hz -0.0207236 0.00509742
+ 1.416e+11Hz -0.0206798 0.00514402
+ 1.417e+11Hz -0.0206355 0.00519066
+ 1.418e+11Hz -0.0205907 0.00523734
+ 1.419e+11Hz -0.0205455 0.00528406
+ 1.42e+11Hz -0.0204997 0.0053308
+ 1.421e+11Hz -0.0204535 0.00537756
+ 1.422e+11Hz -0.0204067 0.00542433
+ 1.423e+11Hz -0.0203595 0.00547111
+ 1.424e+11Hz -0.0203117 0.00551787
+ 1.425e+11Hz -0.0202634 0.00556462
+ 1.426e+11Hz -0.0202146 0.00561135
+ 1.427e+11Hz -0.0201652 0.00565804
+ 1.428e+11Hz -0.0201154 0.00570469
+ 1.429e+11Hz -0.0200649 0.00575129
+ 1.43e+11Hz -0.020014 0.00579784
+ 1.431e+11Hz -0.0199625 0.00584431
+ 1.432e+11Hz -0.0199104 0.0058907
+ 1.433e+11Hz -0.0198578 0.00593701
+ 1.434e+11Hz -0.0198046 0.00598321
+ 1.435e+11Hz -0.0197509 0.00602931
+ 1.436e+11Hz -0.0196966 0.00607529
+ 1.437e+11Hz -0.0196417 0.00612115
+ 1.438e+11Hz -0.0195863 0.00616686
+ 1.439e+11Hz -0.0195302 0.00621243
+ 1.44e+11Hz -0.0194737 0.00625783
+ 1.441e+11Hz -0.0194165 0.00630307
+ 1.442e+11Hz -0.0193588 0.00634812
+ 1.443e+11Hz -0.0193004 0.00639299
+ 1.444e+11Hz -0.0192416 0.00643765
+ 1.445e+11Hz -0.0191821 0.00648209
+ 1.446e+11Hz -0.019122 0.00652632
+ 1.447e+11Hz -0.0190614 0.00657031
+ 1.448e+11Hz -0.0190002 0.00661405
+ 1.449e+11Hz -0.0189384 0.00665754
+ 1.45e+11Hz -0.018876 0.00670075
+ 1.451e+11Hz -0.018813 0.00674369
+ 1.452e+11Hz -0.0187495 0.00678634
+ 1.453e+11Hz -0.0186853 0.00682868
+ 1.454e+11Hz -0.0186206 0.00687072
+ 1.455e+11Hz -0.0185553 0.00691243
+ 1.456e+11Hz -0.0184895 0.0069538
+ 1.457e+11Hz -0.0184231 0.00699483
+ 1.458e+11Hz -0.0183561 0.0070355
+ 1.459e+11Hz -0.0182885 0.0070758
+ 1.46e+11Hz -0.0182204 0.00711572
+ 1.461e+11Hz -0.0181517 0.00715525
+ 1.462e+11Hz -0.0180825 0.00719438
+ 1.463e+11Hz -0.0180127 0.00723309
+ 1.464e+11Hz -0.0179423 0.00727138
+ 1.465e+11Hz -0.0178715 0.00730924
+ 1.466e+11Hz -0.0178 0.00734665
+ 1.467e+11Hz -0.0177281 0.00738361
+ 1.468e+11Hz -0.0176556 0.0074201
+ 1.469e+11Hz -0.0175826 0.00745611
+ 1.47e+11Hz -0.017509 0.00749164
+ 1.471e+11Hz -0.017435 0.00752666
+ 1.472e+11Hz -0.0173604 0.00756118
+ 1.473e+11Hz -0.0172853 0.00759519
+ 1.474e+11Hz -0.0172098 0.00762866
+ 1.475e+11Hz -0.0171337 0.0076616
+ 1.476e+11Hz -0.0170572 0.00769399
+ 1.477e+11Hz -0.0169802 0.00772582
+ 1.478e+11Hz -0.0169027 0.00775709
+ 1.479e+11Hz -0.0168248 0.00778778
+ 1.48e+11Hz -0.0167464 0.00781789
+ 1.481e+11Hz -0.0166676 0.00784741
+ 1.482e+11Hz -0.0165883 0.00787632
+ 1.483e+11Hz -0.0165086 0.00790463
+ 1.484e+11Hz -0.0164285 0.00793231
+ 1.485e+11Hz -0.016348 0.00795937
+ 1.486e+11Hz -0.0162671 0.0079858
+ 1.487e+11Hz -0.0161858 0.00801158
+ 1.488e+11Hz -0.0161041 0.00803671
+ 1.489e+11Hz -0.016022 0.00806118
+ 1.49e+11Hz -0.0159396 0.008085
+ 1.491e+11Hz -0.0158568 0.00810813
+ 1.492e+11Hz -0.0157737 0.0081306
+ 1.493e+11Hz -0.0156902 0.00815237
+ 1.494e+11Hz -0.0156064 0.00817346
+ 1.495e+11Hz -0.0155223 0.00819385
+ 1.496e+11Hz -0.0154379 0.00821354
+ 1.497e+11Hz -0.0153532 0.00823252
+ 1.498e+11Hz -0.0152682 0.00825078
+ 1.499e+11Hz -0.015183 0.00826833
+ 1.5e+11Hz -0.0150974 0.00828515
+ 1.501e+11Hz -0.0150117 0.00830125
+ 1.502e+11Hz -0.0149257 0.00831661
+ 1.503e+11Hz -0.0148395 0.00833124
+ 1.504e+11Hz -0.014753 0.00834513
+ 1.505e+11Hz -0.0146664 0.00835827
+ 1.506e+11Hz -0.0145795 0.00837066
+ 1.507e+11Hz -0.0144925 0.00838231
+ 1.508e+11Hz -0.0144053 0.0083932
+ 1.509e+11Hz -0.014318 0.00840334
+ 1.51e+11Hz -0.0142305 0.00841272
+ 1.511e+11Hz -0.0141429 0.00842133
+ 1.512e+11Hz -0.0140551 0.00842919
+ 1.513e+11Hz -0.0139673 0.00843628
+ 1.514e+11Hz -0.0138793 0.00844261
+ 1.515e+11Hz -0.0137912 0.00844817
+ 1.516e+11Hz -0.0137031 0.00845296
+ 1.517e+11Hz -0.0136149 0.00845699
+ 1.518e+11Hz -0.0135267 0.00846025
+ 1.519e+11Hz -0.0134384 0.00846274
+ 1.52e+11Hz -0.01335 0.00846446
+ 1.521e+11Hz -0.0132617 0.00846541
+ 1.522e+11Hz -0.0131733 0.0084656
+ 1.523e+11Hz -0.013085 0.00846502
+ 1.524e+11Hz -0.0129967 0.00846368
+ 1.525e+11Hz -0.0129084 0.00846157
+ 1.526e+11Hz -0.0128201 0.0084587
+ 1.527e+11Hz -0.0127319 0.00845507
+ 1.528e+11Hz -0.0126437 0.00845069
+ 1.529e+11Hz -0.0125556 0.00844555
+ 1.53e+11Hz -0.0124676 0.00843965
+ 1.531e+11Hz -0.0123797 0.008433
+ 1.532e+11Hz -0.0122919 0.00842561
+ 1.533e+11Hz -0.0122042 0.00841747
+ 1.534e+11Hz -0.0121166 0.00840859
+ 1.535e+11Hz -0.0120292 0.00839898
+ 1.536e+11Hz -0.0119419 0.00838863
+ 1.537e+11Hz -0.0118547 0.00837755
+ 1.538e+11Hz -0.0117678 0.00836574
+ 1.539e+11Hz -0.011681 0.00835321
+ 1.54e+11Hz -0.0115943 0.00833997
+ 1.541e+11Hz -0.0115079 0.00832601
+ 1.542e+11Hz -0.0114217 0.00831135
+ 1.543e+11Hz -0.0113357 0.00829598
+ 1.544e+11Hz -0.0112499 0.00827992
+ 1.545e+11Hz -0.0111644 0.00826317
+ 1.546e+11Hz -0.0110791 0.00824573
+ 1.547e+11Hz -0.010994 0.00822761
+ 1.548e+11Hz -0.0109092 0.00820881
+ 1.549e+11Hz -0.0108246 0.00818935
+ 1.55e+11Hz -0.0107404 0.00816922
+ 1.551e+11Hz -0.0106564 0.00814844
+ 1.552e+11Hz -0.0105727 0.00812701
+ 1.553e+11Hz -0.0104893 0.00810493
+ 1.554e+11Hz -0.0104062 0.00808222
+ 1.555e+11Hz -0.0103234 0.00805888
+ 1.556e+11Hz -0.010241 0.00803491
+ 1.557e+11Hz -0.0101589 0.00801033
+ 1.558e+11Hz -0.0100771 0.00798514
+ 1.559e+11Hz -0.00999559 0.00795935
+ 1.56e+11Hz -0.00991448 0.00793296
+ 1.561e+11Hz -0.00983372 0.00790598
+ 1.562e+11Hz -0.00975332 0.00787842
+ 1.563e+11Hz -0.00967328 0.00785029
+ 1.564e+11Hz -0.00959362 0.0078216
+ 1.565e+11Hz -0.00951433 0.00779234
+ 1.566e+11Hz -0.00943542 0.00776254
+ 1.567e+11Hz -0.00935689 0.00773219
+ 1.568e+11Hz -0.00927876 0.00770131
+ 1.569e+11Hz -0.00920103 0.00766989
+ 1.57e+11Hz -0.00912369 0.00763796
+ 1.571e+11Hz -0.00904676 0.00760552
+ 1.572e+11Hz -0.00897024 0.00757257
+ 1.573e+11Hz -0.00889413 0.00753913
+ 1.574e+11Hz -0.00881843 0.0075052
+ 1.575e+11Hz -0.00874316 0.00747078
+ 1.576e+11Hz -0.00866831 0.0074359
+ 1.577e+11Hz -0.00859389 0.00740055
+ 1.578e+11Hz -0.0085199 0.00736474
+ 1.579e+11Hz -0.00844634 0.00732848
+ 1.58e+11Hz -0.00837322 0.00729178
+ 1.581e+11Hz -0.00830054 0.00725464
+ 1.582e+11Hz -0.0082283 0.00721708
+ 1.583e+11Hz -0.0081565 0.0071791
+ 1.584e+11Hz -0.00808515 0.00714071
+ 1.585e+11Hz -0.00801424 0.00710191
+ 1.586e+11Hz -0.00794379 0.00706272
+ 1.587e+11Hz -0.00787378 0.00702314
+ 1.588e+11Hz -0.00780423 0.00698319
+ 1.589e+11Hz -0.00773513 0.00694285
+ 1.59e+11Hz -0.00766649 0.00690216
+ 1.591e+11Hz -0.0075983 0.0068611
+ 1.592e+11Hz -0.00753057 0.00681969
+ 1.593e+11Hz -0.0074633 0.00677794
+ 1.594e+11Hz -0.00739648 0.00673586
+ 1.595e+11Hz -0.00733013 0.00669344
+ 1.596e+11Hz -0.00726423 0.0066507
+ 1.597e+11Hz -0.0071988 0.00660765
+ 1.598e+11Hz -0.00713382 0.00656429
+ 1.599e+11Hz -0.0070693 0.00652063
+ 1.6e+11Hz -0.00700524 0.00647667
+ 1.601e+11Hz -0.00694165 0.00643242
+ 1.602e+11Hz -0.00687851 0.0063879
+ 1.603e+11Hz -0.00681582 0.0063431
+ 1.604e+11Hz -0.0067536 0.00629803
+ 1.605e+11Hz -0.00669184 0.00625269
+ 1.606e+11Hz -0.00663053 0.00620711
+ 1.607e+11Hz -0.00656967 0.00616127
+ 1.608e+11Hz -0.00650927 0.00611519
+ 1.609e+11Hz -0.00644933 0.00606888
+ 1.61e+11Hz -0.00638984 0.00602233
+ 1.611e+11Hz -0.0063308 0.00597556
+ 1.612e+11Hz -0.00627221 0.00592856
+ 1.613e+11Hz -0.00621407 0.00588136
+ 1.614e+11Hz -0.00615637 0.00583394
+ 1.615e+11Hz -0.00609913 0.00578633
+ 1.616e+11Hz -0.00604233 0.00573851
+ 1.617e+11Hz -0.00598597 0.00569051
+ 1.618e+11Hz -0.00593005 0.00564231
+ 1.619e+11Hz -0.00587457 0.00559394
+ 1.62e+11Hz -0.00581954 0.00554538
+ 1.621e+11Hz -0.00576493 0.00549666
+ 1.622e+11Hz -0.00571077 0.00544777
+ 1.623e+11Hz -0.00565703 0.00539872
+ 1.624e+11Hz -0.00560373 0.00534951
+ 1.625e+11Hz -0.00555085 0.00530015
+ 1.626e+11Hz -0.0054984 0.00525063
+ 1.627e+11Hz -0.00544638 0.00520098
+ 1.628e+11Hz -0.00539478 0.00515119
+ 1.629e+11Hz -0.0053436 0.00510126
+ 1.63e+11Hz -0.00529284 0.0050512
+ 1.631e+11Hz -0.0052425 0.00500101
+ 1.632e+11Hz -0.00519257 0.0049507
+ 1.633e+11Hz -0.00514306 0.00490027
+ 1.634e+11Hz -0.00509395 0.00484972
+ 1.635e+11Hz -0.00504525 0.00479907
+ 1.636e+11Hz -0.00499696 0.0047483
+ 1.637e+11Hz -0.00494908 0.00469743
+ 1.638e+11Hz -0.00490159 0.00464646
+ 1.639e+11Hz -0.00485451 0.0045954
+ 1.64e+11Hz -0.00480782 0.00454424
+ 1.641e+11Hz -0.00476153 0.00449299
+ 1.642e+11Hz -0.00471563 0.00444165
+ 1.643e+11Hz -0.00467012 0.00439023
+ 1.644e+11Hz -0.004625 0.00433873
+ 1.645e+11Hz -0.00458027 0.00428715
+ 1.646e+11Hz -0.00453592 0.00423549
+ 1.647e+11Hz -0.00449195 0.00418377
+ 1.648e+11Hz -0.00444837 0.00413197
+ 1.649e+11Hz -0.00440516 0.00408011
+ 1.65e+11Hz -0.00436232 0.00402819
+ 1.651e+11Hz -0.00431987 0.0039762
+ 1.652e+11Hz -0.00427778 0.00392416
+ 1.653e+11Hz -0.00423606 0.00387206
+ 1.654e+11Hz -0.00419471 0.00381991
+ 1.655e+11Hz -0.00415373 0.00376771
+ 1.656e+11Hz -0.0041131 0.00371547
+ 1.657e+11Hz -0.00407284 0.00366317
+ 1.658e+11Hz -0.00403294 0.00361084
+ 1.659e+11Hz -0.0039934 0.00355846
+ 1.66e+11Hz -0.00395421 0.00350605
+ 1.661e+11Hz -0.00391537 0.0034536
+ 1.662e+11Hz -0.00387689 0.00340112
+ 1.663e+11Hz -0.00383875 0.00334861
+ 1.664e+11Hz -0.00380096 0.00329607
+ 1.665e+11Hz -0.00376352 0.0032435
+ 1.666e+11Hz -0.00372642 0.00319091
+ 1.667e+11Hz -0.00368966 0.00313829
+ 1.668e+11Hz -0.00365324 0.00308566
+ 1.669e+11Hz -0.00361716 0.003033
+ 1.67e+11Hz -0.00358141 0.00298034
+ 1.671e+11Hz -0.003546 0.00292765
+ 1.672e+11Hz -0.00351092 0.00287496
+ 1.673e+11Hz -0.00347617 0.00282225
+ 1.674e+11Hz -0.00344175 0.00276954
+ 1.675e+11Hz -0.00340765 0.00271682
+ 1.676e+11Hz -0.00337388 0.0026641
+ 1.677e+11Hz -0.00334043 0.00261137
+ 1.678e+11Hz -0.0033073 0.00255864
+ 1.679e+11Hz -0.0032745 0.00250592
+ 1.68e+11Hz -0.003242 0.0024532
+ 1.681e+11Hz -0.00320983 0.00240048
+ 1.682e+11Hz -0.00317796 0.00234777
+ 1.683e+11Hz -0.00314641 0.00229507
+ 1.684e+11Hz -0.00311517 0.00224238
+ 1.685e+11Hz -0.00308424 0.0021897
+ 1.686e+11Hz -0.00305361 0.00213704
+ 1.687e+11Hz -0.00302329 0.00208439
+ 1.688e+11Hz -0.00299327 0.00203176
+ 1.689e+11Hz -0.00296355 0.00197915
+ 1.69e+11Hz -0.00293413 0.00192656
+ 1.691e+11Hz -0.00290501 0.00187399
+ 1.692e+11Hz -0.00287618 0.00182145
+ 1.693e+11Hz -0.00284765 0.00176893
+ 1.694e+11Hz -0.00281941 0.00171644
+ 1.695e+11Hz -0.00279146 0.00166398
+ 1.696e+11Hz -0.0027638 0.00161156
+ 1.697e+11Hz -0.00273642 0.00155916
+ 1.698e+11Hz -0.00270933 0.0015068
+ 1.699e+11Hz -0.00268252 0.00145447
+ 1.7e+11Hz -0.00265599 0.00140219
+ 1.701e+11Hz -0.00262975 0.00134994
+ 1.702e+11Hz -0.00260377 0.00129773
+ 1.703e+11Hz -0.00257808 0.00124556
+ 1.704e+11Hz -0.00255265 0.00119344
+ 1.705e+11Hz -0.0025275 0.00114136
+ 1.706e+11Hz -0.00250262 0.00108933
+ 1.707e+11Hz -0.00247801 0.00103735
+ 1.708e+11Hz -0.00245366 0.000985415
+ 1.709e+11Hz -0.00242957 0.000933532
+ 1.71e+11Hz -0.00240575 0.000881702
+ 1.711e+11Hz -0.00238219 0.000829926
+ 1.712e+11Hz -0.00235888 0.000778204
+ 1.713e+11Hz -0.00233583 0.000726539
+ 1.714e+11Hz -0.00231304 0.000674932
+ 1.715e+11Hz -0.00229049 0.000623384
+ 1.716e+11Hz -0.0022682 0.000571896
+ 1.717e+11Hz -0.00224615 0.000520469
+ 1.718e+11Hz -0.00222435 0.000469105
+ 1.719e+11Hz -0.00220279 0.000417805
+ 1.72e+11Hz -0.00218148 0.000366571
+ 1.721e+11Hz -0.0021604 0.000315402
+ 1.722e+11Hz -0.00213956 0.000264301
+ 1.723e+11Hz -0.00211896 0.000213268
+ 1.724e+11Hz -0.00209859 0.000162304
+ 1.725e+11Hz -0.00207845 0.000111411
+ 1.726e+11Hz -0.00205854 6.05895e-05
+ 1.727e+11Hz -0.00203886 9.84029e-06
+ 1.728e+11Hz -0.0020194 -4.08356e-05
+ 1.729e+11Hz -0.00200017 -9.14372e-05
+ 1.73e+11Hz -0.00198115 -0.000141964
+ 1.731e+11Hz -0.00196235 -0.000192414
+ 1.732e+11Hz -0.00194377 -0.000242788
+ 1.733e+11Hz -0.00192541 -0.000293084
+ 1.734e+11Hz -0.00190726 -0.000343302
+ 1.735e+11Hz -0.00188931 -0.000393441
+ 1.736e+11Hz -0.00187158 -0.000443501
+ 1.737e+11Hz -0.00185405 -0.00049348
+ 1.738e+11Hz -0.00183672 -0.000543378
+ 1.739e+11Hz -0.00181959 -0.000593195
+ 1.74e+11Hz -0.00180267 -0.00064293
+ 1.741e+11Hz -0.00178594 -0.000692582
+ 1.742e+11Hz -0.0017694 -0.000742152
+ 1.743e+11Hz -0.00175306 -0.000791638
+ 1.744e+11Hz -0.00173691 -0.00084104
+ 1.745e+11Hz -0.00172095 -0.000890358
+ 1.746e+11Hz -0.00170518 -0.000939592
+ 1.747e+11Hz -0.00168959 -0.000988741
+ 1.748e+11Hz -0.00167418 -0.0010378
+ 1.749e+11Hz -0.00165895 -0.00108678
+ 1.75e+11Hz -0.0016439 -0.00113568
+ 1.751e+11Hz -0.00162903 -0.00118448
+ 1.752e+11Hz -0.00161433 -0.00123321
+ 1.753e+11Hz -0.00159981 -0.00128184
+ 1.754e+11Hz -0.00158545 -0.00133039
+ 1.755e+11Hz -0.00157127 -0.00137885
+ 1.756e+11Hz -0.00155725 -0.00142723
+ 1.757e+11Hz -0.0015434 -0.00147552
+ 1.758e+11Hz -0.00152971 -0.00152373
+ 1.759e+11Hz -0.00151618 -0.00157185
+ 1.76e+11Hz -0.00150281 -0.00161988
+ 1.761e+11Hz -0.0014896 -0.00166783
+ 1.762e+11Hz -0.00147654 -0.00171569
+ 1.763e+11Hz -0.00146364 -0.00176347
+ 1.764e+11Hz -0.00145089 -0.00181116
+ 1.765e+11Hz -0.00143829 -0.00185876
+ 1.766e+11Hz -0.00142584 -0.00190628
+ 1.767e+11Hz -0.00141353 -0.00195372
+ 1.768e+11Hz -0.00140138 -0.00200107
+ 1.769e+11Hz -0.00138936 -0.00204833
+ 1.77e+11Hz -0.00137749 -0.00209551
+ 1.771e+11Hz -0.00136576 -0.00214261
+ 1.772e+11Hz -0.00135418 -0.00218962
+ 1.773e+11Hz -0.00134272 -0.00223655
+ 1.774e+11Hz -0.00133141 -0.0022834
+ 1.775e+11Hz -0.00132023 -0.00233017
+ 1.776e+11Hz -0.00130918 -0.00237685
+ 1.777e+11Hz -0.00129827 -0.00242345
+ 1.778e+11Hz -0.00128749 -0.00246996
+ 1.779e+11Hz -0.00127684 -0.0025164
+ 1.78e+11Hz -0.00126632 -0.00256276
+ 1.781e+11Hz -0.00125592 -0.00260903
+ 1.782e+11Hz -0.00124565 -0.00265522
+ 1.783e+11Hz -0.00123551 -0.00270133
+ 1.784e+11Hz -0.00122549 -0.00274736
+ 1.785e+11Hz -0.00121559 -0.00279332
+ 1.786e+11Hz -0.00120581 -0.00283919
+ 1.787e+11Hz -0.00119616 -0.00288498
+ 1.788e+11Hz -0.00118662 -0.00293069
+ 1.789e+11Hz -0.0011772 -0.00297633
+ 1.79e+11Hz -0.0011679 -0.00302188
+ 1.791e+11Hz -0.00115872 -0.00306736
+ 1.792e+11Hz -0.00114965 -0.00311276
+ 1.793e+11Hz -0.0011407 -0.00315807
+ 1.794e+11Hz -0.00113186 -0.00320332
+ 1.795e+11Hz -0.00112313 -0.00324848
+ 1.796e+11Hz -0.00111451 -0.00329356
+ 1.797e+11Hz -0.00110601 -0.00333857
+ 1.798e+11Hz -0.00109761 -0.0033835
+ 1.799e+11Hz -0.00108932 -0.00342835
+ 1.8e+11Hz -0.00108114 -0.00347312
+ 1.801e+11Hz -0.00107307 -0.00351782
+ 1.802e+11Hz -0.0010651 -0.00356244
+ 1.803e+11Hz -0.00105724 -0.00360697
+ 1.804e+11Hz -0.00104949 -0.00365144
+ 1.805e+11Hz -0.00104183 -0.00369582
+ 1.806e+11Hz -0.00103428 -0.00374012
+ 1.807e+11Hz -0.00102683 -0.00378435
+ 1.808e+11Hz -0.00101949 -0.00382849
+ 1.809e+11Hz -0.00101224 -0.00387256
+ 1.81e+11Hz -0.00100509 -0.00391655
+ 1.811e+11Hz -0.000998037 -0.00396045
+ 1.812e+11Hz -0.000991083 -0.00400428
+ 1.813e+11Hz -0.000984224 -0.00404803
+ 1.814e+11Hz -0.000977461 -0.00409169
+ 1.815e+11Hz -0.000970792 -0.00413528
+ 1.816e+11Hz -0.000964215 -0.00417878
+ 1.817e+11Hz -0.00095773 -0.0042222
+ 1.818e+11Hz -0.000951336 -0.00426554
+ 1.819e+11Hz -0.000945031 -0.00430879
+ 1.82e+11Hz -0.000938815 -0.00435196
+ 1.821e+11Hz -0.000932686 -0.00439505
+ 1.822e+11Hz -0.000926643 -0.00443805
+ 1.823e+11Hz -0.000920684 -0.00448097
+ 1.824e+11Hz -0.000914809 -0.0045238
+ 1.825e+11Hz -0.000909015 -0.00456654
+ 1.826e+11Hz -0.000903302 -0.00460919
+ 1.827e+11Hz -0.000897668 -0.00465176
+ 1.828e+11Hz -0.000892112 -0.00469424
+ 1.829e+11Hz -0.000886631 -0.00473663
+ 1.83e+11Hz -0.000881224 -0.00477893
+ 1.831e+11Hz -0.00087589 -0.00482113
+ 1.832e+11Hz -0.000870627 -0.00486325
+ 1.833e+11Hz -0.000865432 -0.00490527
+ 1.834e+11Hz -0.000860305 -0.0049472
+ 1.835e+11Hz -0.000855243 -0.00498904
+ 1.836e+11Hz -0.000850245 -0.00503078
+ 1.837e+11Hz -0.000845307 -0.00507243
+ 1.838e+11Hz -0.000840428 -0.00511398
+ 1.839e+11Hz -0.000835607 -0.00515544
+ 1.84e+11Hz -0.000830839 -0.0051968
+ 1.841e+11Hz -0.000826125 -0.00523806
+ 1.842e+11Hz -0.00082146 -0.00527922
+ 1.843e+11Hz -0.000816842 -0.00532029
+ 1.844e+11Hz -0.00081227 -0.00536125
+ 1.845e+11Hz -0.000807739 -0.00540212
+ 1.846e+11Hz -0.000803249 -0.00544288
+ 1.847e+11Hz -0.000798795 -0.00548355
+ 1.848e+11Hz -0.000794375 -0.00552411
+ 1.849e+11Hz -0.000789987 -0.00556457
+ 1.85e+11Hz -0.000785626 -0.00560493
+ 1.851e+11Hz -0.000781291 -0.00564519
+ 1.852e+11Hz -0.000776978 -0.00568534
+ 1.853e+11Hz -0.000772684 -0.0057254
+ 1.854e+11Hz -0.000768406 -0.00576535
+ 1.855e+11Hz -0.00076414 -0.0058052
+ 1.856e+11Hz -0.000759882 -0.00584495
+ 1.857e+11Hz -0.000755631 -0.00588459
+ 1.858e+11Hz -0.000751381 -0.00592414
+ 1.859e+11Hz -0.00074713 -0.00596358
+ 1.86e+11Hz -0.000742874 -0.00600292
+ 1.861e+11Hz -0.000738609 -0.00604216
+ 1.862e+11Hz -0.000734331 -0.0060813
+ 1.863e+11Hz -0.000730037 -0.00612034
+ 1.864e+11Hz -0.000725722 -0.00615929
+ 1.865e+11Hz -0.000721383 -0.00619813
+ 1.866e+11Hz -0.000717016 -0.00623688
+ 1.867e+11Hz -0.000712617 -0.00627554
+ 1.868e+11Hz -0.000708181 -0.0063141
+ 1.869e+11Hz -0.000703705 -0.00635256
+ 1.87e+11Hz -0.000699184 -0.00639094
+ 1.871e+11Hz -0.000694614 -0.00642923
+ 1.872e+11Hz -0.000689991 -0.00646742
+ 1.873e+11Hz -0.000685311 -0.00650554
+ 1.874e+11Hz -0.00068057 -0.00654356
+ 1.875e+11Hz -0.000675762 -0.00658151
+ 1.876e+11Hz -0.000670885 -0.00661938
+ 1.877e+11Hz -0.000665933 -0.00665717
+ 1.878e+11Hz -0.000660902 -0.00669488
+ 1.879e+11Hz -0.000655788 -0.00673252
+ 1.88e+11Hz -0.000650586 -0.0067701
+ 1.881e+11Hz -0.000645292 -0.0068076
+ 1.882e+11Hz -0.000639903 -0.00684505
+ 1.883e+11Hz -0.000634412 -0.00688243
+ 1.884e+11Hz -0.000628817 -0.00691976
+ 1.885e+11Hz -0.000623112 -0.00695703
+ 1.886e+11Hz -0.000617294 -0.00699426
+ 1.887e+11Hz -0.000611359 -0.00703144
+ 1.888e+11Hz -0.000605301 -0.00706858
+ 1.889e+11Hz -0.000599118 -0.00710568
+ 1.89e+11Hz -0.000592804 -0.00714275
+ 1.891e+11Hz -0.000586356 -0.0071798
+ 1.892e+11Hz -0.000579771 -0.00721682
+ 1.893e+11Hz -0.000573043 -0.00725382
+ 1.894e+11Hz -0.000566169 -0.00729081
+ 1.895e+11Hz -0.000559145 -0.00732779
+ 1.896e+11Hz -0.000551968 -0.00736477
+ 1.897e+11Hz -0.000544634 -0.00740175
+ 1.898e+11Hz -0.00053714 -0.00743875
+ 1.899e+11Hz -0.000529482 -0.00747575
+ 1.9e+11Hz -0.000521656 -0.00751278
+ 1.901e+11Hz -0.00051366 -0.00754984
+ 1.902e+11Hz -0.000505491 -0.00758693
+ 1.903e+11Hz -0.000497145 -0.00762406
+ 1.904e+11Hz -0.00048862 -0.00766123
+ 1.905e+11Hz -0.000479913 -0.00769846
+ 1.906e+11Hz -0.000471022 -0.00773576
+ 1.907e+11Hz -0.000461944 -0.00777312
+ 1.908e+11Hz -0.000452677 -0.00781055
+ 1.909e+11Hz -0.000443219 -0.00784807
+ 1.91e+11Hz -0.000433568 -0.00788568
+ 1.911e+11Hz -0.000423722 -0.00792339
+ 1.912e+11Hz -0.00041368 -0.0079612
+ 1.913e+11Hz -0.00040344 -0.00799913
+ 1.914e+11Hz -0.000393001 -0.00803718
+ 1.915e+11Hz -0.000382363 -0.00807536
+ 1.916e+11Hz -0.000371524 -0.00811367
+ 1.917e+11Hz -0.000360484 -0.00815214
+ 1.918e+11Hz -0.000349242 -0.00819076
+ 1.919e+11Hz -0.000337798 -0.00822955
+ 1.92e+11Hz -0.000326153 -0.00826851
+ 1.921e+11Hz -0.000314307 -0.00830765
+ 1.922e+11Hz -0.000302259 -0.00834698
+ 1.923e+11Hz -0.000290012 -0.00838651
+ 1.924e+11Hz -0.000277566 -0.00842625
+ 1.925e+11Hz -0.000264921 -0.00846622
+ 1.926e+11Hz -0.000252081 -0.0085064
+ 1.927e+11Hz -0.000239046 -0.00854683
+ 1.928e+11Hz -0.000225818 -0.0085875
+ 1.929e+11Hz -0.0002124 -0.00862843
+ 1.93e+11Hz -0.000198794 -0.00866962
+ 1.931e+11Hz -0.000185003 -0.00871109
+ 1.932e+11Hz -0.00017103 -0.00875284
+ 1.933e+11Hz -0.000156879 -0.00879488
+ 1.934e+11Hz -0.000142552 -0.00883723
+ 1.935e+11Hz -0.000128054 -0.00887989
+ 1.936e+11Hz -0.00011339 -0.00892287
+ 1.937e+11Hz -9.85621e-05 -0.00896618
+ 1.938e+11Hz -8.35767e-05 -0.00900983
+ 1.939e+11Hz -6.84385e-05 -0.00905384
+ 1.94e+11Hz -5.31526e-05 -0.0090982
+ 1.941e+11Hz -3.77246e-05 -0.00914293
+ 1.942e+11Hz -2.21604e-05 -0.00918804
+ 1.943e+11Hz -6.46614e-06 -0.00923354
+ 1.944e+11Hz 9.3518e-06 -0.00927943
+ 1.945e+11Hz 2.52867e-05 -0.00932573
+ 1.946e+11Hz 4.13316e-05 -0.00937244
+ 1.947e+11Hz 5.74792e-05 -0.00941958
+ 1.948e+11Hz 7.37219e-05 -0.00946714
+ 1.949e+11Hz 9.0052e-05 -0.00951515
+ 1.95e+11Hz 0.000106461 -0.0095636
+ 1.951e+11Hz 0.000122941 -0.00961251
+ 1.952e+11Hz 0.000139483 -0.00966189
+ 1.953e+11Hz 0.000156079 -0.00971174
+ 1.954e+11Hz 0.000172718 -0.00976207
+ 1.955e+11Hz 0.000189392 -0.00981289
+ 1.956e+11Hz 0.00020609 -0.0098642
+ 1.957e+11Hz 0.000222803 -0.00991602
+ 1.958e+11Hz 0.000239521 -0.00996835
+ 1.959e+11Hz 0.000256232 -0.0100212
+ 1.96e+11Hz 0.000272927 -0.0100746
+ 1.961e+11Hz 0.000289593 -0.0101285
+ 1.962e+11Hz 0.000306221 -0.0101829
+ 1.963e+11Hz 0.000322797 -0.0102379
+ 1.964e+11Hz 0.000339312 -0.0102934
+ 1.965e+11Hz 0.000355752 -0.0103495
+ 1.966e+11Hz 0.000372105 -0.0104061
+ 1.967e+11Hz 0.00038836 -0.0104633
+ 1.968e+11Hz 0.000404503 -0.0105211
+ 1.969e+11Hz 0.000420522 -0.0105794
+ 1.97e+11Hz 0.000436404 -0.0106383
+ 1.971e+11Hz 0.000452135 -0.0106978
+ 1.972e+11Hz 0.000467702 -0.0107579
+ 1.973e+11Hz 0.000483093 -0.0108186
+ 1.974e+11Hz 0.000498292 -0.0108798
+ 1.975e+11Hz 0.000513287 -0.0109417
+ 1.976e+11Hz 0.000528063 -0.0110041
+ 1.977e+11Hz 0.000542607 -0.0110672
+ 1.978e+11Hz 0.000556903 -0.0111308
+ 1.979e+11Hz 0.000570938 -0.011195
+ 1.98e+11Hz 0.000584697 -0.0112599
+ 1.981e+11Hz 0.000598166 -0.0113253
+ 1.982e+11Hz 0.000611331 -0.0113913
+ 1.983e+11Hz 0.000624175 -0.0114579
+ 1.984e+11Hz 0.000636685 -0.0115252
+ 1.985e+11Hz 0.000648846 -0.011593
+ 1.986e+11Hz 0.000660642 -0.0116614
+ 1.987e+11Hz 0.00067206 -0.0117304
+ 1.988e+11Hz 0.000683083 -0.0118
+ 1.989e+11Hz 0.000693697 -0.0118702
+ 1.99e+11Hz 0.000703887 -0.011941
+ 1.991e+11Hz 0.000713638 -0.0120124
+ 1.992e+11Hz 0.000722935 -0.0120843
+ 1.993e+11Hz 0.000731763 -0.0121569
+ 1.994e+11Hz 0.000740107 -0.01223
+ 1.995e+11Hz 0.000747952 -0.0123036
+ 1.996e+11Hz 0.000755283 -0.0123778
+ 1.997e+11Hz 0.000762086 -0.0124526
+ 1.998e+11Hz 0.000768346 -0.0125279
+ 1.999e+11Hz 0.000774049 -0.0126038
+ 2e+11Hz 0.000779179 -0.0126802
+ 2.001e+11Hz 0.000783722 -0.0127571
+ 2.002e+11Hz 0.000787665 -0.0128346
+ 2.003e+11Hz 0.000790993 -0.0129125
+ 2.004e+11Hz 0.000793692 -0.012991
+ 2.005e+11Hz 0.000795748 -0.01307
+ 2.006e+11Hz 0.000797148 -0.0131494
+ 2.007e+11Hz 0.000797878 -0.0132293
+ 2.008e+11Hz 0.000797925 -0.0133097
+ 2.009e+11Hz 0.000797276 -0.0133906
+ 2.01e+11Hz 0.000795917 -0.0134719
+ 2.011e+11Hz 0.000793837 -0.0135536
+ 2.012e+11Hz 0.000791023 -0.0136358
+ 2.013e+11Hz 0.000787462 -0.0137183
+ 2.014e+11Hz 0.000783143 -0.0138013
+ 2.015e+11Hz 0.000778053 -0.0138846
+ 2.016e+11Hz 0.000772183 -0.0139684
+ 2.017e+11Hz 0.000765519 -0.0140525
+ 2.018e+11Hz 0.000758052 -0.0141369
+ 2.019e+11Hz 0.000749772 -0.0142217
+ 2.02e+11Hz 0.000740666 -0.0143068
+ 2.021e+11Hz 0.000730727 -0.0143922
+ 2.022e+11Hz 0.000719944 -0.0144779
+ 2.023e+11Hz 0.000708307 -0.0145639
+ 2.024e+11Hz 0.000695809 -0.0146501
+ 2.025e+11Hz 0.00068244 -0.0147366
+ 2.026e+11Hz 0.000668192 -0.0148233
+ 2.027e+11Hz 0.000653057 -0.0149102
+ 2.028e+11Hz 0.000637027 -0.0149974
+ 2.029e+11Hz 0.000620096 -0.0150847
+ 2.03e+11Hz 0.000602257 -0.0151722
+ 2.031e+11Hz 0.000583503 -0.0152598
+ 2.032e+11Hz 0.000563829 -0.0153476
+ 2.033e+11Hz 0.000543228 -0.0154355
+ 2.034e+11Hz 0.000521696 -0.0155235
+ 2.035e+11Hz 0.000499228 -0.0156116
+ 2.036e+11Hz 0.000475819 -0.0156998
+ 2.037e+11Hz 0.000451465 -0.015788
+ 2.038e+11Hz 0.000426163 -0.0158762
+ 2.039e+11Hz 0.00039991 -0.0159645
+ 2.04e+11Hz 0.000372704 -0.0160527
+ 2.041e+11Hz 0.000344541 -0.0161409
+ 2.042e+11Hz 0.00031542 -0.0162291
+ 2.043e+11Hz 0.000285339 -0.0163172
+ 2.044e+11Hz 0.000254299 -0.0164053
+ 2.045e+11Hz 0.000222297 -0.0164933
+ 2.046e+11Hz 0.000189335 -0.0165811
+ 2.047e+11Hz 0.000155412 -0.0166689
+ 2.048e+11Hz 0.00012053 -0.0167564
+ 2.049e+11Hz 8.46886e-05 -0.0168438
+ 2.05e+11Hz 4.78907e-05 -0.0169311
+ 2.051e+11Hz 1.0138e-05 -0.0170181
+ 2.052e+11Hz -2.85667e-05 -0.0171049
+ 2.053e+11Hz -6.82207e-05 -0.0171915
+ 2.054e+11Hz -0.00010882 -0.0172778
+ 2.055e+11Hz -0.000150362 -0.0173638
+ 2.056e+11Hz -0.000192841 -0.0174496
+ 2.057e+11Hz -0.000236253 -0.0175351
+ 2.058e+11Hz -0.000280593 -0.0176202
+ 2.059e+11Hz -0.000325855 -0.017705
+ 2.06e+11Hz -0.000372033 -0.0177894
+ 2.061e+11Hz -0.000419121 -0.0178734
+ 2.062e+11Hz -0.000467112 -0.0179571
+ 2.063e+11Hz -0.000515999 -0.0180403
+ 2.064e+11Hz -0.000565774 -0.0181231
+ 2.065e+11Hz -0.00061643 -0.0182055
+ 2.066e+11Hz -0.000667958 -0.0182874
+ 2.067e+11Hz -0.000720348 -0.0183689
+ 2.068e+11Hz -0.000773593 -0.0184498
+ 2.069e+11Hz -0.000827683 -0.0185303
+ 2.07e+11Hz -0.000882607 -0.0186102
+ 2.071e+11Hz -0.000938356 -0.0186896
+ 2.072e+11Hz -0.000994919 -0.0187684
+ 2.073e+11Hz -0.00105229 -0.0188467
+ 2.074e+11Hz -0.00111044 -0.0189244
+ 2.075e+11Hz -0.00116938 -0.0190015
+ 2.076e+11Hz -0.00122909 -0.019078
+ 2.077e+11Hz -0.00128955 -0.0191539
+ 2.078e+11Hz -0.00135076 -0.0192291
+ 2.079e+11Hz -0.0014127 -0.0193038
+ 2.08e+11Hz -0.00147536 -0.0193777
+ 2.081e+11Hz -0.00153873 -0.019451
+ 2.082e+11Hz -0.00160278 -0.0195236
+ 2.083e+11Hz -0.00166752 -0.0195955
+ 2.084e+11Hz -0.00173291 -0.0196668
+ 2.085e+11Hz -0.00179896 -0.0197373
+ 2.086e+11Hz -0.00186565 -0.019807
+ 2.087e+11Hz -0.00193295 -0.0198761
+ 2.088e+11Hz -0.00200086 -0.0199444
+ 2.089e+11Hz -0.00206936 -0.020012
+ 2.09e+11Hz -0.00213844 -0.0200788
+ 2.091e+11Hz -0.00220808 -0.0201449
+ 2.092e+11Hz -0.00227827 -0.0202101
+ 2.093e+11Hz -0.00234898 -0.0202746
+ 2.094e+11Hz -0.00242021 -0.0203383
+ 2.095e+11Hz -0.00249194 -0.0204013
+ 2.096e+11Hz -0.00256415 -0.0204634
+ 2.097e+11Hz -0.00263683 -0.0205247
+ 2.098e+11Hz -0.00270995 -0.0205852
+ 2.099e+11Hz -0.00278352 -0.0206449
+ 2.1e+11Hz -0.0028575 -0.0207037
+ 2.101e+11Hz -0.00293188 -0.0207618
+ 2.102e+11Hz -0.00300665 -0.020819
+ 2.103e+11Hz -0.00308179 -0.0208754
+ 2.104e+11Hz -0.00315728 -0.020931
+ 2.105e+11Hz -0.00323311 -0.0209857
+ 2.106e+11Hz -0.00330926 -0.0210396
+ 2.107e+11Hz -0.00338571 -0.0210926
+ 2.108e+11Hz -0.00346246 -0.0211448
+ 2.109e+11Hz -0.00353947 -0.0211962
+ 2.11e+11Hz -0.00361674 -0.0212467
+ 2.111e+11Hz -0.00369426 -0.0212964
+ 2.112e+11Hz -0.00377199 -0.0213452
+ 2.113e+11Hz -0.00384994 -0.0213932
+ 2.114e+11Hz -0.00392807 -0.0214404
+ 2.115e+11Hz -0.00400639 -0.0214867
+ 2.116e+11Hz -0.00408487 -0.0215322
+ 2.117e+11Hz -0.00416349 -0.0215768
+ 2.118e+11Hz -0.00424224 -0.0216206
+ 2.119e+11Hz -0.00432111 -0.0216636
+ 2.12e+11Hz -0.00440008 -0.0217058
+ 2.121e+11Hz -0.00447914 -0.0217471
+ 2.122e+11Hz -0.00455827 -0.0217876
+ 2.123e+11Hz -0.00463745 -0.0218274
+ 2.124e+11Hz -0.00471668 -0.0218663
+ 2.125e+11Hz -0.00479594 -0.0219043
+ 2.126e+11Hz -0.00487521 -0.0219416
+ 2.127e+11Hz -0.00495448 -0.0219782
+ 2.128e+11Hz -0.00503375 -0.0220139
+ 2.129e+11Hz -0.00511298 -0.0220488
+ 2.13e+11Hz -0.00519218 -0.022083
+ 2.131e+11Hz -0.00527133 -0.0221163
+ 2.132e+11Hz -0.00535041 -0.022149
+ 2.133e+11Hz -0.00542942 -0.0221808
+ 2.134e+11Hz -0.00550835 -0.022212
+ 2.135e+11Hz -0.00558717 -0.0222424
+ 2.136e+11Hz -0.00566588 -0.022272
+ 2.137e+11Hz -0.00574447 -0.0223009
+ 2.138e+11Hz -0.00582293 -0.0223291
+ 2.139e+11Hz -0.00590124 -0.0223566
+ 2.14e+11Hz -0.0059794 -0.0223834
+ 2.141e+11Hz -0.0060574 -0.0224096
+ 2.142e+11Hz -0.00613523 -0.022435
+ 2.143e+11Hz -0.00621287 -0.0224597
+ 2.144e+11Hz -0.00629032 -0.0224838
+ 2.145e+11Hz -0.00636756 -0.0225073
+ 2.146e+11Hz -0.0064446 -0.0225301
+ 2.147e+11Hz -0.00652142 -0.0225522
+ 2.148e+11Hz -0.00659801 -0.0225737
+ 2.149e+11Hz -0.00667437 -0.0225947
+ 2.15e+11Hz -0.00675049 -0.022615
+ 2.151e+11Hz -0.00682636 -0.0226347
+ 2.152e+11Hz -0.00690198 -0.0226538
+ 2.153e+11Hz -0.00697733 -0.0226724
+ 2.154e+11Hz -0.00705241 -0.0226903
+ 2.155e+11Hz -0.00712722 -0.0227078
+ 2.156e+11Hz -0.00720175 -0.0227247
+ 2.157e+11Hz -0.007276 -0.022741
+ 2.158e+11Hz -0.00734995 -0.0227568
+ 2.159e+11Hz -0.00742361 -0.0227721
+ 2.16e+11Hz -0.00749697 -0.022787
+ 2.161e+11Hz -0.00757003 -0.0228013
+ 2.162e+11Hz -0.00764278 -0.0228151
+ 2.163e+11Hz -0.00771521 -0.0228285
+ 2.164e+11Hz -0.00778733 -0.0228413
+ 2.165e+11Hz -0.00785913 -0.0228538
+ 2.166e+11Hz -0.00793061 -0.0228658
+ 2.167e+11Hz -0.00800177 -0.0228774
+ 2.168e+11Hz -0.0080726 -0.0228885
+ 2.169e+11Hz -0.0081431 -0.0228992
+ 2.17e+11Hz -0.00821327 -0.0229096
+ 2.171e+11Hz -0.00828311 -0.0229195
+ 2.172e+11Hz -0.00835261 -0.0229291
+ 2.173e+11Hz -0.00842178 -0.0229383
+ 2.174e+11Hz -0.00849061 -0.0229471
+ 2.175e+11Hz -0.00855911 -0.0229556
+ 2.176e+11Hz -0.00862727 -0.0229637
+ 2.177e+11Hz -0.00869509 -0.0229715
+ 2.178e+11Hz -0.00876257 -0.022979
+ 2.179e+11Hz -0.00882972 -0.0229861
+ 2.18e+11Hz -0.00889653 -0.022993
+ 2.181e+11Hz -0.008963 -0.0229996
+ 2.182e+11Hz -0.00902914 -0.0230058
+ 2.183e+11Hz -0.00909494 -0.0230118
+ 2.184e+11Hz -0.0091604 -0.0230175
+ 2.185e+11Hz -0.00922553 -0.023023
+ 2.186e+11Hz -0.00929033 -0.0230282
+ 2.187e+11Hz -0.0093548 -0.0230332
+ 2.188e+11Hz -0.00941894 -0.0230379
+ 2.189e+11Hz -0.00948276 -0.0230424
+ 2.19e+11Hz -0.00954625 -0.0230467
+ 2.191e+11Hz -0.00960941 -0.0230507
+ 2.192e+11Hz -0.00967225 -0.0230546
+ 2.193e+11Hz -0.00973478 -0.0230583
+ 2.194e+11Hz -0.00979699 -0.0230617
+ 2.195e+11Hz -0.00985888 -0.023065
+ 2.196e+11Hz -0.00992046 -0.0230682
+ 2.197e+11Hz -0.00998173 -0.0230711
+ 2.198e+11Hz -0.0100427 -0.0230739
+ 2.199e+11Hz -0.0101034 -0.0230765
+ 2.2e+11Hz -0.0101637 -0.023079
+ 2.201e+11Hz -0.0102238 -0.0230813
+ 2.202e+11Hz -0.0102836 -0.0230835
+ 2.203e+11Hz -0.010343 -0.0230856
+ 2.204e+11Hz -0.0104022 -0.0230876
+ 2.205e+11Hz -0.0104612 -0.0230894
+ 2.206e+11Hz -0.0105198 -0.0230911
+ 2.207e+11Hz -0.0105781 -0.0230927
+ 2.208e+11Hz -0.0106362 -0.0230943
+ 2.209e+11Hz -0.010694 -0.0230957
+ 2.21e+11Hz -0.0107516 -0.023097
+ 2.211e+11Hz -0.0108088 -0.0230982
+ 2.212e+11Hz -0.0108658 -0.0230994
+ 2.213e+11Hz -0.0109226 -0.0231005
+ 2.214e+11Hz -0.0109791 -0.0231015
+ 2.215e+11Hz -0.0110354 -0.0231025
+ 2.216e+11Hz -0.0110914 -0.0231034
+ 2.217e+11Hz -0.0111471 -0.0231042
+ 2.218e+11Hz -0.0112027 -0.023105
+ 2.219e+11Hz -0.011258 -0.0231057
+ 2.22e+11Hz -0.011313 -0.0231064
+ 2.221e+11Hz -0.0113679 -0.0231071
+ 2.222e+11Hz -0.0114225 -0.0231077
+ 2.223e+11Hz -0.0114769 -0.0231083
+ 2.224e+11Hz -0.0115311 -0.0231089
+ 2.225e+11Hz -0.011585 -0.0231094
+ 2.226e+11Hz -0.0116388 -0.0231099
+ 2.227e+11Hz -0.0116923 -0.0231104
+ 2.228e+11Hz -0.0117457 -0.0231109
+ 2.229e+11Hz -0.0117989 -0.0231114
+ 2.23e+11Hz -0.0118518 -0.0231119
+ 2.231e+11Hz -0.0119046 -0.0231124
+ 2.232e+11Hz -0.0119572 -0.0231129
+ 2.233e+11Hz -0.0120096 -0.0231134
+ 2.234e+11Hz -0.0120619 -0.0231139
+ 2.235e+11Hz -0.0121139 -0.0231144
+ 2.236e+11Hz -0.0121658 -0.0231149
+ 2.237e+11Hz -0.0122175 -0.0231155
+ 2.238e+11Hz -0.0122691 -0.0231161
+ 2.239e+11Hz -0.0123205 -0.0231167
+ 2.24e+11Hz -0.0123718 -0.0231173
+ 2.241e+11Hz -0.0124229 -0.023118
+ 2.242e+11Hz -0.0124738 -0.0231187
+ 2.243e+11Hz -0.0125246 -0.0231194
+ 2.244e+11Hz -0.0125753 -0.0231202
+ 2.245e+11Hz -0.0126259 -0.023121
+ 2.246e+11Hz -0.0126763 -0.0231218
+ 2.247e+11Hz -0.0127266 -0.0231228
+ 2.248e+11Hz -0.0127767 -0.0231237
+ 2.249e+11Hz -0.0128268 -0.0231247
+ 2.25e+11Hz -0.0128767 -0.0231258
+ 2.251e+11Hz -0.0129266 -0.023127
+ 2.252e+11Hz -0.0129763 -0.0231282
+ 2.253e+11Hz -0.0130259 -0.0231295
+ 2.254e+11Hz -0.0130755 -0.0231308
+ 2.255e+11Hz -0.0131249 -0.0231322
+ 2.256e+11Hz -0.0131743 -0.0231337
+ 2.257e+11Hz -0.0132235 -0.0231353
+ 2.258e+11Hz -0.0132727 -0.0231369
+ 2.259e+11Hz -0.0133219 -0.0231387
+ 2.26e+11Hz -0.0133709 -0.0231405
+ 2.261e+11Hz -0.0134199 -0.0231424
+ 2.262e+11Hz -0.0134689 -0.0231444
+ 2.263e+11Hz -0.0135178 -0.0231465
+ 2.264e+11Hz -0.0135666 -0.0231487
+ 2.265e+11Hz -0.0136154 -0.023151
+ 2.266e+11Hz -0.0136642 -0.0231534
+ 2.267e+11Hz -0.0137129 -0.0231559
+ 2.268e+11Hz -0.0137617 -0.0231585
+ 2.269e+11Hz -0.0138104 -0.0231612
+ 2.27e+11Hz -0.013859 -0.023164
+ 2.271e+11Hz -0.0139077 -0.0231669
+ 2.272e+11Hz -0.0139564 -0.02317
+ 2.273e+11Hz -0.0140051 -0.0231731
+ 2.274e+11Hz -0.0140538 -0.0231764
+ 2.275e+11Hz -0.0141025 -0.0231798
+ 2.276e+11Hz -0.0141512 -0.0231833
+ 2.277e+11Hz -0.0142 -0.023187
+ 2.278e+11Hz -0.0142488 -0.0231908
+ 2.279e+11Hz -0.0142977 -0.0231947
+ 2.28e+11Hz -0.0143466 -0.0231987
+ 2.281e+11Hz -0.0143955 -0.0232028
+ 2.282e+11Hz -0.0144446 -0.0232071
+ 2.283e+11Hz -0.0144937 -0.0232115
+ 2.284e+11Hz -0.0145429 -0.0232161
+ 2.285e+11Hz -0.0145921 -0.0232208
+ 2.286e+11Hz -0.0146415 -0.0232256
+ 2.287e+11Hz -0.014691 -0.0232305
+ 2.288e+11Hz -0.0147406 -0.0232356
+ 2.289e+11Hz -0.0147903 -0.0232409
+ 2.29e+11Hz -0.0148401 -0.0232462
+ 2.291e+11Hz -0.0148901 -0.0232517
+ 2.292e+11Hz -0.0149402 -0.0232573
+ 2.293e+11Hz -0.0149905 -0.0232631
+ 2.294e+11Hz -0.0150409 -0.023269
+ 2.295e+11Hz -0.0150915 -0.023275
+ 2.296e+11Hz -0.0151423 -0.0232812
+ 2.297e+11Hz -0.0151933 -0.0232874
+ 2.298e+11Hz -0.0152445 -0.0232938
+ 2.299e+11Hz -0.0152959 -0.0233004
+ 2.3e+11Hz -0.0153475 -0.023307
+ 2.301e+11Hz -0.0153993 -0.0233138
+ 2.302e+11Hz -0.0154513 -0.0233207
+ 2.303e+11Hz -0.0155036 -0.0233277
+ 2.304e+11Hz -0.0155562 -0.0233349
+ 2.305e+11Hz -0.015609 -0.0233421
+ 2.306e+11Hz -0.0156621 -0.0233495
+ 2.307e+11Hz -0.0157155 -0.0233569
+ 2.308e+11Hz -0.0157691 -0.0233645
+ 2.309e+11Hz -0.0158231 -0.0233721
+ 2.31e+11Hz -0.0158774 -0.0233798
+ 2.311e+11Hz -0.015932 -0.0233876
+ 2.312e+11Hz -0.0159869 -0.0233955
+ 2.313e+11Hz -0.0160422 -0.0234035
+ 2.314e+11Hz -0.0160978 -0.0234115
+ 2.315e+11Hz -0.0161538 -0.0234196
+ 2.316e+11Hz -0.0162101 -0.0234278
+ 2.317e+11Hz -0.0162668 -0.023436
+ 2.318e+11Hz -0.0163239 -0.0234442
+ 2.319e+11Hz -0.0163815 -0.0234525
+ 2.32e+11Hz -0.0164394 -0.0234608
+ 2.321e+11Hz -0.0164977 -0.0234691
+ 2.322e+11Hz -0.0165565 -0.0234775
+ 2.323e+11Hz -0.0166157 -0.0234858
+ 2.324e+11Hz -0.0166753 -0.0234941
+ 2.325e+11Hz -0.0167354 -0.0235024
+ 2.326e+11Hz -0.016796 -0.0235107
+ 2.327e+11Hz -0.016857 -0.0235189
+ 2.328e+11Hz -0.0169185 -0.0235271
+ 2.329e+11Hz -0.0169805 -0.0235352
+ 2.33e+11Hz -0.017043 -0.0235433
+ 2.331e+11Hz -0.0171059 -0.0235512
+ 2.332e+11Hz -0.0171694 -0.0235591
+ 2.333e+11Hz -0.0172335 -0.0235669
+ 2.334e+11Hz -0.017298 -0.0235746
+ 2.335e+11Hz -0.0173631 -0.0235821
+ 2.336e+11Hz -0.0174287 -0.0235895
+ 2.337e+11Hz -0.0174949 -0.0235967
+ 2.338e+11Hz -0.0175616 -0.0236038
+ 2.339e+11Hz -0.0176288 -0.0236106
+ 2.34e+11Hz -0.0176967 -0.0236173
+ 2.341e+11Hz -0.0177651 -0.0236237
+ 2.342e+11Hz -0.0178341 -0.02363
+ 2.343e+11Hz -0.0179036 -0.023636
+ 2.344e+11Hz -0.0179738 -0.0236417
+ 2.345e+11Hz -0.0180445 -0.0236471
+ 2.346e+11Hz -0.0181158 -0.0236523
+ 2.347e+11Hz -0.0181878 -0.0236571
+ 2.348e+11Hz -0.0182603 -0.0236617
+ 2.349e+11Hz -0.0183334 -0.0236658
+ 2.35e+11Hz -0.0184071 -0.0236697
+ 2.351e+11Hz -0.0184814 -0.0236731
+ 2.352e+11Hz -0.0185564 -0.0236762
+ 2.353e+11Hz -0.0186319 -0.0236788
+ 2.354e+11Hz -0.0187081 -0.0236811
+ 2.355e+11Hz -0.0187848 -0.0236828
+ 2.356e+11Hz -0.0188622 -0.0236842
+ 2.357e+11Hz -0.0189402 -0.023685
+ 2.358e+11Hz -0.0190187 -0.0236853
+ 2.359e+11Hz -0.0190979 -0.0236851
+ 2.36e+11Hz -0.0191777 -0.0236844
+ 2.361e+11Hz -0.0192581 -0.0236831
+ 2.362e+11Hz -0.019339 -0.0236813
+ 2.363e+11Hz -0.0194206 -0.0236788
+ 2.364e+11Hz -0.0195027 -0.0236757
+ 2.365e+11Hz -0.0195855 -0.023672
+ 2.366e+11Hz -0.0196688 -0.0236677
+ 2.367e+11Hz -0.0197527 -0.0236627
+ 2.368e+11Hz -0.0198371 -0.0236569
+ 2.369e+11Hz -0.0199221 -0.0236505
+ 2.37e+11Hz -0.0200076 -0.0236434
+ 2.371e+11Hz -0.0200937 -0.0236355
+ 2.372e+11Hz -0.0201803 -0.0236268
+ 2.373e+11Hz -0.0202675 -0.0236174
+ 2.374e+11Hz -0.0203551 -0.0236071
+ 2.375e+11Hz -0.0204433 -0.023596
+ 2.376e+11Hz -0.0205319 -0.0235841
+ 2.377e+11Hz -0.020621 -0.0235713
+ 2.378e+11Hz -0.0207106 -0.0235577
+ 2.379e+11Hz -0.0208007 -0.0235431
+ 2.38e+11Hz -0.0208911 -0.0235276
+ 2.381e+11Hz -0.0209821 -0.0235112
+ 2.382e+11Hz -0.0210734 -0.0234939
+ 2.383e+11Hz -0.0211651 -0.0234756
+ 2.384e+11Hz -0.0212572 -0.0234563
+ 2.385e+11Hz -0.0213497 -0.023436
+ 2.386e+11Hz -0.0214425 -0.0234146
+ 2.387e+11Hz -0.0215357 -0.0233923
+ 2.388e+11Hz -0.0216291 -0.0233689
+ 2.389e+11Hz -0.0217229 -0.0233444
+ 2.39e+11Hz -0.021817 -0.0233188
+ 2.391e+11Hz -0.0219113 -0.0232922
+ 2.392e+11Hz -0.0220058 -0.0232644
+ 2.393e+11Hz -0.0221006 -0.0232356
+ 2.394e+11Hz -0.0221956 -0.0232055
+ 2.395e+11Hz -0.0222907 -0.0231744
+ 2.396e+11Hz -0.022386 -0.023142
+ 2.397e+11Hz -0.0224814 -0.0231085
+ 2.398e+11Hz -0.022577 -0.0230739
+ 2.399e+11Hz -0.0226726 -0.023038
+ 2.4e+11Hz -0.0227683 -0.0230009
+ 2.401e+11Hz -0.0228641 -0.0229626
+ 2.402e+11Hz -0.0229598 -0.022923
+ 2.403e+11Hz -0.0230556 -0.0228823
+ 2.404e+11Hz -0.0231513 -0.0228402
+ 2.405e+11Hz -0.023247 -0.022797
+ 2.406e+11Hz -0.0233426 -0.0227524
+ 2.407e+11Hz -0.0234381 -0.0227066
+ 2.408e+11Hz -0.0235334 -0.0226596
+ 2.409e+11Hz -0.0236286 -0.0226112
+ 2.41e+11Hz -0.0237236 -0.0225616
+ 2.411e+11Hz -0.0238184 -0.0225107
+ 2.412e+11Hz -0.0239129 -0.0224585
+ 2.413e+11Hz -0.0240072 -0.022405
+ 2.414e+11Hz -0.0241012 -0.0223502
+ 2.415e+11Hz -0.0241948 -0.0222941
+ 2.416e+11Hz -0.0242881 -0.0222367
+ 2.417e+11Hz -0.0243811 -0.0221781
+ 2.418e+11Hz -0.0244736 -0.0221181
+ 2.419e+11Hz -0.0245657 -0.0220568
+ 2.42e+11Hz -0.0246573 -0.0219943
+ 2.421e+11Hz -0.0247484 -0.0219305
+ 2.422e+11Hz -0.024839 -0.0218653
+ 2.423e+11Hz -0.0249291 -0.0217989
+ 2.424e+11Hz -0.0250185 -0.0217313
+ 2.425e+11Hz -0.0251074 -0.0216623
+ 2.426e+11Hz -0.0251956 -0.0215921
+ 2.427e+11Hz -0.0252832 -0.0215207
+ 2.428e+11Hz -0.0253701 -0.021448
+ 2.429e+11Hz -0.0254562 -0.021374
+ 2.43e+11Hz -0.0255416 -0.0212989
+ 2.431e+11Hz -0.0256263 -0.0212225
+ 2.432e+11Hz -0.0257101 -0.0211449
+ 2.433e+11Hz -0.0257931 -0.0210662
+ 2.434e+11Hz -0.0258753 -0.0209862
+ 2.435e+11Hz -0.0259565 -0.0209051
+ 2.436e+11Hz -0.0260369 -0.0208228
+ 2.437e+11Hz -0.0261163 -0.0207394
+ 2.438e+11Hz -0.0261947 -0.0206549
+ 2.439e+11Hz -0.0262722 -0.0205693
+ 2.44e+11Hz -0.0263486 -0.0204826
+ 2.441e+11Hz -0.026424 -0.0203948
+ 2.442e+11Hz -0.0264984 -0.0203059
+ 2.443e+11Hz -0.0265716 -0.0202161
+ 2.444e+11Hz -0.0266438 -0.0201252
+ 2.445e+11Hz -0.0267148 -0.0200333
+ 2.446e+11Hz -0.0267846 -0.0199405
+ 2.447e+11Hz -0.0268533 -0.0198467
+ 2.448e+11Hz -0.0269207 -0.019752
+ 2.449e+11Hz -0.026987 -0.0196564
+ 2.45e+11Hz -0.0270519 -0.0195599
+ 2.451e+11Hz -0.0271157 -0.0194625
+ 2.452e+11Hz -0.0271781 -0.0193643
+ 2.453e+11Hz -0.0272392 -0.0192653
+ 2.454e+11Hz -0.0272991 -0.0191656
+ 2.455e+11Hz -0.0273575 -0.019065
+ 2.456e+11Hz -0.0274146 -0.0189638
+ 2.457e+11Hz -0.0274704 -0.0188618
+ 2.458e+11Hz -0.0275247 -0.0187592
+ 2.459e+11Hz -0.0275777 -0.0186559
+ 2.46e+11Hz -0.0276292 -0.018552
+ 2.461e+11Hz -0.0276793 -0.0184476
+ 2.462e+11Hz -0.0277279 -0.0183426
+ 2.463e+11Hz -0.0277751 -0.018237
+ 2.464e+11Hz -0.0278209 -0.018131
+ 2.465e+11Hz -0.0278651 -0.0180244
+ 2.466e+11Hz -0.0279078 -0.0179175
+ 2.467e+11Hz -0.0279491 -0.0178101
+ 2.468e+11Hz -0.0279888 -0.0177024
+ 2.469e+11Hz -0.028027 -0.0175943
+ 2.47e+11Hz -0.0280637 -0.0174859
+ 2.471e+11Hz -0.0280989 -0.0173773
+ 2.472e+11Hz -0.0281326 -0.0172683
+ 2.473e+11Hz -0.0281647 -0.0171592
+ 2.474e+11Hz -0.0281952 -0.0170499
+ 2.475e+11Hz -0.0282242 -0.0169404
+ 2.476e+11Hz -0.0282517 -0.0168309
+ 2.477e+11Hz -0.0282776 -0.0167212
+ 2.478e+11Hz -0.028302 -0.0166115
+ 2.479e+11Hz -0.0283248 -0.0165017
+ 2.48e+11Hz -0.0283461 -0.016392
+ 2.481e+11Hz -0.0283658 -0.0162823
+ 2.482e+11Hz -0.028384 -0.0161727
+ 2.483e+11Hz -0.0284007 -0.0160632
+ 2.484e+11Hz -0.0284158 -0.0159539
+ 2.485e+11Hz -0.0284294 -0.0158447
+ 2.486e+11Hz -0.0284415 -0.0157357
+ 2.487e+11Hz -0.028452 -0.015627
+ 2.488e+11Hz -0.0284611 -0.0155185
+ 2.489e+11Hz -0.0284687 -0.0154103
+ 2.49e+11Hz -0.0284748 -0.0153025
+ 2.491e+11Hz -0.0284794 -0.015195
+ 2.492e+11Hz -0.0284825 -0.0150879
+ 2.493e+11Hz -0.0284842 -0.0149812
+ 2.494e+11Hz -0.0284845 -0.014875
+ 2.495e+11Hz -0.0284833 -0.0147692
+ 2.496e+11Hz -0.0284807 -0.014664
+ 2.497e+11Hz -0.0284767 -0.0145593
+ 2.498e+11Hz -0.0284714 -0.0144551
+ 2.499e+11Hz -0.0284646 -0.0143516
+ 2.5e+11Hz -0.0284566 -0.0142487
+ 2.501e+11Hz -0.0284471 -0.0141464
+ 2.502e+11Hz -0.0284364 -0.0140448
+ 2.503e+11Hz -0.0284244 -0.0139439
+ 2.504e+11Hz -0.0284111 -0.0138437
+ 2.505e+11Hz -0.0283966 -0.0137442
+ 2.506e+11Hz -0.0283808 -0.0136456
+ 2.507e+11Hz -0.0283638 -0.0135477
+ 2.508e+11Hz -0.0283457 -0.0134506
+ 2.509e+11Hz -0.0283264 -0.0133544
+ 2.51e+11Hz -0.0283059 -0.013259
+ 2.511e+11Hz -0.0282843 -0.0131646
+ 2.512e+11Hz -0.0282616 -0.013071
+ 2.513e+11Hz -0.0282378 -0.0129783
+ 2.514e+11Hz -0.028213 -0.0128866
+ 2.515e+11Hz -0.0281872 -0.0127958
+ 2.516e+11Hz -0.0281604 -0.0127061
+ 2.517e+11Hz -0.0281326 -0.0126173
+ 2.518e+11Hz -0.0281038 -0.0125295
+ 2.519e+11Hz -0.0280742 -0.0124427
+ 2.52e+11Hz -0.0280437 -0.012357
+ 2.521e+11Hz -0.0280123 -0.0122723
+ 2.522e+11Hz -0.02798 -0.0121887
+ 2.523e+11Hz -0.027947 -0.0121061
+ 2.524e+11Hz -0.0279132 -0.0120247
+ 2.525e+11Hz -0.0278786 -0.0119443
+ 2.526e+11Hz -0.0278433 -0.011865
+ 2.527e+11Hz -0.0278074 -0.0117869
+ 2.528e+11Hz -0.0277707 -0.0117099
+ 2.529e+11Hz -0.0277335 -0.011634
+ 2.53e+11Hz -0.0276956 -0.0115592
+ 2.531e+11Hz -0.0276571 -0.0114856
+ 2.532e+11Hz -0.0276181 -0.0114131
+ 2.533e+11Hz -0.0275786 -0.0113418
+ 2.534e+11Hz -0.0275386 -0.0112716
+ 2.535e+11Hz -0.0274981 -0.0112026
+ 2.536e+11Hz -0.0274572 -0.0111348
+ 2.537e+11Hz -0.0274159 -0.0110681
+ 2.538e+11Hz -0.0273743 -0.0110025
+ 2.539e+11Hz -0.0273322 -0.0109382
+ 2.54e+11Hz -0.0272899 -0.0108749
+ 2.541e+11Hz -0.0272473 -0.0108129
+ 2.542e+11Hz -0.0272044 -0.010752
+ 2.543e+11Hz -0.0271613 -0.0106922
+ 2.544e+11Hz -0.027118 -0.0106336
+ 2.545e+11Hz -0.0270745 -0.0105761
+ 2.546e+11Hz -0.0270308 -0.0105197
+ 2.547e+11Hz -0.026987 -0.0104645
+ 2.548e+11Hz -0.0269432 -0.0104104
+ 2.549e+11Hz -0.0268992 -0.0103574
+ 2.55e+11Hz -0.0268552 -0.0103055
+ 2.551e+11Hz -0.0268112 -0.0102547
+ 2.552e+11Hz -0.0267672 -0.0102049
+ 2.553e+11Hz -0.0267232 -0.0101563
+ 2.554e+11Hz -0.0266793 -0.0101087
+ 2.555e+11Hz -0.0266355 -0.0100621
+ 2.556e+11Hz -0.0265917 -0.0100166
+ 2.557e+11Hz -0.0265481 -0.00997215
+ 2.558e+11Hz -0.0265046 -0.00992867
+ 2.559e+11Hz -0.0264613 -0.00988619
+ 2.56e+11Hz -0.0264181 -0.0098447
+ 2.561e+11Hz -0.0263752 -0.00980417
+ 2.562e+11Hz -0.0263325 -0.00976459
+ 2.563e+11Hz -0.0262901 -0.00972594
+ 2.564e+11Hz -0.0262479 -0.00968822
+ 2.565e+11Hz -0.026206 -0.00965139
+ 2.566e+11Hz -0.0261644 -0.00961545
+ 2.567e+11Hz -0.0261231 -0.00958038
+ 2.568e+11Hz -0.0260821 -0.00954616
+ 2.569e+11Hz -0.0260415 -0.00951276
+ 2.57e+11Hz -0.0260013 -0.00948019
+ 2.571e+11Hz -0.0259614 -0.0094484
+ 2.572e+11Hz -0.025922 -0.00941739
+ 2.573e+11Hz -0.0258829 -0.00938713
+ 2.574e+11Hz -0.0258443 -0.00935761
+ 2.575e+11Hz -0.0258061 -0.00932881
+ 2.576e+11Hz -0.0257683 -0.0093007
+ 2.577e+11Hz -0.025731 -0.00927327
+ 2.578e+11Hz -0.0256941 -0.00924649
+ 2.579e+11Hz -0.0256578 -0.00922035
+ 2.58e+11Hz -0.0256219 -0.00919482
+ 2.581e+11Hz -0.0255865 -0.00916988
+ 2.582e+11Hz -0.0255515 -0.00914552
+ 2.583e+11Hz -0.0255171 -0.00912171
+ 2.584e+11Hz -0.0254832 -0.00909844
+ 2.585e+11Hz -0.0254498 -0.00907567
+ 2.586e+11Hz -0.0254169 -0.0090534
+ 2.587e+11Hz -0.0253846 -0.00903159
+ 2.588e+11Hz -0.0253527 -0.00901024
+ 2.589e+11Hz -0.0253214 -0.00898931
+ 2.59e+11Hz -0.0252906 -0.0089688
+ 2.591e+11Hz -0.0252603 -0.00894867
+ 2.592e+11Hz -0.0252306 -0.00892891
+ 2.593e+11Hz -0.0252014 -0.00890951
+ 2.594e+11Hz -0.0251727 -0.00889043
+ 2.595e+11Hz -0.0251446 -0.00887166
+ 2.596e+11Hz -0.0251169 -0.00885318
+ 2.597e+11Hz -0.0250898 -0.00883498
+ 2.598e+11Hz -0.0250632 -0.00881703
+ 2.599e+11Hz -0.0250372 -0.00879931
+ 2.6e+11Hz -0.0250116 -0.00878181
+ 2.601e+11Hz -0.0249865 -0.00876452
+ 2.602e+11Hz -0.024962 -0.0087474
+ 2.603e+11Hz -0.0249379 -0.00873045
+ 2.604e+11Hz -0.0249144 -0.00871365
+ 2.605e+11Hz -0.0248913 -0.00869698
+ 2.606e+11Hz -0.0248687 -0.00868043
+ 2.607e+11Hz -0.0248465 -0.00866398
+ 2.608e+11Hz -0.0248248 -0.00864761
+ 2.609e+11Hz -0.0248036 -0.00863132
+ 2.61e+11Hz -0.0247828 -0.00861508
+ 2.611e+11Hz -0.0247624 -0.00859889
+ 2.612e+11Hz -0.0247425 -0.00858273
+ 2.613e+11Hz -0.024723 -0.00856659
+ 2.614e+11Hz -0.0247039 -0.00855045
+ 2.615e+11Hz -0.0246852 -0.00853431
+ 2.616e+11Hz -0.0246668 -0.00851815
+ 2.617e+11Hz -0.0246488 -0.00850197
+ 2.618e+11Hz -0.0246312 -0.00848574
+ 2.619e+11Hz -0.024614 -0.00846947
+ 2.62e+11Hz -0.0245971 -0.00845314
+ 2.621e+11Hz -0.0245805 -0.00843674
+ 2.622e+11Hz -0.0245642 -0.00842027
+ 2.623e+11Hz -0.0245482 -0.00840372
+ 2.624e+11Hz -0.0245325 -0.00838708
+ 2.625e+11Hz -0.0245171 -0.00837035
+ 2.626e+11Hz -0.0245019 -0.00835352
+ 2.627e+11Hz -0.024487 -0.00833658
+ 2.628e+11Hz -0.0244723 -0.00831953
+ 2.629e+11Hz -0.0244579 -0.00830236
+ 2.63e+11Hz -0.0244437 -0.00828508
+ 2.631e+11Hz -0.0244296 -0.00826767
+ 2.632e+11Hz -0.0244158 -0.00825014
+ 2.633e+11Hz -0.0244021 -0.00823248
+ 2.634e+11Hz -0.0243886 -0.00821469
+ 2.635e+11Hz -0.0243753 -0.00819678
+ 2.636e+11Hz -0.024362 -0.00817873
+ 2.637e+11Hz -0.0243489 -0.00816056
+ 2.638e+11Hz -0.024336 -0.00814225
+ 2.639e+11Hz -0.0243231 -0.00812382
+ 2.64e+11Hz -0.0243103 -0.00810526
+ 2.641e+11Hz -0.0242976 -0.00808657
+ 2.642e+11Hz -0.0242849 -0.00806776
+ 2.643e+11Hz -0.0242723 -0.00804883
+ 2.644e+11Hz -0.0242598 -0.00802979
+ 2.645e+11Hz -0.0242473 -0.00801063
+ 2.646e+11Hz -0.0242348 -0.00799136
+ 2.647e+11Hz -0.0242223 -0.00797199
+ 2.648e+11Hz -0.0242098 -0.00795252
+ 2.649e+11Hz -0.0241973 -0.00793296
+ 2.65e+11Hz -0.0241848 -0.00791331
+ 2.651e+11Hz -0.0241723 -0.00789357
+ 2.652e+11Hz -0.0241597 -0.00787377
+ 2.653e+11Hz -0.0241471 -0.00785389
+ 2.654e+11Hz -0.0241345 -0.00783395
+ 2.655e+11Hz -0.0241218 -0.00781396
+ 2.656e+11Hz -0.024109 -0.00779393
+ 2.657e+11Hz -0.0240961 -0.00777385
+ 2.658e+11Hz -0.0240832 -0.00775375
+ 2.659e+11Hz -0.0240702 -0.00773363
+ 2.66e+11Hz -0.0240571 -0.00771349
+ 2.661e+11Hz -0.024044 -0.00769335
+ 2.662e+11Hz -0.0240307 -0.00767322
+ 2.663e+11Hz -0.0240173 -0.00765311
+ 2.664e+11Hz -0.0240038 -0.00763302
+ 2.665e+11Hz -0.0239903 -0.00761296
+ 2.666e+11Hz -0.0239766 -0.00759295
+ 2.667e+11Hz -0.0239628 -0.007573
+ 2.668e+11Hz -0.0239488 -0.00755311
+ 2.669e+11Hz -0.0239348 -0.0075333
+ 2.67e+11Hz -0.0239207 -0.00751357
+ 2.671e+11Hz -0.0239064 -0.00749394
+ 2.672e+11Hz -0.0238921 -0.00747442
+ 2.673e+11Hz -0.0238776 -0.00745501
+ 2.674e+11Hz -0.023863 -0.00743573
+ 2.675e+11Hz -0.0238483 -0.00741658
+ 2.676e+11Hz -0.0238335 -0.00739758
+ 2.677e+11Hz -0.0238186 -0.00737874
+ 2.678e+11Hz -0.0238035 -0.00736007
+ 2.679e+11Hz -0.0237884 -0.00734157
+ 2.68e+11Hz -0.0237732 -0.00732326
+ 2.681e+11Hz -0.0237579 -0.00730515
+ 2.682e+11Hz -0.0237426 -0.00728724
+ 2.683e+11Hz -0.0237271 -0.00726955
+ 2.684e+11Hz -0.0237116 -0.00725208
+ 2.685e+11Hz -0.023696 -0.00723484
+ 2.686e+11Hz -0.0236804 -0.00721785
+ 2.687e+11Hz -0.0236647 -0.00720111
+ 2.688e+11Hz -0.0236489 -0.00718462
+ 2.689e+11Hz -0.0236332 -0.0071684
+ 2.69e+11Hz -0.0236174 -0.00715246
+ 2.691e+11Hz -0.0236016 -0.00713679
+ 2.692e+11Hz -0.0235857 -0.00712141
+ 2.693e+11Hz -0.0235699 -0.00710633
+ 2.694e+11Hz -0.0235541 -0.00709155
+ 2.695e+11Hz -0.0235383 -0.00707708
+ 2.696e+11Hz -0.0235226 -0.00706291
+ 2.697e+11Hz -0.0235069 -0.00704907
+ 2.698e+11Hz -0.0234913 -0.00703555
+ 2.699e+11Hz -0.0234757 -0.00702235
+ 2.7e+11Hz -0.0234602 -0.00700949
+ 2.701e+11Hz -0.0234448 -0.00699695
+ 2.702e+11Hz -0.0234295 -0.00698476
+ 2.703e+11Hz -0.0234144 -0.00697291
+ 2.704e+11Hz -0.0233993 -0.00696139
+ 2.705e+11Hz -0.0233844 -0.00695022
+ 2.706e+11Hz -0.0233697 -0.0069394
+ 2.707e+11Hz -0.0233552 -0.00692892
+ 2.708e+11Hz -0.0233408 -0.00691878
+ 2.709e+11Hz -0.0233266 -0.00690899
+ 2.71e+11Hz -0.0233127 -0.00689955
+ 2.711e+11Hz -0.0232989 -0.00689045
+ 2.712e+11Hz -0.0232854 -0.00688169
+ 2.713e+11Hz -0.0232722 -0.00687327
+ 2.714e+11Hz -0.0232592 -0.00686518
+ 2.715e+11Hz -0.0232466 -0.00685743
+ 2.716e+11Hz -0.0232342 -0.00685
+ 2.717e+11Hz -0.0232221 -0.00684291
+ 2.718e+11Hz -0.0232104 -0.00683613
+ 2.719e+11Hz -0.023199 -0.00682966
+ 2.72e+11Hz -0.023188 -0.0068235
+ 2.721e+11Hz -0.0231773 -0.00681764
+ 2.722e+11Hz -0.023167 -0.00681208
+ 2.723e+11Hz -0.0231572 -0.0068068
+ 2.724e+11Hz -0.0231477 -0.00680181
+ 2.725e+11Hz -0.0231387 -0.00679708
+ 2.726e+11Hz -0.0231301 -0.00679261
+ 2.727e+11Hz -0.0231219 -0.00678839
+ 2.728e+11Hz -0.0231142 -0.00678441
+ 2.729e+11Hz -0.023107 -0.00678067
+ 2.73e+11Hz -0.0231003 -0.00677714
+ 2.731e+11Hz -0.0230941 -0.00677382
+ 2.732e+11Hz -0.0230885 -0.00677069
+ 2.733e+11Hz -0.0230833 -0.00676774
+ 2.734e+11Hz -0.0230787 -0.00676496
+ 2.735e+11Hz -0.0230746 -0.00676234
+ 2.736e+11Hz -0.0230711 -0.00675986
+ 2.737e+11Hz -0.0230682 -0.0067575
+ 2.738e+11Hz -0.0230659 -0.00675526
+ 2.739e+11Hz -0.0230642 -0.00675311
+ 2.74e+11Hz -0.023063 -0.00675104
+ 2.741e+11Hz -0.0230625 -0.00674903
+ 2.742e+11Hz -0.0230626 -0.00674707
+ 2.743e+11Hz -0.0230633 -0.00674514
+ 2.744e+11Hz -0.0230647 -0.00674322
+ 2.745e+11Hz -0.0230667 -0.0067413
+ 2.746e+11Hz -0.0230693 -0.00673936
+ 2.747e+11Hz -0.0230727 -0.00673737
+ 2.748e+11Hz -0.0230766 -0.00673532
+ 2.749e+11Hz -0.0230813 -0.00673319
+ 2.75e+11Hz -0.0230866 -0.00673096
+ 2.751e+11Hz -0.0230926 -0.00672862
+ 2.752e+11Hz -0.0230993 -0.00672613
+ 2.753e+11Hz -0.0231067 -0.00672349
+ 2.754e+11Hz -0.0231148 -0.00672067
+ 2.755e+11Hz -0.0231235 -0.00671764
+ 2.756e+11Hz -0.023133 -0.0067144
+ 2.757e+11Hz -0.0231431 -0.00671092
+ 2.758e+11Hz -0.0231539 -0.00670717
+ 2.759e+11Hz -0.0231655 -0.00670314
+ 2.76e+11Hz -0.0231777 -0.0066988
+ 2.761e+11Hz -0.0231906 -0.00669414
+ 2.762e+11Hz -0.0232042 -0.00668913
+ 2.763e+11Hz -0.0232185 -0.00668375
+ 2.764e+11Hz -0.0232335 -0.00667798
+ 2.765e+11Hz -0.0232492 -0.00667179
+ 2.766e+11Hz -0.0232655 -0.00666517
+ 2.767e+11Hz -0.0232825 -0.00665809
+ 2.768e+11Hz -0.0233002 -0.00665053
+ 2.769e+11Hz -0.0233185 -0.00664247
+ 2.77e+11Hz -0.0233375 -0.00663389
+ 2.771e+11Hz -0.0233572 -0.00662477
+ 2.772e+11Hz -0.0233774 -0.00661508
+ 2.773e+11Hz -0.0233983 -0.0066048
+ 2.774e+11Hz -0.0234199 -0.00659392
+ 2.775e+11Hz -0.023442 -0.0065824
+ 2.776e+11Hz -0.0234647 -0.00657024
+ 2.777e+11Hz -0.0234881 -0.0065574
+ 2.778e+11Hz -0.023512 -0.00654387
+ 2.779e+11Hz -0.0235364 -0.00652963
+ 2.78e+11Hz -0.0235615 -0.00651466
+ 2.781e+11Hz -0.023587 -0.00649893
+ 2.782e+11Hz -0.0236131 -0.00648243
+ 2.783e+11Hz -0.0236397 -0.00646513
+ 2.784e+11Hz -0.0236668 -0.00644703
+ 2.785e+11Hz -0.0236943 -0.00642809
+ 2.786e+11Hz -0.0237224 -0.0064083
+ 2.787e+11Hz -0.0237509 -0.00638765
+ 2.788e+11Hz -0.0237798 -0.00636611
+ 2.789e+11Hz -0.0238091 -0.00634367
+ 2.79e+11Hz -0.0238388 -0.00632031
+ 2.791e+11Hz -0.0238689 -0.00629601
+ 2.792e+11Hz -0.0238993 -0.00627075
+ 2.793e+11Hz -0.0239301 -0.00624453
+ 2.794e+11Hz -0.0239612 -0.00621732
+ 2.795e+11Hz -0.0239925 -0.00618911
+ 2.796e+11Hz -0.0240242 -0.00615989
+ 2.797e+11Hz -0.0240561 -0.00612964
+ 2.798e+11Hz -0.0240882 -0.00609834
+ 2.799e+11Hz -0.0241205 -0.00606599
+ 2.8e+11Hz -0.024153 -0.00603257
+ 2.801e+11Hz -0.0241857 -0.00599807
+ 2.802e+11Hz -0.0242185 -0.00596247
+ 2.803e+11Hz -0.0242514 -0.00592577
+ 2.804e+11Hz -0.0242844 -0.00588796
+ 2.805e+11Hz -0.0243175 -0.00584902
+ 2.806e+11Hz -0.0243506 -0.00580895
+ 2.807e+11Hz -0.0243837 -0.00576773
+ 2.808e+11Hz -0.0244168 -0.00572537
+ 2.809e+11Hz -0.0244498 -0.00568184
+ 2.81e+11Hz -0.0244828 -0.00563715
+ 2.811e+11Hz -0.0245157 -0.00559129
+ 2.812e+11Hz -0.0245485 -0.00554424
+ 2.813e+11Hz -0.0245811 -0.00549602
+ 2.814e+11Hz -0.0246135 -0.0054466
+ 2.815e+11Hz -0.0246457 -0.005396
+ 2.816e+11Hz -0.0246777 -0.0053442
+ 2.817e+11Hz -0.0247095 -0.00529119
+ 2.818e+11Hz -0.0247409 -0.00523699
+ 2.819e+11Hz -0.0247721 -0.00518159
+ 2.82e+11Hz -0.0248029 -0.00512498
+ 2.821e+11Hz -0.0248333 -0.00506718
+ 2.822e+11Hz -0.0248633 -0.00500816
+ 2.823e+11Hz -0.0248929 -0.00494795
+ 2.824e+11Hz -0.024922 -0.00488654
+ 2.825e+11Hz -0.0249507 -0.00482393
+ 2.826e+11Hz -0.0249788 -0.00476013
+ 2.827e+11Hz -0.0250064 -0.00469514
+ 2.828e+11Hz -0.0250334 -0.00462896
+ 2.829e+11Hz -0.0250598 -0.0045616
+ 2.83e+11Hz -0.0250856 -0.00449307
+ 2.831e+11Hz -0.0251107 -0.00442337
+ 2.832e+11Hz -0.0251351 -0.00435251
+ 2.833e+11Hz -0.0251588 -0.0042805
+ 2.834e+11Hz -0.0251818 -0.00420734
+ 2.835e+11Hz -0.025204 -0.00413305
+ 2.836e+11Hz -0.0252254 -0.00405764
+ 2.837e+11Hz -0.025246 -0.00398111
+ 2.838e+11Hz -0.0252657 -0.00390347
+ 2.839e+11Hz -0.0252845 -0.00382475
+ 2.84e+11Hz -0.0253024 -0.00374494
+ 2.841e+11Hz -0.0253194 -0.00366407
+ 2.842e+11Hz -0.0253355 -0.00358215
+ 2.843e+11Hz -0.0253505 -0.00349918
+ 2.844e+11Hz -0.0253645 -0.0034152
+ 2.845e+11Hz -0.0253775 -0.00333021
+ 2.846e+11Hz -0.0253894 -0.00324422
+ 2.847e+11Hz -0.0254002 -0.00315726
+ 2.848e+11Hz -0.0254099 -0.00306935
+ 2.849e+11Hz -0.0254184 -0.00298049
+ 2.85e+11Hz -0.0254258 -0.00289072
+ 2.851e+11Hz -0.0254319 -0.00280004
+ 2.852e+11Hz -0.0254369 -0.00270848
+ 2.853e+11Hz -0.0254406 -0.00261606
+ 2.854e+11Hz -0.0254431 -0.0025228
+ 2.855e+11Hz -0.0254442 -0.00242872
+ 2.856e+11Hz -0.0254441 -0.00233384
+ 2.857e+11Hz -0.0254426 -0.00223819
+ 2.858e+11Hz -0.0254398 -0.00214178
+ 2.859e+11Hz -0.0254356 -0.00204465
+ 2.86e+11Hz -0.02543 -0.00194681
+ 2.861e+11Hz -0.025423 -0.00184829
+ 2.862e+11Hz -0.0254146 -0.00174912
+ 2.863e+11Hz -0.0254047 -0.00164931
+ 2.864e+11Hz -0.0253933 -0.0015489
+ 2.865e+11Hz -0.0253805 -0.00144792
+ 2.866e+11Hz -0.0253662 -0.00134638
+ 2.867e+11Hz -0.0253503 -0.00124432
+ 2.868e+11Hz -0.0253329 -0.00114176
+ 2.869e+11Hz -0.0253139 -0.00103873
+ 2.87e+11Hz -0.0252934 -0.000935263
+ 2.871e+11Hz -0.0252713 -0.000831383
+ 2.872e+11Hz -0.0252476 -0.00072712
+ 2.873e+11Hz -0.0252222 -0.000622504
+ 2.874e+11Hz -0.0251953 -0.000517563
+ 2.875e+11Hz -0.0251667 -0.00041233
+ 2.876e+11Hz -0.0251365 -0.000306832
+ 2.877e+11Hz -0.0251046 -0.000201102
+ 2.878e+11Hz -0.025071 -9.51702e-05
+ 2.879e+11Hz -0.0250358 1.09327e-05
+ 2.88e+11Hz -0.0249988 0.000117175
+ 2.881e+11Hz -0.0249602 0.000223525
+ 2.882e+11Hz -0.0249199 0.000329951
+ 2.883e+11Hz -0.0248779 0.000436421
+ 2.884e+11Hz -0.0248341 0.000542902
+ 2.885e+11Hz -0.0247886 0.000649363
+ 2.886e+11Hz -0.0247414 0.00075577
+ 2.887e+11Hz -0.0246925 0.00086209
+ 2.888e+11Hz -0.0246418 0.000968292
+ 2.889e+11Hz -0.0245894 0.00107434
+ 2.89e+11Hz -0.0245352 0.00118021
+ 2.891e+11Hz -0.0244793 0.00128585
+ 2.892e+11Hz -0.0244216 0.00139124
+ 2.893e+11Hz -0.0243622 0.00149635
+ 2.894e+11Hz -0.0243011 0.00160114
+ 2.895e+11Hz -0.0242382 0.00170558
+ 2.896e+11Hz -0.0241736 0.00180963
+ 2.897e+11Hz -0.0241072 0.00191326
+ 2.898e+11Hz -0.0240391 0.00201644
+ 2.899e+11Hz -0.0239692 0.00211914
+ 2.9e+11Hz -0.0238977 0.00222131
+ 2.901e+11Hz -0.0238244 0.00232293
+ 2.902e+11Hz -0.0237493 0.00242397
+ 2.903e+11Hz -0.0236726 0.00252439
+ 2.904e+11Hz -0.0235942 0.00262415
+ 2.905e+11Hz -0.023514 0.00272323
+ 2.906e+11Hz -0.0234322 0.00282159
+ 2.907e+11Hz -0.0233487 0.0029192
+ 2.908e+11Hz -0.0232636 0.00301602
+ 2.909e+11Hz -0.0231767 0.00311203
+ 2.91e+11Hz -0.0230883 0.00320719
+ 2.911e+11Hz -0.0229982 0.00330147
+ 2.912e+11Hz -0.0229064 0.00339484
+ 2.913e+11Hz -0.0228131 0.00348727
+ 2.914e+11Hz -0.0227182 0.00357872
+ 2.915e+11Hz -0.0226217 0.00366916
+ 2.916e+11Hz -0.0225236 0.00375857
+ 2.917e+11Hz -0.022424 0.00384691
+ 2.918e+11Hz -0.0223228 0.00393415
+ 2.919e+11Hz -0.0222201 0.00402026
+ 2.92e+11Hz -0.022116 0.00410522
+ 2.921e+11Hz -0.0220103 0.00418899
+ 2.922e+11Hz -0.0219032 0.00427155
+ 2.923e+11Hz -0.0217947 0.00435286
+ 2.924e+11Hz -0.0216847 0.0044329
+ 2.925e+11Hz -0.0215733 0.00451164
+ 2.926e+11Hz -0.0214606 0.00458905
+ 2.927e+11Hz -0.0213465 0.00466511
+ 2.928e+11Hz -0.021231 0.00473979
+ 2.929e+11Hz -0.0211143 0.00481306
+ 2.93e+11Hz -0.0209962 0.0048849
+ 2.931e+11Hz -0.0208769 0.00495528
+ 2.932e+11Hz -0.0207564 0.00502418
+ 2.933e+11Hz -0.0206346 0.00509158
+ 2.934e+11Hz -0.0205117 0.00515744
+ 2.935e+11Hz -0.0203876 0.00522175
+ 2.936e+11Hz -0.0202624 0.00528448
+ 2.937e+11Hz -0.020136 0.00534562
+ 2.938e+11Hz -0.0200086 0.00540513
+ 2.939e+11Hz -0.0198801 0.00546301
+ 2.94e+11Hz -0.0197506 0.00551922
+ 2.941e+11Hz -0.0196201 0.00557375
+ 2.942e+11Hz -0.0194887 0.00562658
+ 2.943e+11Hz -0.0193563 0.00567769
+ 2.944e+11Hz -0.019223 0.00572706
+ 2.945e+11Hz -0.0190888 0.00577468
+ 2.946e+11Hz -0.0189538 0.00582053
+ 2.947e+11Hz -0.0188179 0.00586458
+ 2.948e+11Hz -0.0186813 0.00590683
+ 2.949e+11Hz -0.0185439 0.00594726
+ 2.95e+11Hz -0.0184059 0.00598586
+ 2.951e+11Hz -0.0182671 0.00602261
+ 2.952e+11Hz -0.0181277 0.00605749
+ 2.953e+11Hz -0.0179876 0.00609051
+ 2.954e+11Hz -0.017847 0.00612164
+ 2.955e+11Hz -0.0177058 0.00615087
+ 2.956e+11Hz -0.0175641 0.00617819
+ 2.957e+11Hz -0.0174219 0.0062036
+ 2.958e+11Hz -0.0172793 0.00622708
+ 2.959e+11Hz -0.0171363 0.00624862
+ 2.96e+11Hz -0.0169928 0.00626822
+ 2.961e+11Hz -0.016849 0.00628588
+ 2.962e+11Hz -0.016705 0.00630158
+ 2.963e+11Hz -0.0165606 0.00631531
+ 2.964e+11Hz -0.016416 0.00632708
+ 2.965e+11Hz -0.0162712 0.00633688
+ 2.966e+11Hz -0.0161262 0.00634471
+ 2.967e+11Hz -0.0159811 0.00635056
+ 2.968e+11Hz -0.0158359 0.00635443
+ 2.969e+11Hz -0.0156906 0.00635632
+ 2.97e+11Hz -0.0155453 0.00635623
+ 2.971e+11Hz -0.0154 0.00635416
+ 2.972e+11Hz -0.0152547 0.00635011
+ 2.973e+11Hz -0.0151095 0.00634408
+ 2.974e+11Hz -0.0149644 0.00633608
+ 2.975e+11Hz -0.0148195 0.0063261
+ 2.976e+11Hz -0.0146748 0.00631416
+ 2.977e+11Hz -0.0145302 0.00630025
+ 2.978e+11Hz -0.014386 0.00628438
+ 2.979e+11Hz -0.014242 0.00626656
+ 2.98e+11Hz -0.0140983 0.0062468
+ 2.981e+11Hz -0.013955 0.00622509
+ 2.982e+11Hz -0.0138121 0.00620146
+ 2.983e+11Hz -0.0136696 0.0061759
+ 2.984e+11Hz -0.0135276 0.00614843
+ 2.985e+11Hz -0.0133861 0.00611906
+ 2.986e+11Hz -0.0132451 0.0060878
+ 2.987e+11Hz -0.0131047 0.00605466
+ 2.988e+11Hz -0.0129648 0.00601965
+ 2.989e+11Hz -0.0128256 0.00598279
+ 2.99e+11Hz -0.0126871 0.00594408
+ 2.991e+11Hz -0.0125492 0.00590355
+ 2.992e+11Hz -0.0124121 0.00586121
+ 2.993e+11Hz -0.0122757 0.00581708
+ 2.994e+11Hz -0.0121401 0.00577116
+ 2.995e+11Hz -0.0120053 0.00572349
+ 2.996e+11Hz -0.0118714 0.00567407
+ 2.997e+11Hz -0.0117384 0.00562292
+ 2.998e+11Hz -0.0116062 0.00557007
+ 2.999e+11Hz -0.011475 0.00551552
+ 3e+11Hz -0.0113448 0.00545931
+ ]

A12 %vd(20 3) %vd(12, 3) xfer2
.model xfer2 xfer R_I=true table=[
+ 0Hz 0.990337 0
+ 1e+08Hz 0.990334 -0.0018782
+ 2e+08Hz 0.990325 -0.0037563
+ 3e+08Hz 0.99031 -0.00563423
+ 4e+08Hz 0.99029 -0.00751187
+ 5e+08Hz 0.990263 -0.00938915
+ 6e+08Hz 0.99023 -0.011266
+ 7e+08Hz 0.990191 -0.0131422
+ 8e+08Hz 0.990146 -0.0150179
+ 9e+08Hz 0.990095 -0.0168928
+ 1e+09Hz 0.990039 -0.0187669
+ 1.1e+09Hz 0.989977 -0.0206401
+ 1.2e+09Hz 0.989908 -0.0225123
+ 1.3e+09Hz 0.989834 -0.0243834
+ 1.4e+09Hz 0.989755 -0.0262534
+ 1.5e+09Hz 0.989669 -0.0281221
+ 1.6e+09Hz 0.989578 -0.0299895
+ 1.7e+09Hz 0.989482 -0.0318556
+ 1.8e+09Hz 0.989379 -0.0337201
+ 1.9e+09Hz 0.989272 -0.0355831
+ 2e+09Hz 0.989158 -0.0374445
+ 2.1e+09Hz 0.98904 -0.0393042
+ 2.2e+09Hz 0.988916 -0.0411622
+ 2.3e+09Hz 0.988787 -0.0430183
+ 2.4e+09Hz 0.988652 -0.0448725
+ 2.5e+09Hz 0.988512 -0.0467248
+ 2.6e+09Hz 0.988368 -0.0485751
+ 2.7e+09Hz 0.988218 -0.0504233
+ 2.8e+09Hz 0.988063 -0.0522694
+ 2.9e+09Hz 0.987903 -0.0541133
+ 3e+09Hz 0.987738 -0.055955
+ 3.1e+09Hz 0.987569 -0.0577944
+ 3.2e+09Hz 0.987395 -0.0596315
+ 3.3e+09Hz 0.987216 -0.0614663
+ 3.4e+09Hz 0.987033 -0.0632986
+ 3.5e+09Hz 0.986845 -0.0651285
+ 3.6e+09Hz 0.986653 -0.066956
+ 3.7e+09Hz 0.986457 -0.068781
+ 3.8e+09Hz 0.986256 -0.0706034
+ 3.9e+09Hz 0.986051 -0.0724233
+ 4e+09Hz 0.985842 -0.0742406
+ 4.1e+09Hz 0.985629 -0.0760554
+ 4.2e+09Hz 0.985413 -0.0778675
+ 4.3e+09Hz 0.985192 -0.0796771
+ 4.4e+09Hz 0.984967 -0.081484
+ 4.5e+09Hz 0.984739 -0.0832882
+ 4.6e+09Hz 0.984507 -0.0850898
+ 4.7e+09Hz 0.984272 -0.0868888
+ 4.8e+09Hz 0.984033 -0.0886851
+ 4.9e+09Hz 0.983791 -0.0904788
+ 5e+09Hz 0.983545 -0.0922699
+ 5.1e+09Hz 0.983296 -0.0940583
+ 5.2e+09Hz 0.983044 -0.0958441
+ 5.3e+09Hz 0.982789 -0.0976273
+ 5.4e+09Hz 0.982531 -0.0994079
+ 5.5e+09Hz 0.98227 -0.101186
+ 5.6e+09Hz 0.982006 -0.102961
+ 5.7e+09Hz 0.981739 -0.104734
+ 5.8e+09Hz 0.98147 -0.106505
+ 5.9e+09Hz 0.981197 -0.108273
+ 6e+09Hz 0.980922 -0.110038
+ 6.1e+09Hz 0.980645 -0.111801
+ 6.2e+09Hz 0.980365 -0.113562
+ 6.3e+09Hz 0.980082 -0.11532
+ 6.4e+09Hz 0.979798 -0.117076
+ 6.5e+09Hz 0.97951 -0.11883
+ 6.6e+09Hz 0.979221 -0.120581
+ 6.7e+09Hz 0.978929 -0.122331
+ 6.8e+09Hz 0.978635 -0.124078
+ 6.9e+09Hz 0.978339 -0.125823
+ 7e+09Hz 0.978041 -0.127566
+ 7.1e+09Hz 0.977741 -0.129307
+ 7.2e+09Hz 0.977439 -0.131045
+ 7.3e+09Hz 0.977134 -0.132782
+ 7.4e+09Hz 0.976828 -0.134517
+ 7.5e+09Hz 0.97652 -0.136251
+ 7.6e+09Hz 0.97621 -0.137982
+ 7.7e+09Hz 0.975898 -0.139712
+ 7.8e+09Hz 0.975585 -0.14144
+ 7.9e+09Hz 0.975269 -0.143166
+ 8e+09Hz 0.974952 -0.144891
+ 8.1e+09Hz 0.974633 -0.146614
+ 8.2e+09Hz 0.974312 -0.148336
+ 8.3e+09Hz 0.97399 -0.150056
+ 8.4e+09Hz 0.973666 -0.151775
+ 8.5e+09Hz 0.97334 -0.153493
+ 8.6e+09Hz 0.973012 -0.155209
+ 8.7e+09Hz 0.972683 -0.156924
+ 8.8e+09Hz 0.972352 -0.158638
+ 8.9e+09Hz 0.972019 -0.160351
+ 9e+09Hz 0.971685 -0.162063
+ 9.1e+09Hz 0.971349 -0.163774
+ 9.2e+09Hz 0.971012 -0.165484
+ 9.3e+09Hz 0.970672 -0.167193
+ 9.4e+09Hz 0.970331 -0.168901
+ 9.5e+09Hz 0.969989 -0.170608
+ 9.6e+09Hz 0.969644 -0.172315
+ 9.7e+09Hz 0.969298 -0.174021
+ 9.8e+09Hz 0.96895 -0.175726
+ 9.9e+09Hz 0.968601 -0.17743
+ 1e+10Hz 0.968249 -0.179134
+ 1.01e+10Hz 0.967896 -0.180838
+ 1.02e+10Hz 0.967541 -0.182541
+ 1.03e+10Hz 0.967184 -0.184243
+ 1.04e+10Hz 0.966825 -0.185945
+ 1.05e+10Hz 0.966464 -0.187647
+ 1.06e+10Hz 0.966102 -0.189348
+ 1.07e+10Hz 0.965737 -0.191049
+ 1.08e+10Hz 0.965371 -0.19275
+ 1.09e+10Hz 0.965002 -0.19445
+ 1.1e+10Hz 0.964632 -0.196151
+ 1.11e+10Hz 0.964259 -0.197851
+ 1.12e+10Hz 0.963884 -0.199551
+ 1.13e+10Hz 0.963507 -0.201251
+ 1.14e+10Hz 0.963128 -0.20295
+ 1.15e+10Hz 0.962747 -0.20465
+ 1.16e+10Hz 0.962363 -0.206349
+ 1.17e+10Hz 0.961977 -0.208049
+ 1.18e+10Hz 0.961589 -0.209748
+ 1.19e+10Hz 0.961198 -0.211447
+ 1.2e+10Hz 0.960805 -0.213147
+ 1.21e+10Hz 0.960409 -0.214846
+ 1.22e+10Hz 0.960011 -0.216545
+ 1.23e+10Hz 0.959611 -0.218245
+ 1.24e+10Hz 0.959207 -0.219944
+ 1.25e+10Hz 0.958802 -0.221643
+ 1.26e+10Hz 0.958393 -0.223343
+ 1.27e+10Hz 0.957982 -0.225042
+ 1.28e+10Hz 0.957568 -0.226742
+ 1.29e+10Hz 0.957151 -0.228441
+ 1.3e+10Hz 0.956732 -0.230141
+ 1.31e+10Hz 0.956309 -0.23184
+ 1.32e+10Hz 0.955884 -0.233539
+ 1.33e+10Hz 0.955455 -0.235239
+ 1.34e+10Hz 0.955024 -0.236938
+ 1.35e+10Hz 0.95459 -0.238638
+ 1.36e+10Hz 0.954152 -0.240337
+ 1.37e+10Hz 0.953712 -0.242036
+ 1.38e+10Hz 0.953268 -0.243735
+ 1.39e+10Hz 0.952821 -0.245434
+ 1.4e+10Hz 0.952371 -0.247133
+ 1.41e+10Hz 0.951918 -0.248832
+ 1.42e+10Hz 0.951461 -0.25053
+ 1.43e+10Hz 0.951001 -0.252228
+ 1.44e+10Hz 0.950538 -0.253926
+ 1.45e+10Hz 0.950071 -0.255624
+ 1.46e+10Hz 0.949602 -0.257322
+ 1.47e+10Hz 0.949128 -0.259019
+ 1.48e+10Hz 0.948651 -0.260715
+ 1.49e+10Hz 0.948171 -0.262412
+ 1.5e+10Hz 0.947687 -0.264108
+ 1.51e+10Hz 0.9472 -0.265803
+ 1.52e+10Hz 0.946709 -0.267498
+ 1.53e+10Hz 0.946215 -0.269193
+ 1.54e+10Hz 0.945717 -0.270886
+ 1.55e+10Hz 0.945215 -0.27258
+ 1.56e+10Hz 0.94471 -0.274272
+ 1.57e+10Hz 0.944201 -0.275964
+ 1.58e+10Hz 0.943689 -0.277655
+ 1.59e+10Hz 0.943173 -0.279346
+ 1.6e+10Hz 0.942653 -0.281035
+ 1.61e+10Hz 0.94213 -0.282724
+ 1.62e+10Hz 0.941603 -0.284412
+ 1.63e+10Hz 0.941073 -0.286099
+ 1.64e+10Hz 0.940539 -0.287785
+ 1.65e+10Hz 0.940001 -0.28947
+ 1.66e+10Hz 0.93946 -0.291154
+ 1.67e+10Hz 0.938915 -0.292837
+ 1.68e+10Hz 0.938366 -0.294519
+ 1.69e+10Hz 0.937814 -0.296199
+ 1.7e+10Hz 0.937258 -0.297878
+ 1.71e+10Hz 0.936698 -0.299557
+ 1.72e+10Hz 0.936135 -0.301234
+ 1.73e+10Hz 0.935568 -0.302909
+ 1.74e+10Hz 0.934998 -0.304583
+ 1.75e+10Hz 0.934424 -0.306256
+ 1.76e+10Hz 0.933847 -0.307927
+ 1.77e+10Hz 0.933266 -0.309597
+ 1.78e+10Hz 0.932682 -0.311266
+ 1.79e+10Hz 0.932094 -0.312933
+ 1.8e+10Hz 0.931503 -0.314598
+ 1.81e+10Hz 0.930908 -0.316262
+ 1.82e+10Hz 0.93031 -0.317924
+ 1.83e+10Hz 0.929708 -0.319585
+ 1.84e+10Hz 0.929104 -0.321244
+ 1.85e+10Hz 0.928495 -0.322901
+ 1.86e+10Hz 0.927884 -0.324556
+ 1.87e+10Hz 0.927269 -0.32621
+ 1.88e+10Hz 0.926651 -0.327862
+ 1.89e+10Hz 0.92603 -0.329512
+ 1.9e+10Hz 0.925406 -0.331161
+ 1.91e+10Hz 0.924778 -0.332807
+ 1.92e+10Hz 0.924148 -0.334452
+ 1.93e+10Hz 0.923514 -0.336095
+ 1.94e+10Hz 0.922877 -0.337736
+ 1.95e+10Hz 0.922238 -0.339375
+ 1.96e+10Hz 0.921595 -0.341012
+ 1.97e+10Hz 0.920949 -0.342647
+ 1.98e+10Hz 0.920301 -0.344281
+ 1.99e+10Hz 0.919649 -0.345912
+ 2e+10Hz 0.918995 -0.347542
+ 2.01e+10Hz 0.918338 -0.349169
+ 2.02e+10Hz 0.917678 -0.350795
+ 2.03e+10Hz 0.917015 -0.352419
+ 2.04e+10Hz 0.91635 -0.354041
+ 2.05e+10Hz 0.915682 -0.35566
+ 2.06e+10Hz 0.915011 -0.357278
+ 2.07e+10Hz 0.914338 -0.358894
+ 2.08e+10Hz 0.913662 -0.360508
+ 2.09e+10Hz 0.912984 -0.36212
+ 2.1e+10Hz 0.912303 -0.363731
+ 2.11e+10Hz 0.911619 -0.365339
+ 2.12e+10Hz 0.910933 -0.366945
+ 2.13e+10Hz 0.910245 -0.36855
+ 2.14e+10Hz 0.909554 -0.370153
+ 2.15e+10Hz 0.908861 -0.371753
+ 2.16e+10Hz 0.908166 -0.373352
+ 2.17e+10Hz 0.907468 -0.374949
+ 2.18e+10Hz 0.906768 -0.376545
+ 2.19e+10Hz 0.906066 -0.378138
+ 2.2e+10Hz 0.905361 -0.37973
+ 2.21e+10Hz 0.904655 -0.38132
+ 2.22e+10Hz 0.903946 -0.382908
+ 2.23e+10Hz 0.903235 -0.384495
+ 2.24e+10Hz 0.902522 -0.386079
+ 2.25e+10Hz 0.901806 -0.387663
+ 2.26e+10Hz 0.901089 -0.389244
+ 2.27e+10Hz 0.900369 -0.390824
+ 2.28e+10Hz 0.899647 -0.392402
+ 2.29e+10Hz 0.898923 -0.393979
+ 2.3e+10Hz 0.898198 -0.395554
+ 2.31e+10Hz 0.89747 -0.397128
+ 2.32e+10Hz 0.89674 -0.3987
+ 2.33e+10Hz 0.896008 -0.40027
+ 2.34e+10Hz 0.895274 -0.401839
+ 2.35e+10Hz 0.894538 -0.403407
+ 2.36e+10Hz 0.8938 -0.404973
+ 2.37e+10Hz 0.89306 -0.406538
+ 2.38e+10Hz 0.892317 -0.408102
+ 2.39e+10Hz 0.891573 -0.409664
+ 2.4e+10Hz 0.890827 -0.411225
+ 2.41e+10Hz 0.890079 -0.412785
+ 2.42e+10Hz 0.889329 -0.414343
+ 2.43e+10Hz 0.888577 -0.4159
+ 2.44e+10Hz 0.887822 -0.417456
+ 2.45e+10Hz 0.887066 -0.419011
+ 2.46e+10Hz 0.886308 -0.420565
+ 2.47e+10Hz 0.885548 -0.422117
+ 2.48e+10Hz 0.884785 -0.423669
+ 2.49e+10Hz 0.884021 -0.425219
+ 2.5e+10Hz 0.883254 -0.426768
+ 2.51e+10Hz 0.882486 -0.428316
+ 2.52e+10Hz 0.881715 -0.429864
+ 2.53e+10Hz 0.880942 -0.43141
+ 2.54e+10Hz 0.880167 -0.432955
+ 2.55e+10Hz 0.87939 -0.434499
+ 2.56e+10Hz 0.87861 -0.436043
+ 2.57e+10Hz 0.877829 -0.437585
+ 2.58e+10Hz 0.877045 -0.439126
+ 2.59e+10Hz 0.876259 -0.440667
+ 2.6e+10Hz 0.875471 -0.442207
+ 2.61e+10Hz 0.87468 -0.443745
+ 2.62e+10Hz 0.873887 -0.445283
+ 2.63e+10Hz 0.873092 -0.44682
+ 2.64e+10Hz 0.872295 -0.448357
+ 2.65e+10Hz 0.871495 -0.449892
+ 2.66e+10Hz 0.870693 -0.451427
+ 2.67e+10Hz 0.869888 -0.45296
+ 2.68e+10Hz 0.869081 -0.454493
+ 2.69e+10Hz 0.868271 -0.456025
+ 2.7e+10Hz 0.867459 -0.457557
+ 2.71e+10Hz 0.866644 -0.459087
+ 2.72e+10Hz 0.865827 -0.460617
+ 2.73e+10Hz 0.865008 -0.462146
+ 2.74e+10Hz 0.864185 -0.463674
+ 2.75e+10Hz 0.86336 -0.465201
+ 2.76e+10Hz 0.862533 -0.466727
+ 2.77e+10Hz 0.861703 -0.468253
+ 2.78e+10Hz 0.86087 -0.469778
+ 2.79e+10Hz 0.860034 -0.471301
+ 2.8e+10Hz 0.859195 -0.472825
+ 2.81e+10Hz 0.858354 -0.474347
+ 2.82e+10Hz 0.85751 -0.475868
+ 2.83e+10Hz 0.856663 -0.477388
+ 2.84e+10Hz 0.855814 -0.478908
+ 2.85e+10Hz 0.854961 -0.480427
+ 2.86e+10Hz 0.854106 -0.481944
+ 2.87e+10Hz 0.853247 -0.483461
+ 2.88e+10Hz 0.852386 -0.484977
+ 2.89e+10Hz 0.851522 -0.486492
+ 2.9e+10Hz 0.850654 -0.488006
+ 2.91e+10Hz 0.849784 -0.489519
+ 2.92e+10Hz 0.848911 -0.49103
+ 2.93e+10Hz 0.848034 -0.492541
+ 2.94e+10Hz 0.847155 -0.494051
+ 2.95e+10Hz 0.846273 -0.495559
+ 2.96e+10Hz 0.845387 -0.497067
+ 2.97e+10Hz 0.844498 -0.498573
+ 2.98e+10Hz 0.843606 -0.500078
+ 2.99e+10Hz 0.842711 -0.501582
+ 3e+10Hz 0.841813 -0.503084
+ 3.01e+10Hz 0.840912 -0.504586
+ 3.02e+10Hz 0.840008 -0.506086
+ 3.03e+10Hz 0.8391 -0.507585
+ 3.04e+10Hz 0.838189 -0.509082
+ 3.05e+10Hz 0.837275 -0.510578
+ 3.06e+10Hz 0.836358 -0.512073
+ 3.07e+10Hz 0.835437 -0.513566
+ 3.08e+10Hz 0.834513 -0.515058
+ 3.09e+10Hz 0.833587 -0.516548
+ 3.1e+10Hz 0.832656 -0.518037
+ 3.11e+10Hz 0.831723 -0.519524
+ 3.12e+10Hz 0.830786 -0.521009
+ 3.13e+10Hz 0.829846 -0.522493
+ 3.14e+10Hz 0.828903 -0.523975
+ 3.15e+10Hz 0.827957 -0.525456
+ 3.16e+10Hz 0.827008 -0.526935
+ 3.17e+10Hz 0.826055 -0.528412
+ 3.18e+10Hz 0.825099 -0.529887
+ 3.19e+10Hz 0.82414 -0.531361
+ 3.2e+10Hz 0.823177 -0.532833
+ 3.21e+10Hz 0.822212 -0.534302
+ 3.22e+10Hz 0.821243 -0.53577
+ 3.23e+10Hz 0.820271 -0.537236
+ 3.24e+10Hz 0.819296 -0.5387
+ 3.25e+10Hz 0.818318 -0.540162
+ 3.26e+10Hz 0.817337 -0.541622
+ 3.27e+10Hz 0.816353 -0.54308
+ 3.28e+10Hz 0.815365 -0.544536
+ 3.29e+10Hz 0.814375 -0.54599
+ 3.3e+10Hz 0.813381 -0.547442
+ 3.31e+10Hz 0.812385 -0.548892
+ 3.32e+10Hz 0.811385 -0.550339
+ 3.33e+10Hz 0.810382 -0.551784
+ 3.34e+10Hz 0.809377 -0.553227
+ 3.35e+10Hz 0.808368 -0.554668
+ 3.36e+10Hz 0.807357 -0.556107
+ 3.37e+10Hz 0.806342 -0.557543
+ 3.38e+10Hz 0.805325 -0.558977
+ 3.39e+10Hz 0.804305 -0.560408
+ 3.4e+10Hz 0.803282 -0.561838
+ 3.41e+10Hz 0.802256 -0.563265
+ 3.42e+10Hz 0.801228 -0.564689
+ 3.43e+10Hz 0.800197 -0.566112
+ 3.44e+10Hz 0.799163 -0.567531
+ 3.45e+10Hz 0.798126 -0.568949
+ 3.46e+10Hz 0.797087 -0.570364
+ 3.47e+10Hz 0.796045 -0.571777
+ 3.48e+10Hz 0.795 -0.573187
+ 3.49e+10Hz 0.793953 -0.574594
+ 3.5e+10Hz 0.792903 -0.576
+ 3.51e+10Hz 0.791851 -0.577403
+ 3.52e+10Hz 0.790796 -0.578803
+ 3.53e+10Hz 0.789738 -0.580201
+ 3.54e+10Hz 0.788679 -0.581596
+ 3.55e+10Hz 0.787616 -0.582989
+ 3.56e+10Hz 0.786552 -0.58438
+ 3.57e+10Hz 0.785485 -0.585768
+ 3.58e+10Hz 0.784415 -0.587153
+ 3.59e+10Hz 0.783344 -0.588536
+ 3.6e+10Hz 0.78227 -0.589917
+ 3.61e+10Hz 0.781194 -0.591295
+ 3.62e+10Hz 0.780115 -0.592671
+ 3.63e+10Hz 0.779035 -0.594044
+ 3.64e+10Hz 0.777952 -0.595415
+ 3.65e+10Hz 0.776867 -0.596783
+ 3.66e+10Hz 0.77578 -0.598149
+ 3.67e+10Hz 0.77469 -0.599512
+ 3.68e+10Hz 0.773599 -0.600873
+ 3.69e+10Hz 0.772506 -0.602232
+ 3.7e+10Hz 0.77141 -0.603588
+ 3.71e+10Hz 0.770313 -0.604942
+ 3.72e+10Hz 0.769213 -0.606294
+ 3.73e+10Hz 0.768112 -0.607643
+ 3.74e+10Hz 0.767008 -0.60899
+ 3.75e+10Hz 0.765903 -0.610334
+ 3.76e+10Hz 0.764795 -0.611676
+ 3.77e+10Hz 0.763686 -0.613016
+ 3.78e+10Hz 0.762575 -0.614354
+ 3.79e+10Hz 0.761462 -0.615689
+ 3.8e+10Hz 0.760347 -0.617022
+ 3.81e+10Hz 0.75923 -0.618353
+ 3.82e+10Hz 0.758111 -0.619682
+ 3.83e+10Hz 0.756991 -0.621008
+ 3.84e+10Hz 0.755868 -0.622332
+ 3.85e+10Hz 0.754744 -0.623654
+ 3.86e+10Hz 0.753618 -0.624974
+ 3.87e+10Hz 0.752491 -0.626292
+ 3.88e+10Hz 0.751361 -0.627608
+ 3.89e+10Hz 0.75023 -0.628921
+ 3.9e+10Hz 0.749097 -0.630233
+ 3.91e+10Hz 0.747962 -0.631542
+ 3.92e+10Hz 0.746825 -0.63285
+ 3.93e+10Hz 0.745686 -0.634155
+ 3.94e+10Hz 0.744546 -0.635458
+ 3.95e+10Hz 0.743404 -0.63676
+ 3.96e+10Hz 0.74226 -0.638059
+ 3.97e+10Hz 0.741115 -0.639357
+ 3.98e+10Hz 0.739967 -0.640652
+ 3.99e+10Hz 0.738818 -0.641946
+ 4e+10Hz 0.737667 -0.643238
+ 4.01e+10Hz 0.736515 -0.644528
+ 4.02e+10Hz 0.73536 -0.645816
+ 4.03e+10Hz 0.734204 -0.647102
+ 4.04e+10Hz 0.733045 -0.648387
+ 4.05e+10Hz 0.731885 -0.649669
+ 4.06e+10Hz 0.730724 -0.65095
+ 4.07e+10Hz 0.72956 -0.652229
+ 4.08e+10Hz 0.728395 -0.653506
+ 4.09e+10Hz 0.727227 -0.654782
+ 4.1e+10Hz 0.726058 -0.656055
+ 4.11e+10Hz 0.724887 -0.657327
+ 4.12e+10Hz 0.723714 -0.658597
+ 4.13e+10Hz 0.722539 -0.659866
+ 4.14e+10Hz 0.721362 -0.661133
+ 4.15e+10Hz 0.720183 -0.662398
+ 4.16e+10Hz 0.719003 -0.663661
+ 4.17e+10Hz 0.71782 -0.664923
+ 4.18e+10Hz 0.716635 -0.666183
+ 4.19e+10Hz 0.715448 -0.667441
+ 4.2e+10Hz 0.71426 -0.668698
+ 4.21e+10Hz 0.713069 -0.669953
+ 4.22e+10Hz 0.711876 -0.671207
+ 4.23e+10Hz 0.710681 -0.672458
+ 4.24e+10Hz 0.709485 -0.673708
+ 4.25e+10Hz 0.708286 -0.674957
+ 4.26e+10Hz 0.707084 -0.676203
+ 4.27e+10Hz 0.705881 -0.677448
+ 4.28e+10Hz 0.704676 -0.678692
+ 4.29e+10Hz 0.703468 -0.679934
+ 4.3e+10Hz 0.702259 -0.681174
+ 4.31e+10Hz 0.701047 -0.682412
+ 4.32e+10Hz 0.699832 -0.683649
+ 4.33e+10Hz 0.698616 -0.684884
+ 4.34e+10Hz 0.697397 -0.686117
+ 4.35e+10Hz 0.696177 -0.687349
+ 4.36e+10Hz 0.694953 -0.688579
+ 4.37e+10Hz 0.693728 -0.689807
+ 4.38e+10Hz 0.6925 -0.691033
+ 4.39e+10Hz 0.69127 -0.692258
+ 4.4e+10Hz 0.690038 -0.693481
+ 4.41e+10Hz 0.688803 -0.694702
+ 4.42e+10Hz 0.687566 -0.695922
+ 4.43e+10Hz 0.686326 -0.697139
+ 4.44e+10Hz 0.685084 -0.698355
+ 4.45e+10Hz 0.68384 -0.699569
+ 4.46e+10Hz 0.682593 -0.700781
+ 4.47e+10Hz 0.681344 -0.701991
+ 4.48e+10Hz 0.680092 -0.7032
+ 4.49e+10Hz 0.678838 -0.704406
+ 4.5e+10Hz 0.677581 -0.705611
+ 4.51e+10Hz 0.676322 -0.706814
+ 4.52e+10Hz 0.675061 -0.708014
+ 4.53e+10Hz 0.673797 -0.709213
+ 4.54e+10Hz 0.67253 -0.71041
+ 4.55e+10Hz 0.671261 -0.711605
+ 4.56e+10Hz 0.66999 -0.712797
+ 4.57e+10Hz 0.668716 -0.713988
+ 4.58e+10Hz 0.667439 -0.715177
+ 4.59e+10Hz 0.66616 -0.716363
+ 4.6e+10Hz 0.664878 -0.717548
+ 4.61e+10Hz 0.663594 -0.71873
+ 4.62e+10Hz 0.662307 -0.71991
+ 4.63e+10Hz 0.661018 -0.721088
+ 4.64e+10Hz 0.659726 -0.722264
+ 4.65e+10Hz 0.658432 -0.723437
+ 4.66e+10Hz 0.657135 -0.724609
+ 4.67e+10Hz 0.655836 -0.725778
+ 4.68e+10Hz 0.654534 -0.726944
+ 4.69e+10Hz 0.65323 -0.728109
+ 4.7e+10Hz 0.651923 -0.729271
+ 4.71e+10Hz 0.650613 -0.73043
+ 4.72e+10Hz 0.649302 -0.731588
+ 4.73e+10Hz 0.647987 -0.732743
+ 4.74e+10Hz 0.64667 -0.733895
+ 4.75e+10Hz 0.645351 -0.735045
+ 4.76e+10Hz 0.644029 -0.736193
+ 4.77e+10Hz 0.642705 -0.737338
+ 4.78e+10Hz 0.641378 -0.73848
+ 4.79e+10Hz 0.640049 -0.73962
+ 4.8e+10Hz 0.638717 -0.740758
+ 4.81e+10Hz 0.637383 -0.741893
+ 4.82e+10Hz 0.636047 -0.743025
+ 4.83e+10Hz 0.634708 -0.744154
+ 4.84e+10Hz 0.633367 -0.745282
+ 4.85e+10Hz 0.632023 -0.746406
+ 4.86e+10Hz 0.630678 -0.747528
+ 4.87e+10Hz 0.629329 -0.748647
+ 4.88e+10Hz 0.627979 -0.749763
+ 4.89e+10Hz 0.626626 -0.750877
+ 4.9e+10Hz 0.625271 -0.751987
+ 4.91e+10Hz 0.623914 -0.753096
+ 4.92e+10Hz 0.622554 -0.754201
+ 4.93e+10Hz 0.621193 -0.755304
+ 4.94e+10Hz 0.619829 -0.756403
+ 4.95e+10Hz 0.618463 -0.7575
+ 4.96e+10Hz 0.617095 -0.758595
+ 4.97e+10Hz 0.615724 -0.759686
+ 4.98e+10Hz 0.614352 -0.760774
+ 4.99e+10Hz 0.612977 -0.76186
+ 5e+10Hz 0.6116 -0.762943
+ 5.01e+10Hz 0.610222 -0.764023
+ 5.02e+10Hz 0.608841 -0.7651
+ 5.03e+10Hz 0.607458 -0.766174
+ 5.04e+10Hz 0.606074 -0.767246
+ 5.05e+10Hz 0.604687 -0.768314
+ 5.06e+10Hz 0.603298 -0.76938
+ 5.07e+10Hz 0.601908 -0.770443
+ 5.08e+10Hz 0.600515 -0.771502
+ 5.09e+10Hz 0.599121 -0.772559
+ 5.1e+10Hz 0.597725 -0.773613
+ 5.11e+10Hz 0.596327 -0.774665
+ 5.12e+10Hz 0.594927 -0.775713
+ 5.13e+10Hz 0.593526 -0.776758
+ 5.14e+10Hz 0.592122 -0.777801
+ 5.15e+10Hz 0.590717 -0.77884
+ 5.16e+10Hz 0.58931 -0.779877
+ 5.17e+10Hz 0.587902 -0.780911
+ 5.18e+10Hz 0.586492 -0.781941
+ 5.19e+10Hz 0.58508 -0.782969
+ 5.2e+10Hz 0.583666 -0.783995
+ 5.21e+10Hz 0.582251 -0.785017
+ 5.22e+10Hz 0.580834 -0.786036
+ 5.23e+10Hz 0.579416 -0.787053
+ 5.24e+10Hz 0.577996 -0.788067
+ 5.25e+10Hz 0.576574 -0.789077
+ 5.26e+10Hz 0.575151 -0.790085
+ 5.27e+10Hz 0.573726 -0.791091
+ 5.28e+10Hz 0.5723 -0.792093
+ 5.29e+10Hz 0.570873 -0.793093
+ 5.3e+10Hz 0.569443 -0.794089
+ 5.31e+10Hz 0.568013 -0.795083
+ 5.32e+10Hz 0.566581 -0.796075
+ 5.33e+10Hz 0.565147 -0.797063
+ 5.34e+10Hz 0.563712 -0.798049
+ 5.35e+10Hz 0.562276 -0.799032
+ 5.36e+10Hz 0.560838 -0.800012
+ 5.37e+10Hz 0.559399 -0.80099
+ 5.38e+10Hz 0.557958 -0.801965
+ 5.39e+10Hz 0.556516 -0.802937
+ 5.4e+10Hz 0.555072 -0.803906
+ 5.41e+10Hz 0.553628 -0.804873
+ 5.42e+10Hz 0.552182 -0.805837
+ 5.43e+10Hz 0.550734 -0.806799
+ 5.44e+10Hz 0.549285 -0.807758
+ 5.45e+10Hz 0.547835 -0.808714
+ 5.46e+10Hz 0.546383 -0.809668
+ 5.47e+10Hz 0.54493 -0.810619
+ 5.48e+10Hz 0.543476 -0.811567
+ 5.49e+10Hz 0.54202 -0.812513
+ 5.5e+10Hz 0.540563 -0.813456
+ 5.51e+10Hz 0.539105 -0.814397
+ 5.52e+10Hz 0.537645 -0.815336
+ 5.53e+10Hz 0.536184 -0.816271
+ 5.54e+10Hz 0.534722 -0.817205
+ 5.55e+10Hz 0.533258 -0.818136
+ 5.56e+10Hz 0.531793 -0.819064
+ 5.57e+10Hz 0.530327 -0.81999
+ 5.58e+10Hz 0.528859 -0.820913
+ 5.59e+10Hz 0.52739 -0.821834
+ 5.6e+10Hz 0.52592 -0.822753
+ 5.61e+10Hz 0.524448 -0.823669
+ 5.62e+10Hz 0.522975 -0.824582
+ 5.63e+10Hz 0.5215 -0.825494
+ 5.64e+10Hz 0.520024 -0.826402
+ 5.65e+10Hz 0.518547 -0.827309
+ 5.66e+10Hz 0.517068 -0.828213
+ 5.67e+10Hz 0.515588 -0.829115
+ 5.68e+10Hz 0.514106 -0.830014
+ 5.69e+10Hz 0.512623 -0.830911
+ 5.7e+10Hz 0.511139 -0.831805
+ 5.71e+10Hz 0.509653 -0.832697
+ 5.72e+10Hz 0.508166 -0.833587
+ 5.73e+10Hz 0.506677 -0.834475
+ 5.74e+10Hz 0.505187 -0.83536
+ 5.75e+10Hz 0.503695 -0.836242
+ 5.76e+10Hz 0.502202 -0.837123
+ 5.77e+10Hz 0.500707 -0.838001
+ 5.78e+10Hz 0.499211 -0.838876
+ 5.79e+10Hz 0.497713 -0.83975
+ 5.8e+10Hz 0.496214 -0.840621
+ 5.81e+10Hz 0.494713 -0.841489
+ 5.82e+10Hz 0.493211 -0.842355
+ 5.83e+10Hz 0.491707 -0.843219
+ 5.84e+10Hz 0.490201 -0.844081
+ 5.85e+10Hz 0.488694 -0.84494
+ 5.86e+10Hz 0.487186 -0.845797
+ 5.87e+10Hz 0.485675 -0.846651
+ 5.88e+10Hz 0.484163 -0.847503
+ 5.89e+10Hz 0.48265 -0.848353
+ 5.9e+10Hz 0.481135 -0.8492
+ 5.91e+10Hz 0.479618 -0.850045
+ 5.92e+10Hz 0.478099 -0.850887
+ 5.93e+10Hz 0.476579 -0.851727
+ 5.94e+10Hz 0.475058 -0.852565
+ 5.95e+10Hz 0.473534 -0.8534
+ 5.96e+10Hz 0.472009 -0.854232
+ 5.97e+10Hz 0.470482 -0.855062
+ 5.98e+10Hz 0.468954 -0.85589
+ 5.99e+10Hz 0.467423 -0.856715
+ 6e+10Hz 0.465891 -0.857538
+ 6.01e+10Hz 0.464357 -0.858358
+ 6.02e+10Hz 0.462822 -0.859176
+ 6.03e+10Hz 0.461285 -0.859991
+ 6.04e+10Hz 0.459746 -0.860803
+ 6.05e+10Hz 0.458205 -0.861613
+ 6.06e+10Hz 0.456663 -0.862421
+ 6.07e+10Hz 0.455119 -0.863225
+ 6.08e+10Hz 0.453573 -0.864028
+ 6.09e+10Hz 0.452025 -0.864827
+ 6.1e+10Hz 0.450475 -0.865624
+ 6.11e+10Hz 0.448924 -0.866418
+ 6.12e+10Hz 0.447371 -0.86721
+ 6.13e+10Hz 0.445816 -0.867999
+ 6.14e+10Hz 0.44426 -0.868785
+ 6.15e+10Hz 0.442701 -0.869568
+ 6.16e+10Hz 0.441141 -0.870349
+ 6.17e+10Hz 0.43958 -0.871126
+ 6.18e+10Hz 0.438016 -0.871902
+ 6.19e+10Hz 0.436451 -0.872674
+ 6.2e+10Hz 0.434883 -0.873443
+ 6.21e+10Hz 0.433315 -0.87421
+ 6.22e+10Hz 0.431744 -0.874974
+ 6.23e+10Hz 0.430172 -0.875734
+ 6.24e+10Hz 0.428597 -0.876492
+ 6.25e+10Hz 0.427022 -0.877247
+ 6.26e+10Hz 0.425444 -0.877999
+ 6.27e+10Hz 0.423865 -0.878749
+ 6.28e+10Hz 0.422284 -0.879495
+ 6.29e+10Hz 0.420701 -0.880238
+ 6.3e+10Hz 0.419117 -0.880978
+ 6.31e+10Hz 0.417531 -0.881716
+ 6.32e+10Hz 0.415943 -0.88245
+ 6.33e+10Hz 0.414354 -0.883181
+ 6.34e+10Hz 0.412763 -0.883909
+ 6.35e+10Hz 0.41117 -0.884634
+ 6.36e+10Hz 0.409576 -0.885356
+ 6.37e+10Hz 0.40798 -0.886074
+ 6.38e+10Hz 0.406382 -0.88679
+ 6.39e+10Hz 0.404783 -0.887503
+ 6.4e+10Hz 0.403183 -0.888212
+ 6.41e+10Hz 0.401581 -0.888918
+ 6.42e+10Hz 0.399977 -0.889621
+ 6.43e+10Hz 0.398372 -0.890321
+ 6.44e+10Hz 0.396765 -0.891017
+ 6.45e+10Hz 0.395157 -0.891711
+ 6.46e+10Hz 0.393547 -0.892401
+ 6.47e+10Hz 0.391936 -0.893088
+ 6.48e+10Hz 0.390324 -0.893771
+ 6.49e+10Hz 0.38871 -0.894452
+ 6.5e+10Hz 0.387094 -0.895129
+ 6.51e+10Hz 0.385478 -0.895803
+ 6.52e+10Hz 0.383859 -0.896473
+ 6.53e+10Hz 0.38224 -0.89714
+ 6.54e+10Hz 0.380619 -0.897804
+ 6.55e+10Hz 0.378997 -0.898465
+ 6.56e+10Hz 0.377374 -0.899122
+ 6.57e+10Hz 0.375749 -0.899776
+ 6.58e+10Hz 0.374123 -0.900427
+ 6.59e+10Hz 0.372496 -0.901074
+ 6.6e+10Hz 0.370868 -0.901718
+ 6.61e+10Hz 0.369238 -0.902358
+ 6.62e+10Hz 0.367608 -0.902996
+ 6.63e+10Hz 0.365976 -0.903629
+ 6.64e+10Hz 0.364343 -0.90426
+ 6.65e+10Hz 0.362709 -0.904887
+ 6.66e+10Hz 0.361074 -0.905511
+ 6.67e+10Hz 0.359437 -0.906131
+ 6.68e+10Hz 0.3578 -0.906748
+ 6.69e+10Hz 0.356162 -0.907362
+ 6.7e+10Hz 0.354522 -0.907972
+ 6.71e+10Hz 0.352882 -0.908579
+ 6.72e+10Hz 0.351241 -0.909183
+ 6.73e+10Hz 0.349599 -0.909783
+ 6.74e+10Hz 0.347955 -0.91038
+ 6.75e+10Hz 0.346311 -0.910974
+ 6.76e+10Hz 0.344666 -0.911564
+ 6.77e+10Hz 0.34302 -0.912151
+ 6.78e+10Hz 0.341374 -0.912735
+ 6.79e+10Hz 0.339726 -0.913315
+ 6.8e+10Hz 0.338077 -0.913892
+ 6.81e+10Hz 0.336428 -0.914466
+ 6.82e+10Hz 0.334778 -0.915036
+ 6.83e+10Hz 0.333127 -0.915603
+ 6.84e+10Hz 0.331475 -0.916167
+ 6.85e+10Hz 0.329823 -0.916727
+ 6.86e+10Hz 0.32817 -0.917284
+ 6.87e+10Hz 0.326516 -0.917838
+ 6.88e+10Hz 0.324861 -0.918389
+ 6.89e+10Hz 0.323206 -0.918936
+ 6.9e+10Hz 0.32155 -0.91948
+ 6.91e+10Hz 0.319893 -0.920021
+ 6.92e+10Hz 0.318236 -0.920559
+ 6.93e+10Hz 0.316578 -0.921093
+ 6.94e+10Hz 0.314919 -0.921625
+ 6.95e+10Hz 0.31326 -0.922153
+ 6.96e+10Hz 0.3116 -0.922678
+ 6.97e+10Hz 0.309939 -0.923199
+ 6.98e+10Hz 0.308278 -0.923718
+ 6.99e+10Hz 0.306616 -0.924233
+ 7e+10Hz 0.304954 -0.924745
+ 7.01e+10Hz 0.303291 -0.925254
+ 7.02e+10Hz 0.301627 -0.92576
+ 7.03e+10Hz 0.299963 -0.926263
+ 7.04e+10Hz 0.298298 -0.926763
+ 7.05e+10Hz 0.296633 -0.92726
+ 7.06e+10Hz 0.294967 -0.927753
+ 7.07e+10Hz 0.293301 -0.928244
+ 7.08e+10Hz 0.291634 -0.928731
+ 7.09e+10Hz 0.289966 -0.929215
+ 7.1e+10Hz 0.288298 -0.929697
+ 7.11e+10Hz 0.286629 -0.930175
+ 7.12e+10Hz 0.28496 -0.93065
+ 7.13e+10Hz 0.28329 -0.931122
+ 7.14e+10Hz 0.28162 -0.931591
+ 7.15e+10Hz 0.279949 -0.932058
+ 7.16e+10Hz 0.278278 -0.932521
+ 7.17e+10Hz 0.276606 -0.932981
+ 7.18e+10Hz 0.274934 -0.933438
+ 7.19e+10Hz 0.273261 -0.933892
+ 7.2e+10Hz 0.271587 -0.934344
+ 7.21e+10Hz 0.269913 -0.934792
+ 7.22e+10Hz 0.268239 -0.935237
+ 7.23e+10Hz 0.266564 -0.93568
+ 7.24e+10Hz 0.264888 -0.936119
+ 7.25e+10Hz 0.263212 -0.936556
+ 7.26e+10Hz 0.261535 -0.936989
+ 7.27e+10Hz 0.259858 -0.93742
+ 7.28e+10Hz 0.25818 -0.937848
+ 7.29e+10Hz 0.256502 -0.938272
+ 7.3e+10Hz 0.254823 -0.938694
+ 7.31e+10Hz 0.253143 -0.939113
+ 7.32e+10Hz 0.251463 -0.939529
+ 7.33e+10Hz 0.249782 -0.939942
+ 7.34e+10Hz 0.248101 -0.940353
+ 7.35e+10Hz 0.246419 -0.94076
+ 7.36e+10Hz 0.244737 -0.941164
+ 7.37e+10Hz 0.243054 -0.941566
+ 7.38e+10Hz 0.24137 -0.941964
+ 7.39e+10Hz 0.239686 -0.94236
+ 7.4e+10Hz 0.238001 -0.942753
+ 7.41e+10Hz 0.236315 -0.943143
+ 7.42e+10Hz 0.234629 -0.943529
+ 7.43e+10Hz 0.232943 -0.943913
+ 7.44e+10Hz 0.231255 -0.944295
+ 7.45e+10Hz 0.229568 -0.944673
+ 7.46e+10Hz 0.227879 -0.945048
+ 7.47e+10Hz 0.22619 -0.94542
+ 7.48e+10Hz 0.2245 -0.94579
+ 7.49e+10Hz 0.22281 -0.946156
+ 7.5e+10Hz 0.221119 -0.94652
+ 7.51e+10Hz 0.219427 -0.94688
+ 7.52e+10Hz 0.217735 -0.947238
+ 7.53e+10Hz 0.216042 -0.947592
+ 7.54e+10Hz 0.214348 -0.947944
+ 7.55e+10Hz 0.212654 -0.948293
+ 7.56e+10Hz 0.210959 -0.948638
+ 7.57e+10Hz 0.209263 -0.948981
+ 7.58e+10Hz 0.207567 -0.949321
+ 7.59e+10Hz 0.20587 -0.949657
+ 7.6e+10Hz 0.204172 -0.949991
+ 7.61e+10Hz 0.202474 -0.950322
+ 7.62e+10Hz 0.200775 -0.950649
+ 7.63e+10Hz 0.199076 -0.950974
+ 7.64e+10Hz 0.197376 -0.951295
+ 7.65e+10Hz 0.195675 -0.951614
+ 7.66e+10Hz 0.193973 -0.951929
+ 7.67e+10Hz 0.192271 -0.952241
+ 7.68e+10Hz 0.190569 -0.952551
+ 7.69e+10Hz 0.188865 -0.952857
+ 7.7e+10Hz 0.187161 -0.95316
+ 7.71e+10Hz 0.185457 -0.953459
+ 7.72e+10Hz 0.183751 -0.953756
+ 7.73e+10Hz 0.182045 -0.95405
+ 7.74e+10Hz 0.180339 -0.95434
+ 7.75e+10Hz 0.178632 -0.954627
+ 7.76e+10Hz 0.176924 -0.954911
+ 7.77e+10Hz 0.175216 -0.955192
+ 7.78e+10Hz 0.173507 -0.95547
+ 7.79e+10Hz 0.171797 -0.955744
+ 7.8e+10Hz 0.170087 -0.956015
+ 7.81e+10Hz 0.168377 -0.956283
+ 7.82e+10Hz 0.166666 -0.956548
+ 7.83e+10Hz 0.164954 -0.95681
+ 7.84e+10Hz 0.163241 -0.957068
+ 7.85e+10Hz 0.161529 -0.957323
+ 7.86e+10Hz 0.159815 -0.957574
+ 7.87e+10Hz 0.158102 -0.957823
+ 7.88e+10Hz 0.156387 -0.958068
+ 7.89e+10Hz 0.154672 -0.958309
+ 7.9e+10Hz 0.152957 -0.958548
+ 7.91e+10Hz 0.151241 -0.958783
+ 7.92e+10Hz 0.149525 -0.959014
+ 7.93e+10Hz 0.147809 -0.959243
+ 7.94e+10Hz 0.146092 -0.959468
+ 7.95e+10Hz 0.144374 -0.959689
+ 7.96e+10Hz 0.142656 -0.959907
+ 7.97e+10Hz 0.140938 -0.960122
+ 7.98e+10Hz 0.139219 -0.960334
+ 7.99e+10Hz 0.137501 -0.960542
+ 8e+10Hz 0.135781 -0.960746
+ 8.01e+10Hz 0.134062 -0.960947
+ 8.02e+10Hz 0.132342 -0.961145
+ 8.03e+10Hz 0.130622 -0.961339
+ 8.04e+10Hz 0.128901 -0.96153
+ 8.05e+10Hz 0.127181 -0.961718
+ 8.06e+10Hz 0.12546 -0.961902
+ 8.07e+10Hz 0.123739 -0.962082
+ 8.08e+10Hz 0.122017 -0.962259
+ 8.09e+10Hz 0.120296 -0.962433
+ 8.1e+10Hz 0.118574 -0.962603
+ 8.11e+10Hz 0.116852 -0.96277
+ 8.12e+10Hz 0.11513 -0.962933
+ 8.13e+10Hz 0.113408 -0.963093
+ 8.14e+10Hz 0.111686 -0.963249
+ 8.15e+10Hz 0.109964 -0.963402
+ 8.16e+10Hz 0.108242 -0.963552
+ 8.17e+10Hz 0.10652 -0.963698
+ 8.18e+10Hz 0.104797 -0.96384
+ 8.19e+10Hz 0.103075 -0.963979
+ 8.2e+10Hz 0.101353 -0.964114
+ 8.21e+10Hz 0.0996305 -0.964247
+ 8.22e+10Hz 0.0979084 -0.964375
+ 8.23e+10Hz 0.0961863 -0.9645
+ 8.24e+10Hz 0.0944643 -0.964622
+ 8.25e+10Hz 0.0927424 -0.96474
+ 8.26e+10Hz 0.0910206 -0.964855
+ 8.27e+10Hz 0.089299 -0.964966
+ 8.28e+10Hz 0.0875776 -0.965074
+ 8.29e+10Hz 0.0858563 -0.965179
+ 8.3e+10Hz 0.0841353 -0.96528
+ 8.31e+10Hz 0.0824144 -0.965377
+ 8.32e+10Hz 0.0806938 -0.965472
+ 8.33e+10Hz 0.0789735 -0.965562
+ 8.34e+10Hz 0.0772534 -0.96565
+ 8.35e+10Hz 0.0755336 -0.965734
+ 8.36e+10Hz 0.0738141 -0.965815
+ 8.37e+10Hz 0.0720949 -0.965892
+ 8.38e+10Hz 0.070376 -0.965966
+ 8.39e+10Hz 0.0686576 -0.966036
+ 8.4e+10Hz 0.0669394 -0.966103
+ 8.41e+10Hz 0.0652217 -0.966167
+ 8.42e+10Hz 0.0635043 -0.966228
+ 8.43e+10Hz 0.0617874 -0.966285
+ 8.44e+10Hz 0.0600708 -0.966339
+ 8.45e+10Hz 0.0583547 -0.966389
+ 8.46e+10Hz 0.0566391 -0.966437
+ 8.47e+10Hz 0.0549239 -0.966481
+ 8.48e+10Hz 0.0532092 -0.966521
+ 8.49e+10Hz 0.051495 -0.966559
+ 8.5e+10Hz 0.0497813 -0.966593
+ 8.51e+10Hz 0.0480681 -0.966624
+ 8.52e+10Hz 0.0463554 -0.966652
+ 8.53e+10Hz 0.0446432 -0.966677
+ 8.54e+10Hz 0.0429316 -0.966698
+ 8.55e+10Hz 0.0412206 -0.966716
+ 8.56e+10Hz 0.0395101 -0.966731
+ 8.57e+10Hz 0.0378002 -0.966743
+ 8.58e+10Hz 0.0360908 -0.966752
+ 8.59e+10Hz 0.0343821 -0.966758
+ 8.6e+10Hz 0.0326739 -0.96676
+ 8.61e+10Hz 0.0309664 -0.96676
+ 8.62e+10Hz 0.0292595 -0.966756
+ 8.63e+10Hz 0.0275532 -0.966749
+ 8.64e+10Hz 0.0258475 -0.966739
+ 8.65e+10Hz 0.0241425 -0.966727
+ 8.66e+10Hz 0.0224381 -0.966711
+ 8.67e+10Hz 0.0207344 -0.966692
+ 8.68e+10Hz 0.0190313 -0.96667
+ 8.69e+10Hz 0.0173289 -0.966645
+ 8.7e+10Hz 0.0156271 -0.966617
+ 8.71e+10Hz 0.013926 -0.966586
+ 8.72e+10Hz 0.0122256 -0.966552
+ 8.73e+10Hz 0.0105259 -0.966516
+ 8.74e+10Hz 0.00882678 -0.966476
+ 8.75e+10Hz 0.0071284 -0.966433
+ 8.76e+10Hz 0.0054307 -0.966388
+ 8.77e+10Hz 0.00373368 -0.966339
+ 8.78e+10Hz 0.00203736 -0.966288
+ 8.79e+10Hz 0.000341723 -0.966234
+ 8.8e+10Hz -0.00135322 -0.966176
+ 8.81e+10Hz -0.00304746 -0.966116
+ 8.82e+10Hz -0.00474101 -0.966054
+ 8.83e+10Hz -0.00643386 -0.965988
+ 8.84e+10Hz -0.00812602 -0.96592
+ 8.85e+10Hz -0.00981748 -0.965848
+ 8.86e+10Hz -0.0115082 -0.965774
+ 8.87e+10Hz -0.0131983 -0.965698
+ 8.88e+10Hz -0.0148877 -0.965618
+ 8.89e+10Hz -0.0165763 -0.965536
+ 8.9e+10Hz -0.0182643 -0.965451
+ 8.91e+10Hz -0.0199516 -0.965363
+ 8.92e+10Hz -0.0216382 -0.965272
+ 8.93e+10Hz -0.023324 -0.965179
+ 8.94e+10Hz -0.0250092 -0.965083
+ 8.95e+10Hz -0.0266937 -0.964984
+ 8.96e+10Hz -0.0283775 -0.964883
+ 8.97e+10Hz -0.0300607 -0.964778
+ 8.98e+10Hz -0.0317431 -0.964672
+ 8.99e+10Hz -0.0334249 -0.964562
+ 9e+10Hz -0.0351059 -0.96445
+ 9.01e+10Hz -0.0367863 -0.964335
+ 9.02e+10Hz -0.038466 -0.964217
+ 9.03e+10Hz -0.040145 -0.964097
+ 9.04e+10Hz -0.0418234 -0.963975
+ 9.05e+10Hz -0.0435011 -0.963849
+ 9.06e+10Hz -0.0451781 -0.963721
+ 9.07e+10Hz -0.0468544 -0.96359
+ 9.08e+10Hz -0.0485301 -0.963457
+ 9.09e+10Hz -0.0502051 -0.963321
+ 9.1e+10Hz -0.0518795 -0.963183
+ 9.11e+10Hz -0.0535531 -0.963041
+ 9.12e+10Hz -0.0552262 -0.962898
+ 9.13e+10Hz -0.0568985 -0.962751
+ 9.14e+10Hz -0.0585702 -0.962602
+ 9.15e+10Hz -0.0602413 -0.962451
+ 9.16e+10Hz -0.0619117 -0.962297
+ 9.17e+10Hz -0.0635815 -0.96214
+ 9.18e+10Hz -0.0652506 -0.961981
+ 9.19e+10Hz -0.066919 -0.961819
+ 9.2e+10Hz -0.0685869 -0.961655
+ 9.21e+10Hz -0.070254 -0.961488
+ 9.22e+10Hz -0.0719206 -0.961318
+ 9.23e+10Hz -0.0735865 -0.961146
+ 9.24e+10Hz -0.0752517 -0.960971
+ 9.25e+10Hz -0.0769163 -0.960794
+ 9.26e+10Hz -0.0785803 -0.960615
+ 9.27e+10Hz -0.0802437 -0.960432
+ 9.28e+10Hz -0.0819064 -0.960247
+ 9.29e+10Hz -0.0835684 -0.96006
+ 9.3e+10Hz -0.0852299 -0.95987
+ 9.31e+10Hz -0.0868907 -0.959678
+ 9.32e+10Hz -0.0885509 -0.959483
+ 9.33e+10Hz -0.0902104 -0.959285
+ 9.34e+10Hz -0.0918693 -0.959085
+ 9.35e+10Hz -0.0935276 -0.958883
+ 9.36e+10Hz -0.0951852 -0.958678
+ 9.37e+10Hz -0.0968422 -0.95847
+ 9.38e+10Hz -0.0984986 -0.95826
+ 9.39e+10Hz -0.100154 -0.958047
+ 9.4e+10Hz -0.101809 -0.957832
+ 9.41e+10Hz -0.103464 -0.957614
+ 9.42e+10Hz -0.105118 -0.957394
+ 9.43e+10Hz -0.106771 -0.957172
+ 9.44e+10Hz -0.108424 -0.956946
+ 9.45e+10Hz -0.110076 -0.956719
+ 9.46e+10Hz -0.111727 -0.956488
+ 9.47e+10Hz -0.113377 -0.956256
+ 9.48e+10Hz -0.115027 -0.95602
+ 9.49e+10Hz -0.116677 -0.955783
+ 9.5e+10Hz -0.118326 -0.955543
+ 9.51e+10Hz -0.119974 -0.9553
+ 9.52e+10Hz -0.121621 -0.955055
+ 9.53e+10Hz -0.123268 -0.954807
+ 9.54e+10Hz -0.124914 -0.954557
+ 9.55e+10Hz -0.12656 -0.954304
+ 9.56e+10Hz -0.128205 -0.954049
+ 9.57e+10Hz -0.129849 -0.953791
+ 9.58e+10Hz -0.131492 -0.953531
+ 9.59e+10Hz -0.133135 -0.953269
+ 9.6e+10Hz -0.134777 -0.953004
+ 9.61e+10Hz -0.136419 -0.952736
+ 9.62e+10Hz -0.13806 -0.952466
+ 9.63e+10Hz -0.1397 -0.952194
+ 9.64e+10Hz -0.14134 -0.951919
+ 9.65e+10Hz -0.142979 -0.951642
+ 9.66e+10Hz -0.144617 -0.951362
+ 9.67e+10Hz -0.146255 -0.95108
+ 9.68e+10Hz -0.147892 -0.950795
+ 9.69e+10Hz -0.149528 -0.950508
+ 9.7e+10Hz -0.151164 -0.950219
+ 9.71e+10Hz -0.152799 -0.949927
+ 9.72e+10Hz -0.154433 -0.949633
+ 9.73e+10Hz -0.156067 -0.949336
+ 9.74e+10Hz -0.1577 -0.949037
+ 9.75e+10Hz -0.159332 -0.948735
+ 9.76e+10Hz -0.160964 -0.948431
+ 9.77e+10Hz -0.162595 -0.948125
+ 9.78e+10Hz -0.164225 -0.947816
+ 9.79e+10Hz -0.165855 -0.947505
+ 9.8e+10Hz -0.167484 -0.947191
+ 9.81e+10Hz -0.169112 -0.946875
+ 9.82e+10Hz -0.17074 -0.946557
+ 9.83e+10Hz -0.172367 -0.946236
+ 9.84e+10Hz -0.173993 -0.945913
+ 9.85e+10Hz -0.175619 -0.945588
+ 9.86e+10Hz -0.177244 -0.94526
+ 9.87e+10Hz -0.178868 -0.94493
+ 9.88e+10Hz -0.180492 -0.944598
+ 9.89e+10Hz -0.182115 -0.944263
+ 9.9e+10Hz -0.183737 -0.943926
+ 9.91e+10Hz -0.185359 -0.943586
+ 9.92e+10Hz -0.18698 -0.943244
+ 9.93e+10Hz -0.1886 -0.9429
+ 9.94e+10Hz -0.19022 -0.942554
+ 9.95e+10Hz -0.191839 -0.942205
+ 9.96e+10Hz -0.193458 -0.941854
+ 9.97e+10Hz -0.195076 -0.941501
+ 9.98e+10Hz -0.196693 -0.941145
+ 9.99e+10Hz -0.19831 -0.940787
+ 1e+11Hz -0.199926 -0.940427
+ 1.001e+11Hz -0.201541 -0.940064
+ 1.002e+11Hz -0.203156 -0.939699
+ 1.003e+11Hz -0.20477 -0.939332
+ 1.004e+11Hz -0.206384 -0.938962
+ 1.005e+11Hz -0.207997 -0.938591
+ 1.006e+11Hz -0.209609 -0.938217
+ 1.007e+11Hz -0.211221 -0.93784
+ 1.008e+11Hz -0.212832 -0.937462
+ 1.009e+11Hz -0.214443 -0.937081
+ 1.01e+11Hz -0.216053 -0.936698
+ 1.011e+11Hz -0.217662 -0.936312
+ 1.012e+11Hz -0.219271 -0.935925
+ 1.013e+11Hz -0.22088 -0.935535
+ 1.014e+11Hz -0.222488 -0.935143
+ 1.015e+11Hz -0.224095 -0.934748
+ 1.016e+11Hz -0.225702 -0.934351
+ 1.017e+11Hz -0.227308 -0.933952
+ 1.018e+11Hz -0.228914 -0.933551
+ 1.019e+11Hz -0.230519 -0.933148
+ 1.02e+11Hz -0.232124 -0.932742
+ 1.021e+11Hz -0.233728 -0.932334
+ 1.022e+11Hz -0.235332 -0.931924
+ 1.023e+11Hz -0.236935 -0.931511
+ 1.024e+11Hz -0.238538 -0.931096
+ 1.025e+11Hz -0.24014 -0.930679
+ 1.026e+11Hz -0.241742 -0.930259
+ 1.027e+11Hz -0.243343 -0.929838
+ 1.028e+11Hz -0.244944 -0.929414
+ 1.029e+11Hz -0.246544 -0.928988
+ 1.03e+11Hz -0.248145 -0.928559
+ 1.031e+11Hz -0.249744 -0.928128
+ 1.032e+11Hz -0.251343 -0.927695
+ 1.033e+11Hz -0.252942 -0.92726
+ 1.034e+11Hz -0.25454 -0.926822
+ 1.035e+11Hz -0.256138 -0.926382
+ 1.036e+11Hz -0.257736 -0.925939
+ 1.037e+11Hz -0.259333 -0.925495
+ 1.038e+11Hz -0.26093 -0.925048
+ 1.039e+11Hz -0.262526 -0.924598
+ 1.04e+11Hz -0.264122 -0.924146
+ 1.041e+11Hz -0.265718 -0.923692
+ 1.042e+11Hz -0.267313 -0.923236
+ 1.043e+11Hz -0.268908 -0.922777
+ 1.044e+11Hz -0.270503 -0.922316
+ 1.045e+11Hz -0.272097 -0.921852
+ 1.046e+11Hz -0.273691 -0.921386
+ 1.047e+11Hz -0.275285 -0.920918
+ 1.048e+11Hz -0.276878 -0.920447
+ 1.049e+11Hz -0.278471 -0.919974
+ 1.05e+11Hz -0.280064 -0.919498
+ 1.051e+11Hz -0.281656 -0.91902
+ 1.052e+11Hz -0.283248 -0.918539
+ 1.053e+11Hz -0.28484 -0.918056
+ 1.054e+11Hz -0.286431 -0.917571
+ 1.055e+11Hz -0.288022 -0.917083
+ 1.056e+11Hz -0.289613 -0.916592
+ 1.057e+11Hz -0.291203 -0.916099
+ 1.058e+11Hz -0.292793 -0.915604
+ 1.059e+11Hz -0.294383 -0.915106
+ 1.06e+11Hz -0.295973 -0.914605
+ 1.061e+11Hz -0.297562 -0.914102
+ 1.062e+11Hz -0.299151 -0.913596
+ 1.063e+11Hz -0.30074 -0.913088
+ 1.064e+11Hz -0.302328 -0.912577
+ 1.065e+11Hz -0.303916 -0.912063
+ 1.066e+11Hz -0.305504 -0.911547
+ 1.067e+11Hz -0.307091 -0.911028
+ 1.068e+11Hz -0.308678 -0.910507
+ 1.069e+11Hz -0.310265 -0.909983
+ 1.07e+11Hz -0.311852 -0.909456
+ 1.071e+11Hz -0.313438 -0.908926
+ 1.072e+11Hz -0.315024 -0.908394
+ 1.073e+11Hz -0.316609 -0.907859
+ 1.074e+11Hz -0.318195 -0.907321
+ 1.075e+11Hz -0.31978 -0.906781
+ 1.076e+11Hz -0.321364 -0.906238
+ 1.077e+11Hz -0.322948 -0.905692
+ 1.078e+11Hz -0.324532 -0.905143
+ 1.079e+11Hz -0.326116 -0.904592
+ 1.08e+11Hz -0.327699 -0.904037
+ 1.081e+11Hz -0.329282 -0.90348
+ 1.082e+11Hz -0.330864 -0.90292
+ 1.083e+11Hz -0.332446 -0.902357
+ 1.084e+11Hz -0.334028 -0.901791
+ 1.085e+11Hz -0.335609 -0.901222
+ 1.086e+11Hz -0.33719 -0.900651
+ 1.087e+11Hz -0.33877 -0.900076
+ 1.088e+11Hz -0.34035 -0.899499
+ 1.089e+11Hz -0.34193 -0.898919
+ 1.09e+11Hz -0.343509 -0.898335
+ 1.091e+11Hz -0.345087 -0.897749
+ 1.092e+11Hz -0.346665 -0.89716
+ 1.093e+11Hz -0.348243 -0.896568
+ 1.094e+11Hz -0.34982 -0.895972
+ 1.095e+11Hz -0.351396 -0.895374
+ 1.096e+11Hz -0.352972 -0.894773
+ 1.097e+11Hz -0.354548 -0.894169
+ 1.098e+11Hz -0.356122 -0.893562
+ 1.099e+11Hz -0.357697 -0.892951
+ 1.1e+11Hz -0.35927 -0.892338
+ 1.101e+11Hz -0.360844 -0.891721
+ 1.102e+11Hz -0.362416 -0.891102
+ 1.103e+11Hz -0.363988 -0.890479
+ 1.104e+11Hz -0.365559 -0.889854
+ 1.105e+11Hz -0.367129 -0.889225
+ 1.106e+11Hz -0.368699 -0.888593
+ 1.107e+11Hz -0.370268 -0.887958
+ 1.108e+11Hz -0.371837 -0.88732
+ 1.109e+11Hz -0.373404 -0.886679
+ 1.11e+11Hz -0.374971 -0.886034
+ 1.111e+11Hz -0.376537 -0.885387
+ 1.112e+11Hz -0.378103 -0.884736
+ 1.113e+11Hz -0.379667 -0.884082
+ 1.114e+11Hz -0.381231 -0.883425
+ 1.115e+11Hz -0.382794 -0.882765
+ 1.116e+11Hz -0.384356 -0.882102
+ 1.117e+11Hz -0.385917 -0.881436
+ 1.118e+11Hz -0.387477 -0.880766
+ 1.119e+11Hz -0.389036 -0.880093
+ 1.12e+11Hz -0.390594 -0.879418
+ 1.121e+11Hz -0.392152 -0.878739
+ 1.122e+11Hz -0.393708 -0.878056
+ 1.123e+11Hz -0.395264 -0.877371
+ 1.124e+11Hz -0.396818 -0.876682
+ 1.125e+11Hz -0.398371 -0.875991
+ 1.126e+11Hz -0.399924 -0.875296
+ 1.127e+11Hz -0.401475 -0.874598
+ 1.128e+11Hz -0.403025 -0.873897
+ 1.129e+11Hz -0.404574 -0.873192
+ 1.13e+11Hz -0.406122 -0.872485
+ 1.131e+11Hz -0.407669 -0.871774
+ 1.132e+11Hz -0.409215 -0.87106
+ 1.133e+11Hz -0.410759 -0.870343
+ 1.134e+11Hz -0.412302 -0.869623
+ 1.135e+11Hz -0.413845 -0.8689
+ 1.136e+11Hz -0.415385 -0.868174
+ 1.137e+11Hz -0.416925 -0.867444
+ 1.138e+11Hz -0.418463 -0.866711
+ 1.139e+11Hz -0.42 -0.865976
+ 1.14e+11Hz -0.421536 -0.865237
+ 1.141e+11Hz -0.423071 -0.864495
+ 1.142e+11Hz -0.424604 -0.86375
+ 1.143e+11Hz -0.426136 -0.863002
+ 1.144e+11Hz -0.427666 -0.862251
+ 1.145e+11Hz -0.429195 -0.861496
+ 1.146e+11Hz -0.430723 -0.860739
+ 1.147e+11Hz -0.432249 -0.859979
+ 1.148e+11Hz -0.433774 -0.859215
+ 1.149e+11Hz -0.435298 -0.858449
+ 1.15e+11Hz -0.43682 -0.857679
+ 1.151e+11Hz -0.43834 -0.856907
+ 1.152e+11Hz -0.43986 -0.856131
+ 1.153e+11Hz -0.441377 -0.855353
+ 1.154e+11Hz -0.442893 -0.854571
+ 1.155e+11Hz -0.444408 -0.853786
+ 1.156e+11Hz -0.445921 -0.852999
+ 1.157e+11Hz -0.447433 -0.852209
+ 1.158e+11Hz -0.448943 -0.851415
+ 1.159e+11Hz -0.450451 -0.850619
+ 1.16e+11Hz -0.451958 -0.84982
+ 1.161e+11Hz -0.453464 -0.849018
+ 1.162e+11Hz -0.454967 -0.848213
+ 1.163e+11Hz -0.45647 -0.847405
+ 1.164e+11Hz -0.45797 -0.846594
+ 1.165e+11Hz -0.459469 -0.84578
+ 1.166e+11Hz -0.460967 -0.844964
+ 1.167e+11Hz -0.462462 -0.844144
+ 1.168e+11Hz -0.463956 -0.843322
+ 1.169e+11Hz -0.465449 -0.842497
+ 1.17e+11Hz -0.46694 -0.841669
+ 1.171e+11Hz -0.468429 -0.840839
+ 1.172e+11Hz -0.469917 -0.840005
+ 1.173e+11Hz -0.471402 -0.839169
+ 1.174e+11Hz -0.472887 -0.83833
+ 1.175e+11Hz -0.474369 -0.837488
+ 1.176e+11Hz -0.47585 -0.836644
+ 1.177e+11Hz -0.477329 -0.835797
+ 1.178e+11Hz -0.478807 -0.834947
+ 1.179e+11Hz -0.480282 -0.834094
+ 1.18e+11Hz -0.481756 -0.833239
+ 1.181e+11Hz -0.483229 -0.832381
+ 1.182e+11Hz -0.4847 -0.83152
+ 1.183e+11Hz -0.486169 -0.830657
+ 1.184e+11Hz -0.487636 -0.829791
+ 1.185e+11Hz -0.489101 -0.828923
+ 1.186e+11Hz -0.490565 -0.828051
+ 1.187e+11Hz -0.492027 -0.827177
+ 1.188e+11Hz -0.493488 -0.826301
+ 1.189e+11Hz -0.494947 -0.825422
+ 1.19e+11Hz -0.496404 -0.82454
+ 1.191e+11Hz -0.497859 -0.823656
+ 1.192e+11Hz -0.499312 -0.822769
+ 1.193e+11Hz -0.500764 -0.82188
+ 1.194e+11Hz -0.502214 -0.820988
+ 1.195e+11Hz -0.503663 -0.820093
+ 1.196e+11Hz -0.505109 -0.819196
+ 1.197e+11Hz -0.506554 -0.818296
+ 1.198e+11Hz -0.507998 -0.817394
+ 1.199e+11Hz -0.509439 -0.81649
+ 1.2e+11Hz -0.510879 -0.815582
+ 1.201e+11Hz -0.512317 -0.814673
+ 1.202e+11Hz -0.513753 -0.81376
+ 1.203e+11Hz -0.515188 -0.812846
+ 1.204e+11Hz -0.516621 -0.811928
+ 1.205e+11Hz -0.518052 -0.811009
+ 1.206e+11Hz -0.519482 -0.810086
+ 1.207e+11Hz -0.52091 -0.809162
+ 1.208e+11Hz -0.522336 -0.808235
+ 1.209e+11Hz -0.52376 -0.807305
+ 1.21e+11Hz -0.525183 -0.806373
+ 1.211e+11Hz -0.526604 -0.805438
+ 1.212e+11Hz -0.528023 -0.804501
+ 1.213e+11Hz -0.52944 -0.803562
+ 1.214e+11Hz -0.530856 -0.80262
+ 1.215e+11Hz -0.53227 -0.801675
+ 1.216e+11Hz -0.533683 -0.800729
+ 1.217e+11Hz -0.535093 -0.799779
+ 1.218e+11Hz -0.536502 -0.798827
+ 1.219e+11Hz -0.53791 -0.797873
+ 1.22e+11Hz -0.539315 -0.796917
+ 1.221e+11Hz -0.540719 -0.795958
+ 1.222e+11Hz -0.542121 -0.794996
+ 1.223e+11Hz -0.543522 -0.794032
+ 1.224e+11Hz -0.54492 -0.793066
+ 1.225e+11Hz -0.546317 -0.792097
+ 1.226e+11Hz -0.547713 -0.791126
+ 1.227e+11Hz -0.549106 -0.790152
+ 1.228e+11Hz -0.550498 -0.789176
+ 1.229e+11Hz -0.551888 -0.788197
+ 1.23e+11Hz -0.553277 -0.787216
+ 1.231e+11Hz -0.554663 -0.786233
+ 1.232e+11Hz -0.556048 -0.785247
+ 1.233e+11Hz -0.557432 -0.784258
+ 1.234e+11Hz -0.558813 -0.783268
+ 1.235e+11Hz -0.560193 -0.782274
+ 1.236e+11Hz -0.561571 -0.781279
+ 1.237e+11Hz -0.562948 -0.780281
+ 1.238e+11Hz -0.564322 -0.77928
+ 1.239e+11Hz -0.565695 -0.778277
+ 1.24e+11Hz -0.567066 -0.777271
+ 1.241e+11Hz -0.568436 -0.776264
+ 1.242e+11Hz -0.569803 -0.775253
+ 1.243e+11Hz -0.571169 -0.77424
+ 1.244e+11Hz -0.572533 -0.773225
+ 1.245e+11Hz -0.573896 -0.772208
+ 1.246e+11Hz -0.575256 -0.771187
+ 1.247e+11Hz -0.576615 -0.770165
+ 1.248e+11Hz -0.577972 -0.76914
+ 1.249e+11Hz -0.579327 -0.768112
+ 1.25e+11Hz -0.580681 -0.767082
+ 1.251e+11Hz -0.582032 -0.76605
+ 1.252e+11Hz -0.583382 -0.765015
+ 1.253e+11Hz -0.58473 -0.763978
+ 1.254e+11Hz -0.586076 -0.762938
+ 1.255e+11Hz -0.587421 -0.761896
+ 1.256e+11Hz -0.588763 -0.760851
+ 1.257e+11Hz -0.590104 -0.759804
+ 1.258e+11Hz -0.591443 -0.758754
+ 1.259e+11Hz -0.59278 -0.757702
+ 1.26e+11Hz -0.594115 -0.756648
+ 1.261e+11Hz -0.595448 -0.755591
+ 1.262e+11Hz -0.596779 -0.754531
+ 1.263e+11Hz -0.598109 -0.753469
+ 1.264e+11Hz -0.599436 -0.752405
+ 1.265e+11Hz -0.600762 -0.751338
+ 1.266e+11Hz -0.602086 -0.750269
+ 1.267e+11Hz -0.603407 -0.749197
+ 1.268e+11Hz -0.604727 -0.748123
+ 1.269e+11Hz -0.606045 -0.747047
+ 1.27e+11Hz -0.607361 -0.745968
+ 1.271e+11Hz -0.608675 -0.744886
+ 1.272e+11Hz -0.609987 -0.743802
+ 1.273e+11Hz -0.611297 -0.742716
+ 1.274e+11Hz -0.612605 -0.741627
+ 1.275e+11Hz -0.613911 -0.740536
+ 1.276e+11Hz -0.615215 -0.739443
+ 1.277e+11Hz -0.616517 -0.738347
+ 1.278e+11Hz -0.617817 -0.737248
+ 1.279e+11Hz -0.619114 -0.736147
+ 1.28e+11Hz -0.62041 -0.735044
+ 1.281e+11Hz -0.621704 -0.733938
+ 1.282e+11Hz -0.622996 -0.732831
+ 1.283e+11Hz -0.624285 -0.73172
+ 1.284e+11Hz -0.625573 -0.730607
+ 1.285e+11Hz -0.626858 -0.729492
+ 1.286e+11Hz -0.628141 -0.728375
+ 1.287e+11Hz -0.629422 -0.727255
+ 1.288e+11Hz -0.630701 -0.726133
+ 1.289e+11Hz -0.631978 -0.725008
+ 1.29e+11Hz -0.633253 -0.723881
+ 1.291e+11Hz -0.634525 -0.722752
+ 1.292e+11Hz -0.635795 -0.721621
+ 1.293e+11Hz -0.637064 -0.720487
+ 1.294e+11Hz -0.638329 -0.719351
+ 1.295e+11Hz -0.639593 -0.718212
+ 1.296e+11Hz -0.640855 -0.717072
+ 1.297e+11Hz -0.642114 -0.715929
+ 1.298e+11Hz -0.643371 -0.714783
+ 1.299e+11Hz -0.644626 -0.713636
+ 1.3e+11Hz -0.645878 -0.712486
+ 1.301e+11Hz -0.647129 -0.711334
+ 1.302e+11Hz -0.648377 -0.71018
+ 1.303e+11Hz -0.649623 -0.709024
+ 1.304e+11Hz -0.650866 -0.707865
+ 1.305e+11Hz -0.652108 -0.706704
+ 1.306e+11Hz -0.653347 -0.705542
+ 1.307e+11Hz -0.654583 -0.704376
+ 1.308e+11Hz -0.655818 -0.703209
+ 1.309e+11Hz -0.65705 -0.70204
+ 1.31e+11Hz -0.65828 -0.700868
+ 1.311e+11Hz -0.659507 -0.699695
+ 1.312e+11Hz -0.660732 -0.698519
+ 1.313e+11Hz -0.661955 -0.697341
+ 1.314e+11Hz -0.663175 -0.696161
+ 1.315e+11Hz -0.664394 -0.694979
+ 1.316e+11Hz -0.665609 -0.693795
+ 1.317e+11Hz -0.666823 -0.692609
+ 1.318e+11Hz -0.668034 -0.691421
+ 1.319e+11Hz -0.669243 -0.690231
+ 1.32e+11Hz -0.670449 -0.689039
+ 1.321e+11Hz -0.671654 -0.687845
+ 1.322e+11Hz -0.672855 -0.686648
+ 1.323e+11Hz -0.674055 -0.68545
+ 1.324e+11Hz -0.675252 -0.68425
+ 1.325e+11Hz -0.676447 -0.683048
+ 1.326e+11Hz -0.677639 -0.681844
+ 1.327e+11Hz -0.678829 -0.680639
+ 1.328e+11Hz -0.680017 -0.679431
+ 1.329e+11Hz -0.681202 -0.678221
+ 1.33e+11Hz -0.682385 -0.67701
+ 1.331e+11Hz -0.683565 -0.675796
+ 1.332e+11Hz -0.684744 -0.674581
+ 1.333e+11Hz -0.68592 -0.673364
+ 1.334e+11Hz -0.687093 -0.672145
+ 1.335e+11Hz -0.688264 -0.670925
+ 1.336e+11Hz -0.689433 -0.669702
+ 1.337e+11Hz -0.6906 -0.668478
+ 1.338e+11Hz -0.691764 -0.667252
+ 1.339e+11Hz -0.692926 -0.666024
+ 1.34e+11Hz -0.694085 -0.664794
+ 1.341e+11Hz -0.695243 -0.663563
+ 1.342e+11Hz -0.696397 -0.66233
+ 1.343e+11Hz -0.69755 -0.661095
+ 1.344e+11Hz -0.6987 -0.659858
+ 1.345e+11Hz -0.699848 -0.65862
+ 1.346e+11Hz -0.700994 -0.65738
+ 1.347e+11Hz -0.702137 -0.656138
+ 1.348e+11Hz -0.703278 -0.654895
+ 1.349e+11Hz -0.704417 -0.65365
+ 1.35e+11Hz -0.705554 -0.652403
+ 1.351e+11Hz -0.706688 -0.651155
+ 1.352e+11Hz -0.70782 -0.649905
+ 1.353e+11Hz -0.708949 -0.648653
+ 1.354e+11Hz -0.710077 -0.6474
+ 1.355e+11Hz -0.711202 -0.646145
+ 1.356e+11Hz -0.712325 -0.644888
+ 1.357e+11Hz -0.713446 -0.64363
+ 1.358e+11Hz -0.714564 -0.642371
+ 1.359e+11Hz -0.715681 -0.641109
+ 1.36e+11Hz -0.716795 -0.639846
+ 1.361e+11Hz -0.717906 -0.638582
+ 1.362e+11Hz -0.719016 -0.637316
+ 1.363e+11Hz -0.720124 -0.636048
+ 1.364e+11Hz -0.721229 -0.634779
+ 1.365e+11Hz -0.722332 -0.633508
+ 1.366e+11Hz -0.723433 -0.632236
+ 1.367e+11Hz -0.724532 -0.630962
+ 1.368e+11Hz -0.725628 -0.629686
+ 1.369e+11Hz -0.726723 -0.628409
+ 1.37e+11Hz -0.727815 -0.62713
+ 1.371e+11Hz -0.728905 -0.62585
+ 1.372e+11Hz -0.729993 -0.624569
+ 1.373e+11Hz -0.731079 -0.623285
+ 1.374e+11Hz -0.732163 -0.622001
+ 1.375e+11Hz -0.733245 -0.620714
+ 1.376e+11Hz -0.734325 -0.619426
+ 1.377e+11Hz -0.735402 -0.618137
+ 1.378e+11Hz -0.736478 -0.616846
+ 1.379e+11Hz -0.737551 -0.615553
+ 1.38e+11Hz -0.738623 -0.614259
+ 1.381e+11Hz -0.739692 -0.612964
+ 1.382e+11Hz -0.740759 -0.611667
+ 1.383e+11Hz -0.741825 -0.610368
+ 1.384e+11Hz -0.742888 -0.609068
+ 1.385e+11Hz -0.743949 -0.607766
+ 1.386e+11Hz -0.745008 -0.606463
+ 1.387e+11Hz -0.746065 -0.605158
+ 1.388e+11Hz -0.74712 -0.603851
+ 1.389e+11Hz -0.748174 -0.602544
+ 1.39e+11Hz -0.749225 -0.601234
+ 1.391e+11Hz -0.750274 -0.599923
+ 1.392e+11Hz -0.751321 -0.59861
+ 1.393e+11Hz -0.752366 -0.597296
+ 1.394e+11Hz -0.753409 -0.59598
+ 1.395e+11Hz -0.754451 -0.594663
+ 1.396e+11Hz -0.75549 -0.593344
+ 1.397e+11Hz -0.756527 -0.592023
+ 1.398e+11Hz -0.757562 -0.590701
+ 1.399e+11Hz -0.758596 -0.589377
+ 1.4e+11Hz -0.759627 -0.588052
+ 1.401e+11Hz -0.760657 -0.586725
+ 1.402e+11Hz -0.761684 -0.585397
+ 1.403e+11Hz -0.76271 -0.584066
+ 1.404e+11Hz -0.763733 -0.582735
+ 1.405e+11Hz -0.764755 -0.581401
+ 1.406e+11Hz -0.765775 -0.580066
+ 1.407e+11Hz -0.766792 -0.578729
+ 1.408e+11Hz -0.767808 -0.577391
+ 1.409e+11Hz -0.768822 -0.576051
+ 1.41e+11Hz -0.769834 -0.57471
+ 1.411e+11Hz -0.770844 -0.573366
+ 1.412e+11Hz -0.771852 -0.572021
+ 1.413e+11Hz -0.772858 -0.570675
+ 1.414e+11Hz -0.773863 -0.569326
+ 1.415e+11Hz -0.774865 -0.567976
+ 1.416e+11Hz -0.775865 -0.566625
+ 1.417e+11Hz -0.776864 -0.565271
+ 1.418e+11Hz -0.77786 -0.563916
+ 1.419e+11Hz -0.778855 -0.562559
+ 1.42e+11Hz -0.779848 -0.561201
+ 1.421e+11Hz -0.780838 -0.55984
+ 1.422e+11Hz -0.781827 -0.558478
+ 1.423e+11Hz -0.782814 -0.557115
+ 1.424e+11Hz -0.783799 -0.555749
+ 1.425e+11Hz -0.784782 -0.554382
+ 1.426e+11Hz -0.785762 -0.553013
+ 1.427e+11Hz -0.786741 -0.551642
+ 1.428e+11Hz -0.787718 -0.55027
+ 1.429e+11Hz -0.788694 -0.548895
+ 1.43e+11Hz -0.789667 -0.547519
+ 1.431e+11Hz -0.790638 -0.546141
+ 1.432e+11Hz -0.791607 -0.544762
+ 1.433e+11Hz -0.792574 -0.54338
+ 1.434e+11Hz -0.793539 -0.541997
+ 1.435e+11Hz -0.794502 -0.540612
+ 1.436e+11Hz -0.795463 -0.539225
+ 1.437e+11Hz -0.796423 -0.537836
+ 1.438e+11Hz -0.79738 -0.536446
+ 1.439e+11Hz -0.798335 -0.535053
+ 1.44e+11Hz -0.799288 -0.533659
+ 1.441e+11Hz -0.800239 -0.532263
+ 1.442e+11Hz -0.801188 -0.530865
+ 1.443e+11Hz -0.802135 -0.529465
+ 1.444e+11Hz -0.80308 -0.528064
+ 1.445e+11Hz -0.804023 -0.52666
+ 1.446e+11Hz -0.804964 -0.525255
+ 1.447e+11Hz -0.805903 -0.523848
+ 1.448e+11Hz -0.806839 -0.522439
+ 1.449e+11Hz -0.807774 -0.521028
+ 1.45e+11Hz -0.808706 -0.519615
+ 1.451e+11Hz -0.809637 -0.5182
+ 1.452e+11Hz -0.810565 -0.516784
+ 1.453e+11Hz -0.811491 -0.515365
+ 1.454e+11Hz -0.812415 -0.513945
+ 1.455e+11Hz -0.813337 -0.512523
+ 1.456e+11Hz -0.814257 -0.511098
+ 1.457e+11Hz -0.815175 -0.509672
+ 1.458e+11Hz -0.81609 -0.508244
+ 1.459e+11Hz -0.817003 -0.506815
+ 1.46e+11Hz -0.817914 -0.505383
+ 1.461e+11Hz -0.818823 -0.503949
+ 1.462e+11Hz -0.81973 -0.502514
+ 1.463e+11Hz -0.820635 -0.501076
+ 1.464e+11Hz -0.821537 -0.499637
+ 1.465e+11Hz -0.822437 -0.498195
+ 1.466e+11Hz -0.823335 -0.496752
+ 1.467e+11Hz -0.824231 -0.495307
+ 1.468e+11Hz -0.825124 -0.49386
+ 1.469e+11Hz -0.826015 -0.492411
+ 1.47e+11Hz -0.826904 -0.49096
+ 1.471e+11Hz -0.827791 -0.489507
+ 1.472e+11Hz -0.828675 -0.488053
+ 1.473e+11Hz -0.829557 -0.486596
+ 1.474e+11Hz -0.830437 -0.485137
+ 1.475e+11Hz -0.831314 -0.483677
+ 1.476e+11Hz -0.83219 -0.482214
+ 1.477e+11Hz -0.833062 -0.48075
+ 1.478e+11Hz -0.833933 -0.479284
+ 1.479e+11Hz -0.834801 -0.477816
+ 1.48e+11Hz -0.835667 -0.476346
+ 1.481e+11Hz -0.83653 -0.474874
+ 1.482e+11Hz -0.837391 -0.4734
+ 1.483e+11Hz -0.83825 -0.471924
+ 1.484e+11Hz -0.839106 -0.470446
+ 1.485e+11Hz -0.83996 -0.468967
+ 1.486e+11Hz -0.840811 -0.467485
+ 1.487e+11Hz -0.84166 -0.466002
+ 1.488e+11Hz -0.842507 -0.464516
+ 1.489e+11Hz -0.843351 -0.463029
+ 1.49e+11Hz -0.844193 -0.46154
+ 1.491e+11Hz -0.845032 -0.460049
+ 1.492e+11Hz -0.845869 -0.458556
+ 1.493e+11Hz -0.846703 -0.457061
+ 1.494e+11Hz -0.847535 -0.455564
+ 1.495e+11Hz -0.848364 -0.454065
+ 1.496e+11Hz -0.849191 -0.452565
+ 1.497e+11Hz -0.850015 -0.451062
+ 1.498e+11Hz -0.850837 -0.449558
+ 1.499e+11Hz -0.851656 -0.448052
+ 1.5e+11Hz -0.852473 -0.446544
+ 1.501e+11Hz -0.853287 -0.445034
+ 1.502e+11Hz -0.854099 -0.443522
+ 1.503e+11Hz -0.854908 -0.442008
+ 1.504e+11Hz -0.855715 -0.440493
+ 1.505e+11Hz -0.856518 -0.438975
+ 1.506e+11Hz -0.85732 -0.437456
+ 1.507e+11Hz -0.858118 -0.435934
+ 1.508e+11Hz -0.858915 -0.434411
+ 1.509e+11Hz -0.859708 -0.432886
+ 1.51e+11Hz -0.860499 -0.43136
+ 1.511e+11Hz -0.861287 -0.429831
+ 1.512e+11Hz -0.862073 -0.4283
+ 1.513e+11Hz -0.862856 -0.426768
+ 1.514e+11Hz -0.863636 -0.425234
+ 1.515e+11Hz -0.864413 -0.423698
+ 1.516e+11Hz -0.865188 -0.42216
+ 1.517e+11Hz -0.865961 -0.42062
+ 1.518e+11Hz -0.86673 -0.419079
+ 1.519e+11Hz -0.867497 -0.417535
+ 1.52e+11Hz -0.868261 -0.41599
+ 1.521e+11Hz -0.869022 -0.414443
+ 1.522e+11Hz -0.869781 -0.412894
+ 1.523e+11Hz -0.870537 -0.411344
+ 1.524e+11Hz -0.87129 -0.409791
+ 1.525e+11Hz -0.87204 -0.408237
+ 1.526e+11Hz -0.872788 -0.406681
+ 1.527e+11Hz -0.873532 -0.405123
+ 1.528e+11Hz -0.874274 -0.403564
+ 1.529e+11Hz -0.875013 -0.402002
+ 1.53e+11Hz -0.87575 -0.400439
+ 1.531e+11Hz -0.876483 -0.398874
+ 1.532e+11Hz -0.877214 -0.397307
+ 1.533e+11Hz -0.877942 -0.395739
+ 1.534e+11Hz -0.878667 -0.394168
+ 1.535e+11Hz -0.879389 -0.392596
+ 1.536e+11Hz -0.880108 -0.391023
+ 1.537e+11Hz -0.880824 -0.389447
+ 1.538e+11Hz -0.881538 -0.38787
+ 1.539e+11Hz -0.882248 -0.386291
+ 1.54e+11Hz -0.882956 -0.38471
+ 1.541e+11Hz -0.883661 -0.383127
+ 1.542e+11Hz -0.884363 -0.381543
+ 1.543e+11Hz -0.885061 -0.379957
+ 1.544e+11Hz -0.885757 -0.37837
+ 1.545e+11Hz -0.88645 -0.37678
+ 1.546e+11Hz -0.88714 -0.375189
+ 1.547e+11Hz -0.887827 -0.373596
+ 1.548e+11Hz -0.888511 -0.372002
+ 1.549e+11Hz -0.889192 -0.370406
+ 1.55e+11Hz -0.88987 -0.368808
+ 1.551e+11Hz -0.890545 -0.367208
+ 1.552e+11Hz -0.891216 -0.365607
+ 1.553e+11Hz -0.891885 -0.364005
+ 1.554e+11Hz -0.892551 -0.3624
+ 1.555e+11Hz -0.893214 -0.360794
+ 1.556e+11Hz -0.893873 -0.359186
+ 1.557e+11Hz -0.89453 -0.357577
+ 1.558e+11Hz -0.895183 -0.355966
+ 1.559e+11Hz -0.895833 -0.354353
+ 1.56e+11Hz -0.89648 -0.352739
+ 1.561e+11Hz -0.897124 -0.351123
+ 1.562e+11Hz -0.897765 -0.349506
+ 1.563e+11Hz -0.898403 -0.347887
+ 1.564e+11Hz -0.899037 -0.346267
+ 1.565e+11Hz -0.899669 -0.344645
+ 1.566e+11Hz -0.900297 -0.343021
+ 1.567e+11Hz -0.900922 -0.341396
+ 1.568e+11Hz -0.901544 -0.339769
+ 1.569e+11Hz -0.902162 -0.338141
+ 1.57e+11Hz -0.902777 -0.336511
+ 1.571e+11Hz -0.903389 -0.33488
+ 1.572e+11Hz -0.903998 -0.333248
+ 1.573e+11Hz -0.904604 -0.331613
+ 1.574e+11Hz -0.905206 -0.329978
+ 1.575e+11Hz -0.905805 -0.328341
+ 1.576e+11Hz -0.906401 -0.326702
+ 1.577e+11Hz -0.906993 -0.325062
+ 1.578e+11Hz -0.907582 -0.323421
+ 1.579e+11Hz -0.908168 -0.321778
+ 1.58e+11Hz -0.908751 -0.320134
+ 1.581e+11Hz -0.90933 -0.318488
+ 1.582e+11Hz -0.909905 -0.316841
+ 1.583e+11Hz -0.910478 -0.315193
+ 1.584e+11Hz -0.911047 -0.313543
+ 1.585e+11Hz -0.911613 -0.311892
+ 1.586e+11Hz -0.912175 -0.31024
+ 1.587e+11Hz -0.912734 -0.308586
+ 1.588e+11Hz -0.913289 -0.306931
+ 1.589e+11Hz -0.913841 -0.305275
+ 1.59e+11Hz -0.91439 -0.303618
+ 1.591e+11Hz -0.914935 -0.301959
+ 1.592e+11Hz -0.915477 -0.300299
+ 1.593e+11Hz -0.916016 -0.298638
+ 1.594e+11Hz -0.916551 -0.296975
+ 1.595e+11Hz -0.917082 -0.295312
+ 1.596e+11Hz -0.91761 -0.293647
+ 1.597e+11Hz -0.918135 -0.291981
+ 1.598e+11Hz -0.918656 -0.290314
+ 1.599e+11Hz -0.919173 -0.288645
+ 1.6e+11Hz -0.919688 -0.286976
+ 1.601e+11Hz -0.920198 -0.285305
+ 1.602e+11Hz -0.920705 -0.283634
+ 1.603e+11Hz -0.921209 -0.281961
+ 1.604e+11Hz -0.921709 -0.280287
+ 1.605e+11Hz -0.922206 -0.278613
+ 1.606e+11Hz -0.922699 -0.276937
+ 1.607e+11Hz -0.923189 -0.27526
+ 1.608e+11Hz -0.923675 -0.273582
+ 1.609e+11Hz -0.924157 -0.271903
+ 1.61e+11Hz -0.924636 -0.270223
+ 1.611e+11Hz -0.925112 -0.268543
+ 1.612e+11Hz -0.925584 -0.266861
+ 1.613e+11Hz -0.926052 -0.265178
+ 1.614e+11Hz -0.926517 -0.263495
+ 1.615e+11Hz -0.926979 -0.26181
+ 1.616e+11Hz -0.927436 -0.260125
+ 1.617e+11Hz -0.927891 -0.258439
+ 1.618e+11Hz -0.928341 -0.256752
+ 1.619e+11Hz -0.928788 -0.255064
+ 1.62e+11Hz -0.929232 -0.253376
+ 1.621e+11Hz -0.929672 -0.251686
+ 1.622e+11Hz -0.930109 -0.249996
+ 1.623e+11Hz -0.930542 -0.248305
+ 1.624e+11Hz -0.930971 -0.246614
+ 1.625e+11Hz -0.931397 -0.244921
+ 1.626e+11Hz -0.931819 -0.243228
+ 1.627e+11Hz -0.932238 -0.241534
+ 1.628e+11Hz -0.932653 -0.23984
+ 1.629e+11Hz -0.933065 -0.238145
+ 1.63e+11Hz -0.933473 -0.236449
+ 1.631e+11Hz -0.933877 -0.234752
+ 1.632e+11Hz -0.934278 -0.233055
+ 1.633e+11Hz -0.934676 -0.231358
+ 1.634e+11Hz -0.93507 -0.229659
+ 1.635e+11Hz -0.93546 -0.227961
+ 1.636e+11Hz -0.935847 -0.226261
+ 1.637e+11Hz -0.93623 -0.224561
+ 1.638e+11Hz -0.93661 -0.222861
+ 1.639e+11Hz -0.936986 -0.22116
+ 1.64e+11Hz -0.937359 -0.219458
+ 1.641e+11Hz -0.937728 -0.217756
+ 1.642e+11Hz -0.938094 -0.216054
+ 1.643e+11Hz -0.938456 -0.214351
+ 1.644e+11Hz -0.938815 -0.212648
+ 1.645e+11Hz -0.93917 -0.210944
+ 1.646e+11Hz -0.939522 -0.20924
+ 1.647e+11Hz -0.93987 -0.207535
+ 1.648e+11Hz -0.940215 -0.20583
+ 1.649e+11Hz -0.940557 -0.204125
+ 1.65e+11Hz -0.940894 -0.202419
+ 1.651e+11Hz -0.941229 -0.200713
+ 1.652e+11Hz -0.94156 -0.199006
+ 1.653e+11Hz -0.941887 -0.1973
+ 1.654e+11Hz -0.942211 -0.195593
+ 1.655e+11Hz -0.942532 -0.193885
+ 1.656e+11Hz -0.942849 -0.192177
+ 1.657e+11Hz -0.943163 -0.190469
+ 1.658e+11Hz -0.943473 -0.188761
+ 1.659e+11Hz -0.94378 -0.187053
+ 1.66e+11Hz -0.944084 -0.185344
+ 1.661e+11Hz -0.944384 -0.183635
+ 1.662e+11Hz -0.94468 -0.181925
+ 1.663e+11Hz -0.944974 -0.180216
+ 1.664e+11Hz -0.945264 -0.178506
+ 1.665e+11Hz -0.94555 -0.176796
+ 1.666e+11Hz -0.945834 -0.175086
+ 1.667e+11Hz -0.946113 -0.173376
+ 1.668e+11Hz -0.94639 -0.171665
+ 1.669e+11Hz -0.946663 -0.169954
+ 1.67e+11Hz -0.946933 -0.168244
+ 1.671e+11Hz -0.947199 -0.166533
+ 1.672e+11Hz -0.947463 -0.164821
+ 1.673e+11Hz -0.947722 -0.16311
+ 1.674e+11Hz -0.947979 -0.161398
+ 1.675e+11Hz -0.948232 -0.159687
+ 1.676e+11Hz -0.948482 -0.157975
+ 1.677e+11Hz -0.948729 -0.156263
+ 1.678e+11Hz -0.948972 -0.154551
+ 1.679e+11Hz -0.949212 -0.152839
+ 1.68e+11Hz -0.949449 -0.151127
+ 1.681e+11Hz -0.949683 -0.149414
+ 1.682e+11Hz -0.949913 -0.147702
+ 1.683e+11Hz -0.95014 -0.145989
+ 1.684e+11Hz -0.950364 -0.144277
+ 1.685e+11Hz -0.950584 -0.142564
+ 1.686e+11Hz -0.950802 -0.140851
+ 1.687e+11Hz -0.951016 -0.139138
+ 1.688e+11Hz -0.951227 -0.137426
+ 1.689e+11Hz -0.951434 -0.135713
+ 1.69e+11Hz -0.951639 -0.133999
+ 1.691e+11Hz -0.95184 -0.132286
+ 1.692e+11Hz -0.952038 -0.130573
+ 1.693e+11Hz -0.952233 -0.12886
+ 1.694e+11Hz -0.952424 -0.127147
+ 1.695e+11Hz -0.952613 -0.125433
+ 1.696e+11Hz -0.952798 -0.12372
+ 1.697e+11Hz -0.95298 -0.122007
+ 1.698e+11Hz -0.953159 -0.120293
+ 1.699e+11Hz -0.953335 -0.11858
+ 1.7e+11Hz -0.953507 -0.116866
+ 1.701e+11Hz -0.953677 -0.115153
+ 1.702e+11Hz -0.953843 -0.113439
+ 1.703e+11Hz -0.954006 -0.111726
+ 1.704e+11Hz -0.954166 -0.110012
+ 1.705e+11Hz -0.954323 -0.108299
+ 1.706e+11Hz -0.954476 -0.106585
+ 1.707e+11Hz -0.954627 -0.104871
+ 1.708e+11Hz -0.954774 -0.103158
+ 1.709e+11Hz -0.954918 -0.101444
+ 1.71e+11Hz -0.955059 -0.0997304
+ 1.711e+11Hz -0.955197 -0.0980168
+ 1.712e+11Hz -0.955332 -0.0963031
+ 1.713e+11Hz -0.955463 -0.0945895
+ 1.714e+11Hz -0.955592 -0.0928758
+ 1.715e+11Hz -0.955717 -0.0911622
+ 1.716e+11Hz -0.955839 -0.0894486
+ 1.717e+11Hz -0.955958 -0.087735
+ 1.718e+11Hz -0.956074 -0.0860214
+ 1.719e+11Hz -0.956187 -0.0843078
+ 1.72e+11Hz -0.956297 -0.0825942
+ 1.721e+11Hz -0.956403 -0.0808807
+ 1.722e+11Hz -0.956506 -0.0791672
+ 1.723e+11Hz -0.956607 -0.0774537
+ 1.724e+11Hz -0.956704 -0.0757403
+ 1.725e+11Hz -0.956798 -0.0740269
+ 1.726e+11Hz -0.956888 -0.0723135
+ 1.727e+11Hz -0.956976 -0.0706002
+ 1.728e+11Hz -0.957061 -0.0688869
+ 1.729e+11Hz -0.957142 -0.0671736
+ 1.73e+11Hz -0.95722 -0.0654605
+ 1.731e+11Hz -0.957295 -0.0637473
+ 1.732e+11Hz -0.957367 -0.0620343
+ 1.733e+11Hz -0.957436 -0.0603213
+ 1.734e+11Hz -0.957502 -0.0586083
+ 1.735e+11Hz -0.957564 -0.0568955
+ 1.736e+11Hz -0.957623 -0.0551827
+ 1.737e+11Hz -0.95768 -0.05347
+ 1.738e+11Hz -0.957733 -0.0517574
+ 1.739e+11Hz -0.957783 -0.0500449
+ 1.74e+11Hz -0.957829 -0.0483325
+ 1.741e+11Hz -0.957873 -0.0466202
+ 1.742e+11Hz -0.957913 -0.044908
+ 1.743e+11Hz -0.95795 -0.0431959
+ 1.744e+11Hz -0.957985 -0.0414839
+ 1.745e+11Hz -0.958015 -0.0397721
+ 1.746e+11Hz -0.958043 -0.0380604
+ 1.747e+11Hz -0.958068 -0.0363488
+ 1.748e+11Hz -0.958089 -0.0346374
+ 1.749e+11Hz -0.958107 -0.0329261
+ 1.75e+11Hz -0.958122 -0.031215
+ 1.751e+11Hz -0.958134 -0.0295041
+ 1.752e+11Hz -0.958143 -0.0277933
+ 1.753e+11Hz -0.958148 -0.0260827
+ 1.754e+11Hz -0.958151 -0.0243723
+ 1.755e+11Hz -0.95815 -0.0226621
+ 1.756e+11Hz -0.958146 -0.0209521
+ 1.757e+11Hz -0.958139 -0.0192423
+ 1.758e+11Hz -0.958128 -0.0175327
+ 1.759e+11Hz -0.958114 -0.0158234
+ 1.76e+11Hz -0.958098 -0.0141142
+ 1.761e+11Hz -0.958078 -0.0124054
+ 1.762e+11Hz -0.958054 -0.0106967
+ 1.763e+11Hz -0.958028 -0.00898838
+ 1.764e+11Hz -0.957998 -0.00728029
+ 1.765e+11Hz -0.957965 -0.00557247
+ 1.766e+11Hz -0.957929 -0.00386494
+ 1.767e+11Hz -0.95789 -0.0021577
+ 1.768e+11Hz -0.957848 -0.000450775
+ 1.769e+11Hz -0.957802 0.00125584
+ 1.77e+11Hz -0.957753 0.00296213
+ 1.771e+11Hz -0.957701 0.00466809
+ 1.772e+11Hz -0.957646 0.0063737
+ 1.773e+11Hz -0.957587 0.00807897
+ 1.774e+11Hz -0.957526 0.00978386
+ 1.775e+11Hz -0.957461 0.0114884
+ 1.776e+11Hz -0.957393 0.0131925
+ 1.777e+11Hz -0.957322 0.0148963
+ 1.778e+11Hz -0.957247 0.0165996
+ 1.779e+11Hz -0.957169 0.0183026
+ 1.78e+11Hz -0.957089 0.0200051
+ 1.781e+11Hz -0.957004 0.0217072
+ 1.782e+11Hz -0.956917 0.0234088
+ 1.783e+11Hz -0.956827 0.02511
+ 1.784e+11Hz -0.956733 0.0268107
+ 1.785e+11Hz -0.956636 0.028511
+ 1.786e+11Hz -0.956536 0.0302107
+ 1.787e+11Hz -0.956433 0.03191
+ 1.788e+11Hz -0.956327 0.0336088
+ 1.789e+11Hz -0.956217 0.035307
+ 1.79e+11Hz -0.956104 0.0370047
+ 1.791e+11Hz -0.955988 0.0387019
+ 1.792e+11Hz -0.955869 0.0403985
+ 1.793e+11Hz -0.955747 0.0420946
+ 1.794e+11Hz -0.955621 0.0437901
+ 1.795e+11Hz -0.955493 0.0454851
+ 1.796e+11Hz -0.955361 0.0471794
+ 1.797e+11Hz -0.955226 0.0488732
+ 1.798e+11Hz -0.955088 0.0505663
+ 1.799e+11Hz -0.954947 0.0522588
+ 1.8e+11Hz -0.954802 0.0539507
+ 1.801e+11Hz -0.954655 0.055642
+ 1.802e+11Hz -0.954504 0.0573326
+ 1.803e+11Hz -0.95435 0.0590225
+ 1.804e+11Hz -0.954193 0.0607118
+ 1.805e+11Hz -0.954033 0.0624004
+ 1.806e+11Hz -0.95387 0.0640883
+ 1.807e+11Hz -0.953704 0.0657755
+ 1.808e+11Hz -0.953534 0.067462
+ 1.809e+11Hz -0.953362 0.0691478
+ 1.81e+11Hz -0.953186 0.0708329
+ 1.811e+11Hz -0.953008 0.0725172
+ 1.812e+11Hz -0.952826 0.0742008
+ 1.813e+11Hz -0.952641 0.0758836
+ 1.814e+11Hz -0.952453 0.0775657
+ 1.815e+11Hz -0.952262 0.079247
+ 1.816e+11Hz -0.952068 0.0809275
+ 1.817e+11Hz -0.951871 0.0826072
+ 1.818e+11Hz -0.951671 0.0842862
+ 1.819e+11Hz -0.951468 0.0859643
+ 1.82e+11Hz -0.951262 0.0876416
+ 1.821e+11Hz -0.951053 0.0893181
+ 1.822e+11Hz -0.95084 0.0909938
+ 1.823e+11Hz -0.950625 0.0926686
+ 1.824e+11Hz -0.950407 0.0943425
+ 1.825e+11Hz -0.950186 0.0960157
+ 1.826e+11Hz -0.949961 0.0976879
+ 1.827e+11Hz -0.949734 0.0993593
+ 1.828e+11Hz -0.949504 0.10103
+ 1.829e+11Hz -0.949271 0.102699
+ 1.83e+11Hz -0.949035 0.104368
+ 1.831e+11Hz -0.948796 0.106036
+ 1.832e+11Hz -0.948554 0.107703
+ 1.833e+11Hz -0.948309 0.109369
+ 1.834e+11Hz -0.948061 0.111034
+ 1.835e+11Hz -0.94781 0.112698
+ 1.836e+11Hz -0.947556 0.114361
+ 1.837e+11Hz -0.947299 0.116024
+ 1.838e+11Hz -0.94704 0.117685
+ 1.839e+11Hz -0.946777 0.119345
+ 1.84e+11Hz -0.946512 0.121005
+ 1.841e+11Hz -0.946244 0.122663
+ 1.842e+11Hz -0.945972 0.124321
+ 1.843e+11Hz -0.945698 0.125977
+ 1.844e+11Hz -0.945422 0.127633
+ 1.845e+11Hz -0.945142 0.129287
+ 1.846e+11Hz -0.944859 0.130941
+ 1.847e+11Hz -0.944574 0.132594
+ 1.848e+11Hz -0.944286 0.134245
+ 1.849e+11Hz -0.943995 0.135896
+ 1.85e+11Hz -0.943701 0.137545
+ 1.851e+11Hz -0.943404 0.139194
+ 1.852e+11Hz -0.943105 0.140841
+ 1.853e+11Hz -0.942802 0.142487
+ 1.854e+11Hz -0.942497 0.144133
+ 1.855e+11Hz -0.94219 0.145777
+ 1.856e+11Hz -0.941879 0.147421
+ 1.857e+11Hz -0.941566 0.149063
+ 1.858e+11Hz -0.941249 0.150704
+ 1.859e+11Hz -0.940931 0.152344
+ 1.86e+11Hz -0.940609 0.153983
+ 1.861e+11Hz -0.940285 0.155621
+ 1.862e+11Hz -0.939958 0.157258
+ 1.863e+11Hz -0.939628 0.158894
+ 1.864e+11Hz -0.939295 0.160528
+ 1.865e+11Hz -0.93896 0.162162
+ 1.866e+11Hz -0.938622 0.163795
+ 1.867e+11Hz -0.938282 0.165426
+ 1.868e+11Hz -0.937939 0.167056
+ 1.869e+11Hz -0.937593 0.168686
+ 1.87e+11Hz -0.937244 0.170314
+ 1.871e+11Hz -0.936893 0.171941
+ 1.872e+11Hz -0.936539 0.173566
+ 1.873e+11Hz -0.936183 0.175191
+ 1.874e+11Hz -0.935823 0.176815
+ 1.875e+11Hz -0.935462 0.178437
+ 1.876e+11Hz -0.935097 0.180058
+ 1.877e+11Hz -0.93473 0.181679
+ 1.878e+11Hz -0.934361 0.183298
+ 1.879e+11Hz -0.933989 0.184915
+ 1.88e+11Hz -0.933614 0.186532
+ 1.881e+11Hz -0.933237 0.188148
+ 1.882e+11Hz -0.932857 0.189762
+ 1.883e+11Hz -0.932474 0.191375
+ 1.884e+11Hz -0.932089 0.192987
+ 1.885e+11Hz -0.931702 0.194598
+ 1.886e+11Hz -0.931312 0.196208
+ 1.887e+11Hz -0.930919 0.197816
+ 1.888e+11Hz -0.930524 0.199424
+ 1.889e+11Hz -0.930127 0.20103
+ 1.89e+11Hz -0.929727 0.202635
+ 1.891e+11Hz -0.929324 0.204238
+ 1.892e+11Hz -0.928919 0.205841
+ 1.893e+11Hz -0.928512 0.207442
+ 1.894e+11Hz -0.928102 0.209042
+ 1.895e+11Hz -0.927689 0.210641
+ 1.896e+11Hz -0.927275 0.212239
+ 1.897e+11Hz -0.926857 0.213835
+ 1.898e+11Hz -0.926438 0.21543
+ 1.899e+11Hz -0.926016 0.217024
+ 1.9e+11Hz -0.925591 0.218617
+ 1.901e+11Hz -0.925164 0.220209
+ 1.902e+11Hz -0.924735 0.221799
+ 1.903e+11Hz -0.924304 0.223388
+ 1.904e+11Hz -0.92387 0.224976
+ 1.905e+11Hz -0.923433 0.226562
+ 1.906e+11Hz -0.922995 0.228148
+ 1.907e+11Hz -0.922554 0.229732
+ 1.908e+11Hz -0.922111 0.231315
+ 1.909e+11Hz -0.921665 0.232896
+ 1.91e+11Hz -0.921217 0.234477
+ 1.911e+11Hz -0.920767 0.236056
+ 1.912e+11Hz -0.920315 0.237634
+ 1.913e+11Hz -0.91986 0.23921
+ 1.914e+11Hz -0.919403 0.240786
+ 1.915e+11Hz -0.918944 0.24236
+ 1.916e+11Hz -0.918483 0.243933
+ 1.917e+11Hz -0.918019 0.245504
+ 1.918e+11Hz -0.917554 0.247075
+ 1.919e+11Hz -0.917086 0.248644
+ 1.92e+11Hz -0.916616 0.250212
+ 1.921e+11Hz -0.916143 0.251779
+ 1.922e+11Hz -0.915669 0.253344
+ 1.923e+11Hz -0.915192 0.254908
+ 1.924e+11Hz -0.914714 0.256471
+ 1.925e+11Hz -0.914233 0.258033
+ 1.926e+11Hz -0.91375 0.259593
+ 1.927e+11Hz -0.913265 0.261153
+ 1.928e+11Hz -0.912778 0.262711
+ 1.929e+11Hz -0.912289 0.264267
+ 1.93e+11Hz -0.911798 0.265823
+ 1.931e+11Hz -0.911304 0.267377
+ 1.932e+11Hz -0.910809 0.26893
+ 1.933e+11Hz -0.910312 0.270482
+ 1.934e+11Hz -0.909813 0.272033
+ 1.935e+11Hz -0.909311 0.273583
+ 1.936e+11Hz -0.908808 0.275131
+ 1.937e+11Hz -0.908303 0.276678
+ 1.938e+11Hz -0.907796 0.278224
+ 1.939e+11Hz -0.907287 0.279769
+ 1.94e+11Hz -0.906776 0.281313
+ 1.941e+11Hz -0.906263 0.282855
+ 1.942e+11Hz -0.905748 0.284396
+ 1.943e+11Hz -0.905231 0.285937
+ 1.944e+11Hz -0.904713 0.287476
+ 1.945e+11Hz -0.904192 0.289014
+ 1.946e+11Hz -0.90367 0.29055
+ 1.947e+11Hz -0.903145 0.292086
+ 1.948e+11Hz -0.902619 0.293621
+ 1.949e+11Hz -0.902092 0.295154
+ 1.95e+11Hz -0.901562 0.296687
+ 1.951e+11Hz -0.90103 0.298218
+ 1.952e+11Hz -0.900497 0.299749
+ 1.953e+11Hz -0.899962 0.301278
+ 1.954e+11Hz -0.899425 0.302806
+ 1.955e+11Hz -0.898886 0.304333
+ 1.956e+11Hz -0.898346 0.30586
+ 1.957e+11Hz -0.897804 0.307385
+ 1.958e+11Hz -0.89726 0.308909
+ 1.959e+11Hz -0.896714 0.310432
+ 1.96e+11Hz -0.896167 0.311955
+ 1.961e+11Hz -0.895618 0.313476
+ 1.962e+11Hz -0.895067 0.314997
+ 1.963e+11Hz -0.894514 0.316516
+ 1.964e+11Hz -0.89396 0.318035
+ 1.965e+11Hz -0.893404 0.319553
+ 1.966e+11Hz -0.892846 0.32107
+ 1.967e+11Hz -0.892287 0.322586
+ 1.968e+11Hz -0.891726 0.324101
+ 1.969e+11Hz -0.891163 0.325615
+ 1.97e+11Hz -0.890599 0.327129
+ 1.971e+11Hz -0.890033 0.328642
+ 1.972e+11Hz -0.889465 0.330154
+ 1.973e+11Hz -0.888896 0.331665
+ 1.974e+11Hz -0.888325 0.333176
+ 1.975e+11Hz -0.887752 0.334686
+ 1.976e+11Hz -0.887177 0.336195
+ 1.977e+11Hz -0.886601 0.337704
+ 1.978e+11Hz -0.886024 0.339211
+ 1.979e+11Hz -0.885444 0.340719
+ 1.98e+11Hz -0.884863 0.342225
+ 1.981e+11Hz -0.884281 0.343731
+ 1.982e+11Hz -0.883696 0.345237
+ 1.983e+11Hz -0.88311 0.346742
+ 1.984e+11Hz -0.882522 0.348246
+ 1.985e+11Hz -0.881933 0.34975
+ 1.986e+11Hz -0.881342 0.351253
+ 1.987e+11Hz -0.880749 0.352756
+ 1.988e+11Hz -0.880154 0.354258
+ 1.989e+11Hz -0.879558 0.35576
+ 1.99e+11Hz -0.87896 0.357261
+ 1.991e+11Hz -0.878361 0.358762
+ 1.992e+11Hz -0.877759 0.360262
+ 1.993e+11Hz -0.877156 0.361763
+ 1.994e+11Hz -0.876551 0.363262
+ 1.995e+11Hz -0.875945 0.364762
+ 1.996e+11Hz -0.875336 0.366261
+ 1.997e+11Hz -0.874726 0.36776
+ 1.998e+11Hz -0.874114 0.369258
+ 1.999e+11Hz -0.8735 0.370756
+ 2e+11Hz -0.872885 0.372254
+ 2.001e+11Hz -0.872267 0.373752
+ 2.002e+11Hz -0.871648 0.37525
+ 2.003e+11Hz -0.871027 0.376747
+ 2.004e+11Hz -0.870404 0.378244
+ 2.005e+11Hz -0.869779 0.379741
+ 2.006e+11Hz -0.869152 0.381238
+ 2.007e+11Hz -0.868524 0.382734
+ 2.008e+11Hz -0.867893 0.384231
+ 2.009e+11Hz -0.86726 0.385727
+ 2.01e+11Hz -0.866626 0.387223
+ 2.011e+11Hz -0.865989 0.388719
+ 2.012e+11Hz -0.865351 0.390215
+ 2.013e+11Hz -0.86471 0.391711
+ 2.014e+11Hz -0.864067 0.393207
+ 2.015e+11Hz -0.863422 0.394703
+ 2.016e+11Hz -0.862775 0.396198
+ 2.017e+11Hz -0.862126 0.397694
+ 2.018e+11Hz -0.861475 0.39919
+ 2.019e+11Hz -0.860822 0.400686
+ 2.02e+11Hz -0.860166 0.402181
+ 2.021e+11Hz -0.859509 0.403677
+ 2.022e+11Hz -0.858849 0.405173
+ 2.023e+11Hz -0.858186 0.406669
+ 2.024e+11Hz -0.857522 0.408164
+ 2.025e+11Hz -0.856855 0.40966
+ 2.026e+11Hz -0.856186 0.411156
+ 2.027e+11Hz -0.855514 0.412652
+ 2.028e+11Hz -0.85484 0.414148
+ 2.029e+11Hz -0.854163 0.415644
+ 2.03e+11Hz -0.853485 0.41714
+ 2.031e+11Hz -0.852803 0.418636
+ 2.032e+11Hz -0.852119 0.420132
+ 2.033e+11Hz -0.851433 0.421628
+ 2.034e+11Hz -0.850744 0.423124
+ 2.035e+11Hz -0.850053 0.42462
+ 2.036e+11Hz -0.849358 0.426117
+ 2.037e+11Hz -0.848662 0.427613
+ 2.038e+11Hz -0.847962 0.429109
+ 2.039e+11Hz -0.84726 0.430606
+ 2.04e+11Hz -0.846555 0.432102
+ 2.041e+11Hz -0.845848 0.433598
+ 2.042e+11Hz -0.845137 0.435095
+ 2.043e+11Hz -0.844424 0.436591
+ 2.044e+11Hz -0.843708 0.438088
+ 2.045e+11Hz -0.842989 0.439584
+ 2.046e+11Hz -0.842267 0.44108
+ 2.047e+11Hz -0.841542 0.442577
+ 2.048e+11Hz -0.840815 0.444073
+ 2.049e+11Hz -0.840084 0.445569
+ 2.05e+11Hz -0.83935 0.447065
+ 2.051e+11Hz -0.838614 0.448561
+ 2.052e+11Hz -0.837874 0.450057
+ 2.053e+11Hz -0.837131 0.451553
+ 2.054e+11Hz -0.836385 0.453049
+ 2.055e+11Hz -0.835636 0.454545
+ 2.056e+11Hz -0.834884 0.45604
+ 2.057e+11Hz -0.834129 0.457535
+ 2.058e+11Hz -0.83337 0.45903
+ 2.059e+11Hz -0.832608 0.460525
+ 2.06e+11Hz -0.831843 0.462019
+ 2.061e+11Hz -0.831075 0.463514
+ 2.062e+11Hz -0.830303 0.465008
+ 2.063e+11Hz -0.829528 0.466501
+ 2.064e+11Hz -0.82875 0.467995
+ 2.065e+11Hz -0.827968 0.469488
+ 2.066e+11Hz -0.827183 0.47098
+ 2.067e+11Hz -0.826394 0.472472
+ 2.068e+11Hz -0.825602 0.473964
+ 2.069e+11Hz -0.824807 0.475456
+ 2.07e+11Hz -0.824008 0.476946
+ 2.071e+11Hz -0.823206 0.478437
+ 2.072e+11Hz -0.8224 0.479926
+ 2.073e+11Hz -0.821591 0.481416
+ 2.074e+11Hz -0.820778 0.482904
+ 2.075e+11Hz -0.819961 0.484392
+ 2.076e+11Hz -0.819141 0.48588
+ 2.077e+11Hz -0.818318 0.487366
+ 2.078e+11Hz -0.817491 0.488852
+ 2.079e+11Hz -0.81666 0.490338
+ 2.08e+11Hz -0.815825 0.491822
+ 2.081e+11Hz -0.814987 0.493306
+ 2.082e+11Hz -0.814146 0.494788
+ 2.083e+11Hz -0.8133 0.49627
+ 2.084e+11Hz -0.812451 0.497751
+ 2.085e+11Hz -0.811599 0.499232
+ 2.086e+11Hz -0.810742 0.500711
+ 2.087e+11Hz -0.809882 0.502189
+ 2.088e+11Hz -0.809019 0.503666
+ 2.089e+11Hz -0.808151 0.505142
+ 2.09e+11Hz -0.80728 0.506617
+ 2.091e+11Hz -0.806405 0.508091
+ 2.092e+11Hz -0.805527 0.509564
+ 2.093e+11Hz -0.804645 0.511035
+ 2.094e+11Hz -0.803759 0.512505
+ 2.095e+11Hz -0.802869 0.513975
+ 2.096e+11Hz -0.801976 0.515442
+ 2.097e+11Hz -0.801079 0.516909
+ 2.098e+11Hz -0.800178 0.518374
+ 2.099e+11Hz -0.799274 0.519838
+ 2.1e+11Hz -0.798366 0.5213
+ 2.101e+11Hz -0.797454 0.522761
+ 2.102e+11Hz -0.796538 0.52422
+ 2.103e+11Hz -0.795619 0.525678
+ 2.104e+11Hz -0.794696 0.527134
+ 2.105e+11Hz -0.79377 0.528589
+ 2.106e+11Hz -0.792839 0.530042
+ 2.107e+11Hz -0.791906 0.531493
+ 2.108e+11Hz -0.790968 0.532943
+ 2.109e+11Hz -0.790027 0.534391
+ 2.11e+11Hz -0.789082 0.535838
+ 2.111e+11Hz -0.788134 0.537282
+ 2.112e+11Hz -0.787182 0.538725
+ 2.113e+11Hz -0.786226 0.540166
+ 2.114e+11Hz -0.785267 0.541605
+ 2.115e+11Hz -0.784304 0.543043
+ 2.116e+11Hz -0.783338 0.544478
+ 2.117e+11Hz -0.782368 0.545912
+ 2.118e+11Hz -0.781395 0.547343
+ 2.119e+11Hz -0.780418 0.548773
+ 2.12e+11Hz -0.779438 0.5502
+ 2.121e+11Hz -0.778454 0.551626
+ 2.122e+11Hz -0.777467 0.553049
+ 2.123e+11Hz -0.776476 0.554471
+ 2.124e+11Hz -0.775482 0.55589
+ 2.125e+11Hz -0.774484 0.557307
+ 2.126e+11Hz -0.773484 0.558722
+ 2.127e+11Hz -0.772479 0.560135
+ 2.128e+11Hz -0.771472 0.561546
+ 2.129e+11Hz -0.770461 0.562954
+ 2.13e+11Hz -0.769446 0.56436
+ 2.131e+11Hz -0.768429 0.565764
+ 2.132e+11Hz -0.767408 0.567166
+ 2.133e+11Hz -0.766384 0.568565
+ 2.134e+11Hz -0.765357 0.569962
+ 2.135e+11Hz -0.764326 0.571357
+ 2.136e+11Hz -0.763293 0.57275
+ 2.137e+11Hz -0.762256 0.57414
+ 2.138e+11Hz -0.761216 0.575528
+ 2.139e+11Hz -0.760173 0.576913
+ 2.14e+11Hz -0.759127 0.578296
+ 2.141e+11Hz -0.758078 0.579677
+ 2.142e+11Hz -0.757025 0.581055
+ 2.143e+11Hz -0.75597 0.58243
+ 2.144e+11Hz -0.754912 0.583804
+ 2.145e+11Hz -0.753851 0.585175
+ 2.146e+11Hz -0.752786 0.586543
+ 2.147e+11Hz -0.751719 0.587909
+ 2.148e+11Hz -0.750649 0.589272
+ 2.149e+11Hz -0.749576 0.590633
+ 2.15e+11Hz -0.7485 0.591992
+ 2.151e+11Hz -0.747421 0.593348
+ 2.152e+11Hz -0.74634 0.594701
+ 2.153e+11Hz -0.745255 0.596052
+ 2.154e+11Hz -0.744168 0.597401
+ 2.155e+11Hz -0.743078 0.598746
+ 2.156e+11Hz -0.741985 0.60009
+ 2.157e+11Hz -0.74089 0.601431
+ 2.158e+11Hz -0.739792 0.602769
+ 2.159e+11Hz -0.738691 0.604105
+ 2.16e+11Hz -0.737587 0.605438
+ 2.161e+11Hz -0.736481 0.606769
+ 2.162e+11Hz -0.735372 0.608097
+ 2.163e+11Hz -0.734261 0.609422
+ 2.164e+11Hz -0.733147 0.610745
+ 2.165e+11Hz -0.73203 0.612066
+ 2.166e+11Hz -0.730911 0.613384
+ 2.167e+11Hz -0.729789 0.614699
+ 2.168e+11Hz -0.728665 0.616012
+ 2.169e+11Hz -0.727538 0.617322
+ 2.17e+11Hz -0.726409 0.61863
+ 2.171e+11Hz -0.725277 0.619935
+ 2.172e+11Hz -0.724142 0.621238
+ 2.173e+11Hz -0.723006 0.622538
+ 2.174e+11Hz -0.721866 0.623836
+ 2.175e+11Hz -0.720725 0.625131
+ 2.176e+11Hz -0.719581 0.626424
+ 2.177e+11Hz -0.718434 0.627714
+ 2.178e+11Hz -0.717285 0.629001
+ 2.179e+11Hz -0.716134 0.630286
+ 2.18e+11Hz -0.714981 0.631569
+ 2.181e+11Hz -0.713825 0.632848
+ 2.182e+11Hz -0.712666 0.634126
+ 2.183e+11Hz -0.711506 0.635401
+ 2.184e+11Hz -0.710343 0.636673
+ 2.185e+11Hz -0.709177 0.637943
+ 2.186e+11Hz -0.70801 0.63921
+ 2.187e+11Hz -0.70684 0.640475
+ 2.188e+11Hz -0.705667 0.641738
+ 2.189e+11Hz -0.704493 0.642998
+ 2.19e+11Hz -0.703316 0.644255
+ 2.191e+11Hz -0.702137 0.64551
+ 2.192e+11Hz -0.700955 0.646762
+ 2.193e+11Hz -0.699772 0.648012
+ 2.194e+11Hz -0.698586 0.64926
+ 2.195e+11Hz -0.697398 0.650505
+ 2.196e+11Hz -0.696207 0.651747
+ 2.197e+11Hz -0.695015 0.652987
+ 2.198e+11Hz -0.69382 0.654225
+ 2.199e+11Hz -0.692623 0.65546
+ 2.2e+11Hz -0.691423 0.656693
+ 2.201e+11Hz -0.690222 0.657923
+ 2.202e+11Hz -0.689018 0.659151
+ 2.203e+11Hz -0.687812 0.660376
+ 2.204e+11Hz -0.686604 0.661599
+ 2.205e+11Hz -0.685393 0.662819
+ 2.206e+11Hz -0.684181 0.664037
+ 2.207e+11Hz -0.682966 0.665252
+ 2.208e+11Hz -0.681749 0.666465
+ 2.209e+11Hz -0.680529 0.667675
+ 2.21e+11Hz -0.679308 0.668883
+ 2.211e+11Hz -0.678084 0.670089
+ 2.212e+11Hz -0.676858 0.671292
+ 2.213e+11Hz -0.67563 0.672492
+ 2.214e+11Hz -0.674399 0.67369
+ 2.215e+11Hz -0.673167 0.674886
+ 2.216e+11Hz -0.671932 0.676079
+ 2.217e+11Hz -0.670695 0.67727
+ 2.218e+11Hz -0.669456 0.678458
+ 2.219e+11Hz -0.668215 0.679643
+ 2.22e+11Hz -0.666971 0.680826
+ 2.221e+11Hz -0.665725 0.682007
+ 2.222e+11Hz -0.664477 0.683185
+ 2.223e+11Hz -0.663227 0.68436
+ 2.224e+11Hz -0.661975 0.685533
+ 2.225e+11Hz -0.66072 0.686703
+ 2.226e+11Hz -0.659463 0.687871
+ 2.227e+11Hz -0.658204 0.689036
+ 2.228e+11Hz -0.656943 0.690199
+ 2.229e+11Hz -0.65568 0.691359
+ 2.23e+11Hz -0.654414 0.692517
+ 2.231e+11Hz -0.653147 0.693672
+ 2.232e+11Hz -0.651877 0.694824
+ 2.233e+11Hz -0.650605 0.695974
+ 2.234e+11Hz -0.649331 0.697121
+ 2.235e+11Hz -0.648054 0.698265
+ 2.236e+11Hz -0.646776 0.699407
+ 2.237e+11Hz -0.645495 0.700546
+ 2.238e+11Hz -0.644212 0.701683
+ 2.239e+11Hz -0.642927 0.702817
+ 2.24e+11Hz -0.64164 0.703948
+ 2.241e+11Hz -0.64035 0.705076
+ 2.242e+11Hz -0.639059 0.706202
+ 2.243e+11Hz -0.637765 0.707325
+ 2.244e+11Hz -0.636469 0.708445
+ 2.245e+11Hz -0.635172 0.709563
+ 2.246e+11Hz -0.633872 0.710677
+ 2.247e+11Hz -0.63257 0.711789
+ 2.248e+11Hz -0.631265 0.712899
+ 2.249e+11Hz -0.629959 0.714005
+ 2.25e+11Hz -0.628651 0.715109
+ 2.251e+11Hz -0.62734 0.716209
+ 2.252e+11Hz -0.626028 0.717307
+ 2.253e+11Hz -0.624713 0.718402
+ 2.254e+11Hz -0.623397 0.719494
+ 2.255e+11Hz -0.622078 0.720584
+ 2.256e+11Hz -0.620758 0.72167
+ 2.257e+11Hz -0.619435 0.722754
+ 2.258e+11Hz -0.61811 0.723834
+ 2.259e+11Hz -0.616784 0.724912
+ 2.26e+11Hz -0.615455 0.725986
+ 2.261e+11Hz -0.614125 0.727058
+ 2.262e+11Hz -0.612792 0.728127
+ 2.263e+11Hz -0.611458 0.729193
+ 2.264e+11Hz -0.610122 0.730256
+ 2.265e+11Hz -0.608784 0.731315
+ 2.266e+11Hz -0.607444 0.732372
+ 2.267e+11Hz -0.606102 0.733426
+ 2.268e+11Hz -0.604758 0.734477
+ 2.269e+11Hz -0.603412 0.735524
+ 2.27e+11Hz -0.602065 0.736569
+ 2.271e+11Hz -0.600716 0.737611
+ 2.272e+11Hz -0.599365 0.738649
+ 2.273e+11Hz -0.598012 0.739684
+ 2.274e+11Hz -0.596658 0.740717
+ 2.275e+11Hz -0.595302 0.741746
+ 2.276e+11Hz -0.593944 0.742772
+ 2.277e+11Hz -0.592585 0.743795
+ 2.278e+11Hz -0.591223 0.744815
+ 2.279e+11Hz -0.589861 0.745831
+ 2.28e+11Hz -0.588496 0.746845
+ 2.281e+11Hz -0.58713 0.747855
+ 2.282e+11Hz -0.585763 0.748863
+ 2.283e+11Hz -0.584394 0.749867
+ 2.284e+11Hz -0.583023 0.750868
+ 2.285e+11Hz -0.581651 0.751865
+ 2.286e+11Hz -0.580278 0.75286
+ 2.287e+11Hz -0.578903 0.753851
+ 2.288e+11Hz -0.577526 0.75484
+ 2.289e+11Hz -0.576149 0.755825
+ 2.29e+11Hz -0.57477 0.756807
+ 2.291e+11Hz -0.573389 0.757785
+ 2.292e+11Hz -0.572007 0.758761
+ 2.293e+11Hz -0.570624 0.759733
+ 2.294e+11Hz -0.56924 0.760702
+ 2.295e+11Hz -0.567854 0.761668
+ 2.296e+11Hz -0.566467 0.762631
+ 2.297e+11Hz -0.565079 0.763591
+ 2.298e+11Hz -0.563689 0.764547
+ 2.299e+11Hz -0.562299 0.7655
+ 2.3e+11Hz -0.560907 0.76645
+ 2.301e+11Hz -0.559515 0.767397
+ 2.302e+11Hz -0.558121 0.768341
+ 2.303e+11Hz -0.556726 0.769282
+ 2.304e+11Hz -0.55533 0.770219
+ 2.305e+11Hz -0.553933 0.771154
+ 2.306e+11Hz -0.552535 0.772085
+ 2.307e+11Hz -0.551136 0.773013
+ 2.308e+11Hz -0.549736 0.773938
+ 2.309e+11Hz -0.548335 0.77486
+ 2.31e+11Hz -0.546934 0.775779
+ 2.311e+11Hz -0.545531 0.776695
+ 2.312e+11Hz -0.544128 0.777608
+ 2.313e+11Hz -0.542723 0.778517
+ 2.314e+11Hz -0.541318 0.779424
+ 2.315e+11Hz -0.539912 0.780328
+ 2.316e+11Hz -0.538505 0.781228
+ 2.317e+11Hz -0.537098 0.782126
+ 2.318e+11Hz -0.53569 0.78302
+ 2.319e+11Hz -0.534281 0.783912
+ 2.32e+11Hz -0.532871 0.784801
+ 2.321e+11Hz -0.531461 0.785686
+ 2.322e+11Hz -0.53005 0.786569
+ 2.323e+11Hz -0.528639 0.787449
+ 2.324e+11Hz -0.527226 0.788326
+ 2.325e+11Hz -0.525814 0.789201
+ 2.326e+11Hz -0.5244 0.790072
+ 2.327e+11Hz -0.522986 0.79094
+ 2.328e+11Hz -0.521572 0.791806
+ 2.329e+11Hz -0.520157 0.792669
+ 2.33e+11Hz -0.518741 0.793529
+ 2.331e+11Hz -0.517325 0.794386
+ 2.332e+11Hz -0.515908 0.795241
+ 2.333e+11Hz -0.514491 0.796093
+ 2.334e+11Hz -0.513073 0.796942
+ 2.335e+11Hz -0.511655 0.797789
+ 2.336e+11Hz -0.510237 0.798633
+ 2.337e+11Hz -0.508818 0.799474
+ 2.338e+11Hz -0.507398 0.800313
+ 2.339e+11Hz -0.505978 0.801149
+ 2.34e+11Hz -0.504558 0.801982
+ 2.341e+11Hz -0.503137 0.802813
+ 2.342e+11Hz -0.501716 0.803642
+ 2.343e+11Hz -0.500295 0.804468
+ 2.344e+11Hz -0.498873 0.805291
+ 2.345e+11Hz -0.497451 0.806112
+ 2.346e+11Hz -0.496028 0.806931
+ 2.347e+11Hz -0.494605 0.807747
+ 2.348e+11Hz -0.493181 0.808561
+ 2.349e+11Hz -0.491757 0.809372
+ 2.35e+11Hz -0.490333 0.810181
+ 2.351e+11Hz -0.488909 0.810988
+ 2.352e+11Hz -0.487484 0.811792
+ 2.353e+11Hz -0.486058 0.812595
+ 2.354e+11Hz -0.484633 0.813395
+ 2.355e+11Hz -0.483207 0.814192
+ 2.356e+11Hz -0.48178 0.814988
+ 2.357e+11Hz -0.480353 0.815781
+ 2.358e+11Hz -0.478926 0.816572
+ 2.359e+11Hz -0.477499 0.817361
+ 2.36e+11Hz -0.476071 0.818148
+ 2.361e+11Hz -0.474642 0.818933
+ 2.362e+11Hz -0.473213 0.819716
+ 2.363e+11Hz -0.471784 0.820496
+ 2.364e+11Hz -0.470355 0.821275
+ 2.365e+11Hz -0.468925 0.822051
+ 2.366e+11Hz -0.467494 0.822826
+ 2.367e+11Hz -0.466063 0.823598
+ 2.368e+11Hz -0.464632 0.824369
+ 2.369e+11Hz -0.4632 0.825138
+ 2.37e+11Hz -0.461768 0.825904
+ 2.371e+11Hz -0.460335 0.826669
+ 2.372e+11Hz -0.458902 0.827432
+ 2.373e+11Hz -0.457469 0.828193
+ 2.374e+11Hz -0.456035 0.828952
+ 2.375e+11Hz -0.4546 0.829709
+ 2.376e+11Hz -0.453165 0.830465
+ 2.377e+11Hz -0.451729 0.831218
+ 2.378e+11Hz -0.450293 0.83197
+ 2.379e+11Hz -0.448856 0.83272
+ 2.38e+11Hz -0.447419 0.833468
+ 2.381e+11Hz -0.445981 0.834215
+ 2.382e+11Hz -0.444542 0.83496
+ 2.383e+11Hz -0.443103 0.835703
+ 2.384e+11Hz -0.441663 0.836444
+ 2.385e+11Hz -0.440223 0.837183
+ 2.386e+11Hz -0.438782 0.837921
+ 2.387e+11Hz -0.43734 0.838657
+ 2.388e+11Hz -0.435897 0.839392
+ 2.389e+11Hz -0.434454 0.840125
+ 2.39e+11Hz -0.43301 0.840856
+ 2.391e+11Hz -0.431566 0.841585
+ 2.392e+11Hz -0.430121 0.842313
+ 2.393e+11Hz -0.428674 0.843039
+ 2.394e+11Hz -0.427228 0.843764
+ 2.395e+11Hz -0.42578 0.844487
+ 2.396e+11Hz -0.424331 0.845208
+ 2.397e+11Hz -0.422882 0.845928
+ 2.398e+11Hz -0.421432 0.846646
+ 2.399e+11Hz -0.419981 0.847362
+ 2.4e+11Hz -0.418529 0.848077
+ 2.401e+11Hz -0.417076 0.84879
+ 2.402e+11Hz -0.415623 0.849502
+ 2.403e+11Hz -0.414168 0.850212
+ 2.404e+11Hz -0.412713 0.85092
+ 2.405e+11Hz -0.411256 0.851627
+ 2.406e+11Hz -0.409799 0.852333
+ 2.407e+11Hz -0.40834 0.853036
+ 2.408e+11Hz -0.406881 0.853738
+ 2.409e+11Hz -0.40542 0.854439
+ 2.41e+11Hz -0.403959 0.855138
+ 2.411e+11Hz -0.402496 0.855835
+ 2.412e+11Hz -0.401032 0.856531
+ 2.413e+11Hz -0.399568 0.857225
+ 2.414e+11Hz -0.398102 0.857917
+ 2.415e+11Hz -0.396635 0.858608
+ 2.416e+11Hz -0.395167 0.859298
+ 2.417e+11Hz -0.393698 0.859985
+ 2.418e+11Hz -0.392228 0.860671
+ 2.419e+11Hz -0.390756 0.861356
+ 2.42e+11Hz -0.389283 0.862039
+ 2.421e+11Hz -0.387809 0.86272
+ 2.422e+11Hz -0.386334 0.8634
+ 2.423e+11Hz -0.384858 0.864078
+ 2.424e+11Hz -0.38338 0.864754
+ 2.425e+11Hz -0.381902 0.865429
+ 2.426e+11Hz -0.380422 0.866102
+ 2.427e+11Hz -0.37894 0.866773
+ 2.428e+11Hz -0.377458 0.867443
+ 2.429e+11Hz -0.375974 0.868111
+ 2.43e+11Hz -0.374488 0.868778
+ 2.431e+11Hz -0.373002 0.869442
+ 2.432e+11Hz -0.371514 0.870105
+ 2.433e+11Hz -0.370025 0.870767
+ 2.434e+11Hz -0.368534 0.871426
+ 2.435e+11Hz -0.367042 0.872084
+ 2.436e+11Hz -0.365549 0.87274
+ 2.437e+11Hz -0.364054 0.873395
+ 2.438e+11Hz -0.362558 0.874048
+ 2.439e+11Hz -0.36106 0.874699
+ 2.44e+11Hz -0.359561 0.875348
+ 2.441e+11Hz -0.358061 0.875995
+ 2.442e+11Hz -0.356559 0.876641
+ 2.443e+11Hz -0.355055 0.877285
+ 2.444e+11Hz -0.353551 0.877927
+ 2.445e+11Hz -0.352044 0.878568
+ 2.446e+11Hz -0.350537 0.879206
+ 2.447e+11Hz -0.349027 0.879843
+ 2.448e+11Hz -0.347517 0.880478
+ 2.449e+11Hz -0.346004 0.881111
+ 2.45e+11Hz -0.344491 0.881742
+ 2.451e+11Hz -0.342975 0.882371
+ 2.452e+11Hz -0.341459 0.882999
+ 2.453e+11Hz -0.33994 0.883625
+ 2.454e+11Hz -0.338421 0.884248
+ 2.455e+11Hz -0.336899 0.88487
+ 2.456e+11Hz -0.335376 0.88549
+ 2.457e+11Hz -0.333852 0.886108
+ 2.458e+11Hz -0.332326 0.886724
+ 2.459e+11Hz -0.330798 0.887338
+ 2.46e+11Hz -0.329269 0.887951
+ 2.461e+11Hz -0.327738 0.888561
+ 2.462e+11Hz -0.326206 0.889169
+ 2.463e+11Hz -0.324672 0.889776
+ 2.464e+11Hz -0.323136 0.89038
+ 2.465e+11Hz -0.321599 0.890982
+ 2.466e+11Hz -0.32006 0.891583
+ 2.467e+11Hz -0.318519 0.892181
+ 2.468e+11Hz -0.316977 0.892777
+ 2.469e+11Hz -0.315434 0.893372
+ 2.47e+11Hz -0.313888 0.893964
+ 2.471e+11Hz -0.312341 0.894554
+ 2.472e+11Hz -0.310793 0.895142
+ 2.473e+11Hz -0.309242 0.895728
+ 2.474e+11Hz -0.30769 0.896312
+ 2.475e+11Hz -0.306137 0.896894
+ 2.476e+11Hz -0.304581 0.897474
+ 2.477e+11Hz -0.303024 0.898052
+ 2.478e+11Hz -0.301466 0.898627
+ 2.479e+11Hz -0.299905 0.8992
+ 2.48e+11Hz -0.298343 0.899772
+ 2.481e+11Hz -0.29678 0.900341
+ 2.482e+11Hz -0.295214 0.900907
+ 2.483e+11Hz -0.293647 0.901472
+ 2.484e+11Hz -0.292078 0.902035
+ 2.485e+11Hz -0.290507 0.902595
+ 2.486e+11Hz -0.288935 0.903153
+ 2.487e+11Hz -0.287361 0.903709
+ 2.488e+11Hz -0.285785 0.904262
+ 2.489e+11Hz -0.284208 0.904814
+ 2.49e+11Hz -0.282629 0.905363
+ 2.491e+11Hz -0.281048 0.90591
+ 2.492e+11Hz -0.279465 0.906454
+ 2.493e+11Hz -0.27788 0.906996
+ 2.494e+11Hz -0.276294 0.907536
+ 2.495e+11Hz -0.274706 0.908074
+ 2.496e+11Hz -0.273116 0.908609
+ 2.497e+11Hz -0.271525 0.909142
+ 2.498e+11Hz -0.269931 0.909672
+ 2.499e+11Hz -0.268336 0.9102
+ 2.5e+11Hz -0.266739 0.910726
+ 2.501e+11Hz -0.26514 0.911249
+ 2.502e+11Hz -0.26354 0.91177
+ 2.503e+11Hz -0.261937 0.912289
+ 2.504e+11Hz -0.260333 0.912805
+ 2.505e+11Hz -0.258727 0.913318
+ 2.506e+11Hz -0.257119 0.913829
+ 2.507e+11Hz -0.25551 0.914338
+ 2.508e+11Hz -0.253898 0.914844
+ 2.509e+11Hz -0.252285 0.915347
+ 2.51e+11Hz -0.25067 0.915848
+ 2.511e+11Hz -0.249053 0.916346
+ 2.512e+11Hz -0.247434 0.916842
+ 2.513e+11Hz -0.245814 0.917335
+ 2.514e+11Hz -0.244191 0.917826
+ 2.515e+11Hz -0.242567 0.918314
+ 2.516e+11Hz -0.240941 0.918799
+ 2.517e+11Hz -0.239313 0.919282
+ 2.518e+11Hz -0.237683 0.919762
+ 2.519e+11Hz -0.236051 0.920239
+ 2.52e+11Hz -0.234418 0.920714
+ 2.521e+11Hz -0.232782 0.921185
+ 2.522e+11Hz -0.231145 0.921654
+ 2.523e+11Hz -0.229506 0.922121
+ 2.524e+11Hz -0.227865 0.922584
+ 2.525e+11Hz -0.226222 0.923045
+ 2.526e+11Hz -0.224577 0.923502
+ 2.527e+11Hz -0.22293 0.923957
+ 2.528e+11Hz -0.221282 0.924409
+ 2.529e+11Hz -0.219631 0.924859
+ 2.53e+11Hz -0.217979 0.925305
+ 2.531e+11Hz -0.216325 0.925748
+ 2.532e+11Hz -0.214669 0.926188
+ 2.533e+11Hz -0.213011 0.926626
+ 2.534e+11Hz -0.211351 0.92706
+ 2.535e+11Hz -0.20969 0.927491
+ 2.536e+11Hz -0.208026 0.92792
+ 2.537e+11Hz -0.206361 0.928345
+ 2.538e+11Hz -0.204694 0.928767
+ 2.539e+11Hz -0.203025 0.929186
+ 2.54e+11Hz -0.201354 0.929602
+ 2.541e+11Hz -0.199682 0.930014
+ 2.542e+11Hz -0.198007 0.930424
+ 2.543e+11Hz -0.196331 0.93083
+ 2.544e+11Hz -0.194653 0.931233
+ 2.545e+11Hz -0.192973 0.931633
+ 2.546e+11Hz -0.191291 0.932029
+ 2.547e+11Hz -0.189608 0.932422
+ 2.548e+11Hz -0.187923 0.932812
+ 2.549e+11Hz -0.186236 0.933199
+ 2.55e+11Hz -0.184547 0.933582
+ 2.551e+11Hz -0.182856 0.933961
+ 2.552e+11Hz -0.181164 0.934338
+ 2.553e+11Hz -0.17947 0.93471
+ 2.554e+11Hz -0.177774 0.93508
+ 2.555e+11Hz -0.176077 0.935446
+ 2.556e+11Hz -0.174378 0.935808
+ 2.557e+11Hz -0.172677 0.936167
+ 2.558e+11Hz -0.170974 0.936522
+ 2.559e+11Hz -0.16927 0.936873
+ 2.56e+11Hz -0.167564 0.937221
+ 2.561e+11Hz -0.165857 0.937565
+ 2.562e+11Hz -0.164148 0.937906
+ 2.563e+11Hz -0.162437 0.938243
+ 2.564e+11Hz -0.160725 0.938576
+ 2.565e+11Hz -0.159011 0.938906
+ 2.566e+11Hz -0.157296 0.939232
+ 2.567e+11Hz -0.155579 0.939554
+ 2.568e+11Hz -0.153861 0.939872
+ 2.569e+11Hz -0.152141 0.940186
+ 2.57e+11Hz -0.15042 0.940497
+ 2.571e+11Hz -0.148698 0.940803
+ 2.572e+11Hz -0.146974 0.941106
+ 2.573e+11Hz -0.145248 0.941405
+ 2.574e+11Hz -0.143521 0.9417
+ 2.575e+11Hz -0.141793 0.941991
+ 2.576e+11Hz -0.140064 0.942278
+ 2.577e+11Hz -0.138333 0.942561
+ 2.578e+11Hz -0.136601 0.94284
+ 2.579e+11Hz -0.134867 0.943115
+ 2.58e+11Hz -0.133133 0.943386
+ 2.581e+11Hz -0.131397 0.943652
+ 2.582e+11Hz -0.12966 0.943915
+ 2.583e+11Hz -0.127922 0.944174
+ 2.584e+11Hz -0.126183 0.944429
+ 2.585e+11Hz -0.124442 0.944679
+ 2.586e+11Hz -0.122701 0.944926
+ 2.587e+11Hz -0.120959 0.945168
+ 2.588e+11Hz -0.119215 0.945406
+ 2.589e+11Hz -0.117471 0.94564
+ 2.59e+11Hz -0.115725 0.945869
+ 2.591e+11Hz -0.113979 0.946095
+ 2.592e+11Hz -0.112232 0.946316
+ 2.593e+11Hz -0.110484 0.946533
+ 2.594e+11Hz -0.108735 0.946746
+ 2.595e+11Hz -0.106985 0.946955
+ 2.596e+11Hz -0.105235 0.947159
+ 2.597e+11Hz -0.103484 0.947359
+ 2.598e+11Hz -0.101732 0.947555
+ 2.599e+11Hz -0.0999791 0.947746
+ 2.6e+11Hz -0.0982258 0.947934
+ 2.601e+11Hz -0.096472 0.948117
+ 2.602e+11Hz -0.0947175 0.948295
+ 2.603e+11Hz -0.0929624 0.94847
+ 2.604e+11Hz -0.0912069 0.94864
+ 2.605e+11Hz -0.0894508 0.948806
+ 2.606e+11Hz -0.0876943 0.948967
+ 2.607e+11Hz -0.0859373 0.949124
+ 2.608e+11Hz -0.0841799 0.949277
+ 2.609e+11Hz -0.0824222 0.949426
+ 2.61e+11Hz -0.0806641 0.94957
+ 2.611e+11Hz -0.0789057 0.94971
+ 2.612e+11Hz -0.0771471 0.949845
+ 2.613e+11Hz -0.0753881 0.949977
+ 2.614e+11Hz -0.073629 0.950104
+ 2.615e+11Hz -0.0718697 0.950226
+ 2.616e+11Hz -0.0701102 0.950345
+ 2.617e+11Hz -0.0683506 0.950459
+ 2.618e+11Hz -0.0665909 0.950569
+ 2.619e+11Hz -0.0648311 0.950674
+ 2.62e+11Hz -0.0630713 0.950775
+ 2.621e+11Hz -0.0613115 0.950872
+ 2.622e+11Hz -0.0595517 0.950965
+ 2.623e+11Hz -0.0577919 0.951054
+ 2.624e+11Hz -0.0560322 0.951138
+ 2.625e+11Hz -0.0542727 0.951218
+ 2.626e+11Hz -0.0525132 0.951294
+ 2.627e+11Hz -0.0507539 0.951365
+ 2.628e+11Hz -0.0489948 0.951432
+ 2.629e+11Hz -0.047236 0.951496
+ 2.63e+11Hz -0.0454773 0.951554
+ 2.631e+11Hz -0.0437189 0.951609
+ 2.632e+11Hz -0.0419608 0.95166
+ 2.633e+11Hz -0.0402031 0.951706
+ 2.634e+11Hz -0.0384456 0.951749
+ 2.635e+11Hz -0.0366886 0.951787
+ 2.636e+11Hz -0.0349319 0.951821
+ 2.637e+11Hz -0.0331756 0.951851
+ 2.638e+11Hz -0.0314197 0.951877
+ 2.639e+11Hz -0.0296643 0.951899
+ 2.64e+11Hz -0.0279094 0.951916
+ 2.641e+11Hz -0.026155 0.95193
+ 2.642e+11Hz -0.0244011 0.95194
+ 2.643e+11Hz -0.0226477 0.951945
+ 2.644e+11Hz -0.0208949 0.951947
+ 2.645e+11Hz -0.0191427 0.951945
+ 2.646e+11Hz -0.017391 0.951939
+ 2.647e+11Hz -0.01564 0.951928
+ 2.648e+11Hz -0.0138896 0.951914
+ 2.649e+11Hz -0.0121398 0.951896
+ 2.65e+11Hz -0.0103907 0.951874
+ 2.651e+11Hz -0.0086423 0.951849
+ 2.652e+11Hz -0.00689458 0.951819
+ 2.653e+11Hz -0.00514756 0.951785
+ 2.654e+11Hz -0.00340127 0.951748
+ 2.655e+11Hz -0.00165571 0.951707
+ 2.656e+11Hz 8.90999e-05 0.951662
+ 2.657e+11Hz 0.00183314 0.951613
+ 2.658e+11Hz 0.00357641 0.951561
+ 2.659e+11Hz 0.00531889 0.951504
+ 2.66e+11Hz 0.00706058 0.951444
+ 2.661e+11Hz 0.00880145 0.951381
+ 2.662e+11Hz 0.0105415 0.951313
+ 2.663e+11Hz 0.0122807 0.951242
+ 2.664e+11Hz 0.0140191 0.951168
+ 2.665e+11Hz 0.0157566 0.951089
+ 2.666e+11Hz 0.0174933 0.951007
+ 2.667e+11Hz 0.0192291 0.950922
+ 2.668e+11Hz 0.020964 0.950832
+ 2.669e+11Hz 0.0226981 0.95074
+ 2.67e+11Hz 0.0244312 0.950643
+ 2.671e+11Hz 0.0261635 0.950543
+ 2.672e+11Hz 0.0278948 0.95044
+ 2.673e+11Hz 0.0296253 0.950333
+ 2.674e+11Hz 0.0313548 0.950222
+ 2.675e+11Hz 0.0330834 0.950108
+ 2.676e+11Hz 0.0348111 0.949991
+ 2.677e+11Hz 0.0365378 0.94987
+ 2.678e+11Hz 0.0382636 0.949746
+ 2.679e+11Hz 0.0399885 0.949618
+ 2.68e+11Hz 0.0417124 0.949486
+ 2.681e+11Hz 0.0434354 0.949352
+ 2.682e+11Hz 0.0451574 0.949214
+ 2.683e+11Hz 0.0468784 0.949072
+ 2.684e+11Hz 0.0485985 0.948927
+ 2.685e+11Hz 0.0503176 0.948779
+ 2.686e+11Hz 0.0520358 0.948627
+ 2.687e+11Hz 0.053753 0.948472
+ 2.688e+11Hz 0.0554692 0.948314
+ 2.689e+11Hz 0.0571844 0.948152
+ 2.69e+11Hz 0.0588986 0.947987
+ 2.691e+11Hz 0.0606118 0.947819
+ 2.692e+11Hz 0.0623241 0.947647
+ 2.693e+11Hz 0.0640353 0.947472
+ 2.694e+11Hz 0.0657456 0.947294
+ 2.695e+11Hz 0.0674549 0.947112
+ 2.696e+11Hz 0.0691631 0.946928
+ 2.697e+11Hz 0.0708703 0.94674
+ 2.698e+11Hz 0.0725766 0.946548
+ 2.699e+11Hz 0.0742818 0.946354
+ 2.7e+11Hz 0.075986 0.946156
+ 2.701e+11Hz 0.0776892 0.945955
+ 2.702e+11Hz 0.0793913 0.94575
+ 2.703e+11Hz 0.0810924 0.945543
+ 2.704e+11Hz 0.0827925 0.945332
+ 2.705e+11Hz 0.0844915 0.945118
+ 2.706e+11Hz 0.0861895 0.944901
+ 2.707e+11Hz 0.0878865 0.944681
+ 2.708e+11Hz 0.0895824 0.944457
+ 2.709e+11Hz 0.0912772 0.94423
+ 2.71e+11Hz 0.092971 0.944
+ 2.711e+11Hz 0.0946637 0.943767
+ 2.712e+11Hz 0.0963553 0.943531
+ 2.713e+11Hz 0.0980458 0.943291
+ 2.714e+11Hz 0.0997353 0.943048
+ 2.715e+11Hz 0.101424 0.942802
+ 2.716e+11Hz 0.103111 0.942553
+ 2.717e+11Hz 0.104797 0.942301
+ 2.718e+11Hz 0.106482 0.942045
+ 2.719e+11Hz 0.108166 0.941787
+ 2.72e+11Hz 0.109849 0.941525
+ 2.721e+11Hz 0.11153 0.94126
+ 2.722e+11Hz 0.113211 0.940992
+ 2.723e+11Hz 0.11489 0.940721
+ 2.724e+11Hz 0.116568 0.940447
+ 2.725e+11Hz 0.118245 0.940169
+ 2.726e+11Hz 0.119921 0.939889
+ 2.727e+11Hz 0.121595 0.939605
+ 2.728e+11Hz 0.123269 0.939318
+ 2.729e+11Hz 0.124941 0.939028
+ 2.73e+11Hz 0.126612 0.938735
+ 2.731e+11Hz 0.128282 0.938439
+ 2.732e+11Hz 0.12995 0.93814
+ 2.733e+11Hz 0.131617 0.937837
+ 2.734e+11Hz 0.133283 0.937532
+ 2.735e+11Hz 0.134948 0.937223
+ 2.736e+11Hz 0.136611 0.936912
+ 2.737e+11Hz 0.138273 0.936597
+ 2.738e+11Hz 0.139934 0.936279
+ 2.739e+11Hz 0.141593 0.935959
+ 2.74e+11Hz 0.143251 0.935635
+ 2.741e+11Hz 0.144907 0.935308
+ 2.742e+11Hz 0.146563 0.934978
+ 2.743e+11Hz 0.148216 0.934645
+ 2.744e+11Hz 0.149869 0.934309
+ 2.745e+11Hz 0.15152 0.933971
+ 2.746e+11Hz 0.15317 0.933629
+ 2.747e+11Hz 0.154818 0.933284
+ 2.748e+11Hz 0.156464 0.932936
+ 2.749e+11Hz 0.15811 0.932585
+ 2.75e+11Hz 0.159753 0.932232
+ 2.751e+11Hz 0.161396 0.931875
+ 2.752e+11Hz 0.163036 0.931515
+ 2.753e+11Hz 0.164675 0.931153
+ 2.754e+11Hz 0.166313 0.930788
+ 2.755e+11Hz 0.167949 0.930419
+ 2.756e+11Hz 0.169584 0.930048
+ 2.757e+11Hz 0.171217 0.929675
+ 2.758e+11Hz 0.172848 0.929298
+ 2.759e+11Hz 0.174478 0.928918
+ 2.76e+11Hz 0.176106 0.928536
+ 2.761e+11Hz 0.177733 0.928151
+ 2.762e+11Hz 0.179358 0.927763
+ 2.763e+11Hz 0.180981 0.927372
+ 2.764e+11Hz 0.182602 0.926979
+ 2.765e+11Hz 0.184222 0.926583
+ 2.766e+11Hz 0.18584 0.926184
+ 2.767e+11Hz 0.187457 0.925783
+ 2.768e+11Hz 0.189072 0.925379
+ 2.769e+11Hz 0.190685 0.924972
+ 2.77e+11Hz 0.192296 0.924563
+ 2.771e+11Hz 0.193906 0.924151
+ 2.772e+11Hz 0.195514 0.923737
+ 2.773e+11Hz 0.19712 0.92332
+ 2.774e+11Hz 0.198724 0.922901
+ 2.775e+11Hz 0.200327 0.922479
+ 2.776e+11Hz 0.201928 0.922055
+ 2.777e+11Hz 0.203527 0.921628
+ 2.778e+11Hz 0.205124 0.921199
+ 2.779e+11Hz 0.20672 0.920767
+ 2.78e+11Hz 0.208314 0.920333
+ 2.781e+11Hz 0.209906 0.919897
+ 2.782e+11Hz 0.211496 0.919459
+ 2.783e+11Hz 0.213084 0.919018
+ 2.784e+11Hz 0.214671 0.918575
+ 2.785e+11Hz 0.216256 0.918129
+ 2.786e+11Hz 0.217839 0.917682
+ 2.787e+11Hz 0.21942 0.917232
+ 2.788e+11Hz 0.220999 0.91678
+ 2.789e+11Hz 0.222577 0.916327
+ 2.79e+11Hz 0.224152 0.915871
+ 2.791e+11Hz 0.225726 0.915412
+ 2.792e+11Hz 0.227299 0.914952
+ 2.793e+11Hz 0.228869 0.91449
+ 2.794e+11Hz 0.230438 0.914026
+ 2.795e+11Hz 0.232005 0.91356
+ 2.796e+11Hz 0.23357 0.913092
+ 2.797e+11Hz 0.235133 0.912622
+ 2.798e+11Hz 0.236695 0.91215
+ 2.799e+11Hz 0.238255 0.911677
+ 2.8e+11Hz 0.239813 0.911201
+ 2.801e+11Hz 0.24137 0.910724
+ 2.802e+11Hz 0.242925 0.910245
+ 2.803e+11Hz 0.244478 0.909764
+ 2.804e+11Hz 0.246029 0.909282
+ 2.805e+11Hz 0.247579 0.908798
+ 2.806e+11Hz 0.249127 0.908312
+ 2.807e+11Hz 0.250674 0.907824
+ 2.808e+11Hz 0.252219 0.907335
+ 2.809e+11Hz 0.253762 0.906844
+ 2.81e+11Hz 0.255304 0.906352
+ 2.811e+11Hz 0.256844 0.905858
+ 2.812e+11Hz 0.258383 0.905363
+ 2.813e+11Hz 0.25992 0.904866
+ 2.814e+11Hz 0.261456 0.904368
+ 2.815e+11Hz 0.26299 0.903868
+ 2.816e+11Hz 0.264523 0.903367
+ 2.817e+11Hz 0.266055 0.902864
+ 2.818e+11Hz 0.267585 0.90236
+ 2.819e+11Hz 0.269114 0.901855
+ 2.82e+11Hz 0.270641 0.901348
+ 2.821e+11Hz 0.272167 0.90084
+ 2.822e+11Hz 0.273692 0.900331
+ 2.823e+11Hz 0.275215 0.89982
+ 2.824e+11Hz 0.276737 0.899308
+ 2.825e+11Hz 0.278259 0.898795
+ 2.826e+11Hz 0.279778 0.89828
+ 2.827e+11Hz 0.281297 0.897764
+ 2.828e+11Hz 0.282815 0.897247
+ 2.829e+11Hz 0.284331 0.896729
+ 2.83e+11Hz 0.285847 0.896209
+ 2.831e+11Hz 0.287361 0.895688
+ 2.832e+11Hz 0.288875 0.895166
+ 2.833e+11Hz 0.290387 0.894643
+ 2.834e+11Hz 0.291899 0.894118
+ 2.835e+11Hz 0.29341 0.893593
+ 2.836e+11Hz 0.294919 0.893066
+ 2.837e+11Hz 0.296428 0.892538
+ 2.838e+11Hz 0.297937 0.892009
+ 2.839e+11Hz 0.299444 0.891478
+ 2.84e+11Hz 0.300951 0.890947
+ 2.841e+11Hz 0.302457 0.890414
+ 2.842e+11Hz 0.303962 0.88988
+ 2.843e+11Hz 0.305467 0.889345
+ 2.844e+11Hz 0.306971 0.888808
+ 2.845e+11Hz 0.308474 0.888271
+ 2.846e+11Hz 0.309977 0.887732
+ 2.847e+11Hz 0.311479 0.887192
+ 2.848e+11Hz 0.312981 0.886651
+ 2.849e+11Hz 0.314483 0.886108
+ 2.85e+11Hz 0.315984 0.885564
+ 2.851e+11Hz 0.317485 0.885019
+ 2.852e+11Hz 0.318985 0.884473
+ 2.853e+11Hz 0.320485 0.883926
+ 2.854e+11Hz 0.321985 0.883377
+ 2.855e+11Hz 0.323484 0.882827
+ 2.856e+11Hz 0.324984 0.882275
+ 2.857e+11Hz 0.326483 0.881722
+ 2.858e+11Hz 0.327982 0.881168
+ 2.859e+11Hz 0.32948 0.880613
+ 2.86e+11Hz 0.330979 0.880056
+ 2.861e+11Hz 0.332478 0.879497
+ 2.862e+11Hz 0.333976 0.878937
+ 2.863e+11Hz 0.335475 0.878376
+ 2.864e+11Hz 0.336973 0.877813
+ 2.865e+11Hz 0.338471 0.877249
+ 2.866e+11Hz 0.33997 0.876683
+ 2.867e+11Hz 0.341468 0.876115
+ 2.868e+11Hz 0.342967 0.875546
+ 2.869e+11Hz 0.344466 0.874976
+ 2.87e+11Hz 0.345965 0.874403
+ 2.871e+11Hz 0.347464 0.873829
+ 2.872e+11Hz 0.348963 0.873254
+ 2.873e+11Hz 0.350462 0.872676
+ 2.874e+11Hz 0.351962 0.872097
+ 2.875e+11Hz 0.353462 0.871516
+ 2.876e+11Hz 0.354962 0.870933
+ 2.877e+11Hz 0.356462 0.870348
+ 2.878e+11Hz 0.357962 0.869762
+ 2.879e+11Hz 0.359463 0.869173
+ 2.88e+11Hz 0.360964 0.868583
+ 2.881e+11Hz 0.362466 0.86799
+ 2.882e+11Hz 0.363967 0.867396
+ 2.883e+11Hz 0.365469 0.866799
+ 2.884e+11Hz 0.366972 0.8662
+ 2.885e+11Hz 0.368474 0.865599
+ 2.886e+11Hz 0.369977 0.864996
+ 2.887e+11Hz 0.37148 0.864391
+ 2.888e+11Hz 0.372984 0.863784
+ 2.889e+11Hz 0.374488 0.863174
+ 2.89e+11Hz 0.375992 0.862562
+ 2.891e+11Hz 0.377497 0.861947
+ 2.892e+11Hz 0.379002 0.861331
+ 2.893e+11Hz 0.380507 0.860711
+ 2.894e+11Hz 0.382013 0.86009
+ 2.895e+11Hz 0.383519 0.859466
+ 2.896e+11Hz 0.385025 0.858839
+ 2.897e+11Hz 0.386532 0.85821
+ 2.898e+11Hz 0.388039 0.857578
+ 2.899e+11Hz 0.389546 0.856943
+ 2.9e+11Hz 0.391053 0.856306
+ 2.901e+11Hz 0.392561 0.855666
+ 2.902e+11Hz 0.394069 0.855023
+ 2.903e+11Hz 0.395577 0.854378
+ 2.904e+11Hz 0.397086 0.85373
+ 2.905e+11Hz 0.398595 0.853079
+ 2.906e+11Hz 0.400104 0.852425
+ 2.907e+11Hz 0.401613 0.851768
+ 2.908e+11Hz 0.403122 0.851108
+ 2.909e+11Hz 0.404632 0.850445
+ 2.91e+11Hz 0.406142 0.849779
+ 2.911e+11Hz 0.407651 0.849111
+ 2.912e+11Hz 0.409161 0.848439
+ 2.913e+11Hz 0.410671 0.847764
+ 2.914e+11Hz 0.412181 0.847086
+ 2.915e+11Hz 0.413692 0.846405
+ 2.916e+11Hz 0.415202 0.84572
+ 2.917e+11Hz 0.416712 0.845033
+ 2.918e+11Hz 0.418222 0.844342
+ 2.919e+11Hz 0.419732 0.843648
+ 2.92e+11Hz 0.421242 0.842951
+ 2.921e+11Hz 0.422751 0.84225
+ 2.922e+11Hz 0.424261 0.841546
+ 2.923e+11Hz 0.425771 0.840839
+ 2.924e+11Hz 0.42728 0.840128
+ 2.925e+11Hz 0.428789 0.839414
+ 2.926e+11Hz 0.430298 0.838697
+ 2.927e+11Hz 0.431806 0.837976
+ 2.928e+11Hz 0.433315 0.837252
+ 2.929e+11Hz 0.434822 0.836524
+ 2.93e+11Hz 0.43633 0.835793
+ 2.931e+11Hz 0.437837 0.835059
+ 2.932e+11Hz 0.439344 0.834321
+ 2.933e+11Hz 0.44085 0.833579
+ 2.934e+11Hz 0.442355 0.832834
+ 2.935e+11Hz 0.44386 0.832085
+ 2.936e+11Hz 0.445365 0.831333
+ 2.937e+11Hz 0.446869 0.830577
+ 2.938e+11Hz 0.448372 0.829818
+ 2.939e+11Hz 0.449875 0.829055
+ 2.94e+11Hz 0.451377 0.828289
+ 2.941e+11Hz 0.452878 0.827519
+ 2.942e+11Hz 0.454379 0.826745
+ 2.943e+11Hz 0.455878 0.825968
+ 2.944e+11Hz 0.457377 0.825187
+ 2.945e+11Hz 0.458875 0.824403
+ 2.946e+11Hz 0.460372 0.823615
+ 2.947e+11Hz 0.461869 0.822824
+ 2.948e+11Hz 0.463364 0.822029
+ 2.949e+11Hz 0.464858 0.82123
+ 2.95e+11Hz 0.466351 0.820428
+ 2.951e+11Hz 0.467843 0.819622
+ 2.952e+11Hz 0.469335 0.818812
+ 2.953e+11Hz 0.470825 0.817999
+ 2.954e+11Hz 0.472314 0.817183
+ 2.955e+11Hz 0.473801 0.816362
+ 2.956e+11Hz 0.475288 0.815539
+ 2.957e+11Hz 0.476773 0.814711
+ 2.958e+11Hz 0.478257 0.813881
+ 2.959e+11Hz 0.47974 0.813046
+ 2.96e+11Hz 0.481221 0.812208
+ 2.961e+11Hz 0.482702 0.811367
+ 2.962e+11Hz 0.48418 0.810522
+ 2.963e+11Hz 0.485658 0.809674
+ 2.964e+11Hz 0.487134 0.808822
+ 2.965e+11Hz 0.488609 0.807966
+ 2.966e+11Hz 0.490082 0.807107
+ 2.967e+11Hz 0.491553 0.806245
+ 2.968e+11Hz 0.493023 0.805379
+ 2.969e+11Hz 0.494492 0.80451
+ 2.97e+11Hz 0.495959 0.803637
+ 2.971e+11Hz 0.497425 0.802761
+ 2.972e+11Hz 0.498889 0.801882
+ 2.973e+11Hz 0.500351 0.800999
+ 2.974e+11Hz 0.501812 0.800113
+ 2.975e+11Hz 0.503271 0.799224
+ 2.976e+11Hz 0.504728 0.798331
+ 2.977e+11Hz 0.506184 0.797435
+ 2.978e+11Hz 0.507638 0.796535
+ 2.979e+11Hz 0.50909 0.795632
+ 2.98e+11Hz 0.510541 0.794726
+ 2.981e+11Hz 0.51199 0.793817
+ 2.982e+11Hz 0.513437 0.792904
+ 2.983e+11Hz 0.514882 0.791989
+ 2.984e+11Hz 0.516326 0.79107
+ 2.985e+11Hz 0.517768 0.790148
+ 2.986e+11Hz 0.519207 0.789222
+ 2.987e+11Hz 0.520646 0.788294
+ 2.988e+11Hz 0.522082 0.787362
+ 2.989e+11Hz 0.523516 0.786427
+ 2.99e+11Hz 0.524949 0.785489
+ 2.991e+11Hz 0.52638 0.784548
+ 2.992e+11Hz 0.527809 0.783604
+ 2.993e+11Hz 0.529236 0.782657
+ 2.994e+11Hz 0.530661 0.781707
+ 2.995e+11Hz 0.532084 0.780754
+ 2.996e+11Hz 0.533505 0.779797
+ 2.997e+11Hz 0.534925 0.778838
+ 2.998e+11Hz 0.536342 0.777876
+ 2.999e+11Hz 0.537758 0.77691
+ 3e+11Hz 0.539172 0.775942
+ ]

A21 %vd(10 3) %vd(21, 22) xfer3
.model xfer3 xfer R_I=true table=[
+ 0Hz 0.990338 0
+ 1e+08Hz 0.990335 -0.0018782
+ 2e+08Hz 0.990326 -0.00375631
+ 3e+08Hz 0.990311 -0.00563423
+ 4e+08Hz 0.99029 -0.00751188
+ 5e+08Hz 0.990263 -0.00938916
+ 6e+08Hz 0.99023 -0.011266
+ 7e+08Hz 0.990191 -0.0131423
+ 8e+08Hz 0.990146 -0.0150179
+ 9e+08Hz 0.990096 -0.0168928
+ 1e+09Hz 0.990039 -0.0187669
+ 1.1e+09Hz 0.989977 -0.0206401
+ 1.2e+09Hz 0.989909 -0.0225123
+ 1.3e+09Hz 0.989835 -0.0243834
+ 1.4e+09Hz 0.989755 -0.0262534
+ 1.5e+09Hz 0.98967 -0.0281222
+ 1.6e+09Hz 0.989579 -0.0299896
+ 1.7e+09Hz 0.989482 -0.0318556
+ 1.8e+09Hz 0.98938 -0.0337202
+ 1.9e+09Hz 0.989272 -0.0355832
+ 2e+09Hz 0.989159 -0.0374446
+ 2.1e+09Hz 0.98904 -0.0393043
+ 2.2e+09Hz 0.988916 -0.0411622
+ 2.3e+09Hz 0.988787 -0.0430184
+ 2.4e+09Hz 0.988652 -0.0448726
+ 2.5e+09Hz 0.988513 -0.0467249
+ 2.6e+09Hz 0.988368 -0.0485752
+ 2.7e+09Hz 0.988218 -0.0504234
+ 2.8e+09Hz 0.988063 -0.0522695
+ 2.9e+09Hz 0.987903 -0.0541134
+ 3e+09Hz 0.987739 -0.0559551
+ 3.1e+09Hz 0.987569 -0.0577945
+ 3.2e+09Hz 0.987395 -0.0596316
+ 3.3e+09Hz 0.987217 -0.0614664
+ 3.4e+09Hz 0.987033 -0.0632987
+ 3.5e+09Hz 0.986846 -0.0651286
+ 3.6e+09Hz 0.986654 -0.0669561
+ 3.7e+09Hz 0.986457 -0.0687811
+ 3.8e+09Hz 0.986256 -0.0706035
+ 3.9e+09Hz 0.986052 -0.0724234
+ 4e+09Hz 0.985843 -0.0742408
+ 4.1e+09Hz 0.98563 -0.0760555
+ 4.2e+09Hz 0.985413 -0.0778677
+ 4.3e+09Hz 0.985192 -0.0796772
+ 4.4e+09Hz 0.984968 -0.0814841
+ 4.5e+09Hz 0.984739 -0.0832884
+ 4.6e+09Hz 0.984507 -0.08509
+ 4.7e+09Hz 0.984272 -0.0868889
+ 4.8e+09Hz 0.984033 -0.0886853
+ 4.9e+09Hz 0.983791 -0.090479
+ 5e+09Hz 0.983545 -0.09227
+ 5.1e+09Hz 0.983297 -0.0940584
+ 5.2e+09Hz 0.983045 -0.0958442
+ 5.3e+09Hz 0.982789 -0.0976274
+ 5.4e+09Hz 0.982531 -0.099408
+ 5.5e+09Hz 0.98227 -0.101186
+ 5.6e+09Hz 0.982006 -0.102962
+ 5.7e+09Hz 0.981739 -0.104734
+ 5.8e+09Hz 0.98147 -0.106505
+ 5.9e+09Hz 0.981197 -0.108273
+ 6e+09Hz 0.980923 -0.110038
+ 6.1e+09Hz 0.980645 -0.111801
+ 6.2e+09Hz 0.980365 -0.113562
+ 6.3e+09Hz 0.980083 -0.11532
+ 6.4e+09Hz 0.979798 -0.117076
+ 6.5e+09Hz 0.979511 -0.11883
+ 6.6e+09Hz 0.979221 -0.120582
+ 6.7e+09Hz 0.978929 -0.122331
+ 6.8e+09Hz 0.978635 -0.124078
+ 6.9e+09Hz 0.978339 -0.125823
+ 7e+09Hz 0.978041 -0.127566
+ 7.1e+09Hz 0.977741 -0.129307
+ 7.2e+09Hz 0.977439 -0.131046
+ 7.3e+09Hz 0.977134 -0.132783
+ 7.4e+09Hz 0.976828 -0.134518
+ 7.5e+09Hz 0.97652 -0.136251
+ 7.6e+09Hz 0.97621 -0.137982
+ 7.7e+09Hz 0.975898 -0.139712
+ 7.8e+09Hz 0.975585 -0.14144
+ 7.9e+09Hz 0.975269 -0.143166
+ 8e+09Hz 0.974952 -0.144891
+ 8.1e+09Hz 0.974633 -0.146614
+ 8.2e+09Hz 0.974312 -0.148336
+ 8.3e+09Hz 0.97399 -0.150056
+ 8.4e+09Hz 0.973666 -0.151775
+ 8.5e+09Hz 0.97334 -0.153493
+ 8.6e+09Hz 0.973012 -0.15521
+ 8.7e+09Hz 0.972683 -0.156925
+ 8.8e+09Hz 0.972352 -0.158639
+ 8.9e+09Hz 0.97202 -0.160352
+ 9e+09Hz 0.971685 -0.162063
+ 9.1e+09Hz 0.971349 -0.163774
+ 9.2e+09Hz 0.971012 -0.165484
+ 9.3e+09Hz 0.970672 -0.167193
+ 9.4e+09Hz 0.970331 -0.168901
+ 9.5e+09Hz 0.969989 -0.170609
+ 9.6e+09Hz 0.969644 -0.172315
+ 9.7e+09Hz 0.969298 -0.174021
+ 9.8e+09Hz 0.96895 -0.175726
+ 9.9e+09Hz 0.968601 -0.177431
+ 1e+10Hz 0.968249 -0.179135
+ 1.01e+10Hz 0.967896 -0.180838
+ 1.02e+10Hz 0.967541 -0.182541
+ 1.03e+10Hz 0.967184 -0.184243
+ 1.04e+10Hz 0.966825 -0.185946
+ 1.05e+10Hz 0.966464 -0.187647
+ 1.06e+10Hz 0.966102 -0.189348
+ 1.07e+10Hz 0.965737 -0.191049
+ 1.08e+10Hz 0.965371 -0.19275
+ 1.09e+10Hz 0.965002 -0.194451
+ 1.1e+10Hz 0.964632 -0.196151
+ 1.11e+10Hz 0.964259 -0.197851
+ 1.12e+10Hz 0.963884 -0.199551
+ 1.13e+10Hz 0.963507 -0.201251
+ 1.14e+10Hz 0.963128 -0.20295
+ 1.15e+10Hz 0.962747 -0.20465
+ 1.16e+10Hz 0.962363 -0.206349
+ 1.17e+10Hz 0.961977 -0.208049
+ 1.18e+10Hz 0.961589 -0.209748
+ 1.19e+10Hz 0.961198 -0.211448
+ 1.2e+10Hz 0.960805 -0.213147
+ 1.21e+10Hz 0.960409 -0.214846
+ 1.22e+10Hz 0.960011 -0.216546
+ 1.23e+10Hz 0.959611 -0.218245
+ 1.24e+10Hz 0.959207 -0.219944
+ 1.25e+10Hz 0.958802 -0.221644
+ 1.26e+10Hz 0.958393 -0.223343
+ 1.27e+10Hz 0.957982 -0.225042
+ 1.28e+10Hz 0.957568 -0.226742
+ 1.29e+10Hz 0.957151 -0.228441
+ 1.3e+10Hz 0.956731 -0.230141
+ 1.31e+10Hz 0.956309 -0.23184
+ 1.32e+10Hz 0.955884 -0.23354
+ 1.33e+10Hz 0.955455 -0.235239
+ 1.34e+10Hz 0.955024 -0.236938
+ 1.35e+10Hz 0.95459 -0.238638
+ 1.36e+10Hz 0.954152 -0.240337
+ 1.37e+10Hz 0.953712 -0.242036
+ 1.38e+10Hz 0.953268 -0.243735
+ 1.39e+10Hz 0.952821 -0.245434
+ 1.4e+10Hz 0.952371 -0.247133
+ 1.41e+10Hz 0.951918 -0.248832
+ 1.42e+10Hz 0.951461 -0.25053
+ 1.43e+10Hz 0.951001 -0.252228
+ 1.44e+10Hz 0.950538 -0.253927
+ 1.45e+10Hz 0.950071 -0.255624
+ 1.46e+10Hz 0.949601 -0.257322
+ 1.47e+10Hz 0.949128 -0.259019
+ 1.48e+10Hz 0.948651 -0.260716
+ 1.49e+10Hz 0.948171 -0.262412
+ 1.5e+10Hz 0.947687 -0.264108
+ 1.51e+10Hz 0.9472 -0.265803
+ 1.52e+10Hz 0.946709 -0.267498
+ 1.53e+10Hz 0.946215 -0.269193
+ 1.54e+10Hz 0.945717 -0.270886
+ 1.55e+10Hz 0.945215 -0.27258
+ 1.56e+10Hz 0.94471 -0.274272
+ 1.57e+10Hz 0.944201 -0.275964
+ 1.58e+10Hz 0.943689 -0.277655
+ 1.59e+10Hz 0.943173 -0.279346
+ 1.6e+10Hz 0.942653 -0.281035
+ 1.61e+10Hz 0.94213 -0.282724
+ 1.62e+10Hz 0.941603 -0.284412
+ 1.63e+10Hz 0.941073 -0.286099
+ 1.64e+10Hz 0.940539 -0.287785
+ 1.65e+10Hz 0.940001 -0.28947
+ 1.66e+10Hz 0.93946 -0.291154
+ 1.67e+10Hz 0.938914 -0.292837
+ 1.68e+10Hz 0.938366 -0.294519
+ 1.69e+10Hz 0.937813 -0.296199
+ 1.7e+10Hz 0.937258 -0.297878
+ 1.71e+10Hz 0.936698 -0.299557
+ 1.72e+10Hz 0.936135 -0.301233
+ 1.73e+10Hz 0.935568 -0.302909
+ 1.74e+10Hz 0.934998 -0.304583
+ 1.75e+10Hz 0.934424 -0.306256
+ 1.76e+10Hz 0.933847 -0.307927
+ 1.77e+10Hz 0.933266 -0.309597
+ 1.78e+10Hz 0.932682 -0.311266
+ 1.79e+10Hz 0.932094 -0.312933
+ 1.8e+10Hz 0.931503 -0.314598
+ 1.81e+10Hz 0.930908 -0.316262
+ 1.82e+10Hz 0.93031 -0.317924
+ 1.83e+10Hz 0.929708 -0.319585
+ 1.84e+10Hz 0.929104 -0.321244
+ 1.85e+10Hz 0.928495 -0.322901
+ 1.86e+10Hz 0.927884 -0.324556
+ 1.87e+10Hz 0.927269 -0.32621
+ 1.88e+10Hz 0.926651 -0.327862
+ 1.89e+10Hz 0.92603 -0.329512
+ 1.9e+10Hz 0.925406 -0.331161
+ 1.91e+10Hz 0.924778 -0.332807
+ 1.92e+10Hz 0.924148 -0.334452
+ 1.93e+10Hz 0.923514 -0.336095
+ 1.94e+10Hz 0.922877 -0.337736
+ 1.95e+10Hz 0.922238 -0.339375
+ 1.96e+10Hz 0.921595 -0.341012
+ 1.97e+10Hz 0.920949 -0.342647
+ 1.98e+10Hz 0.920301 -0.344281
+ 1.99e+10Hz 0.919649 -0.345912
+ 2e+10Hz 0.918995 -0.347542
+ 2.01e+10Hz 0.918338 -0.349169
+ 2.02e+10Hz 0.917678 -0.350795
+ 2.03e+10Hz 0.917015 -0.352419
+ 2.04e+10Hz 0.91635 -0.35404
+ 2.05e+10Hz 0.915682 -0.35566
+ 2.06e+10Hz 0.915011 -0.357278
+ 2.07e+10Hz 0.914338 -0.358894
+ 2.08e+10Hz 0.913662 -0.360508
+ 2.09e+10Hz 0.912984 -0.36212
+ 2.1e+10Hz 0.912303 -0.363731
+ 2.11e+10Hz 0.911619 -0.365339
+ 2.12e+10Hz 0.910933 -0.366945
+ 2.13e+10Hz 0.910245 -0.36855
+ 2.14e+10Hz 0.909554 -0.370152
+ 2.15e+10Hz 0.908861 -0.371753
+ 2.16e+10Hz 0.908166 -0.373352
+ 2.17e+10Hz 0.907468 -0.374949
+ 2.18e+10Hz 0.906768 -0.376545
+ 2.19e+10Hz 0.906066 -0.378138
+ 2.2e+10Hz 0.905362 -0.37973
+ 2.21e+10Hz 0.904655 -0.38132
+ 2.22e+10Hz 0.903946 -0.382908
+ 2.23e+10Hz 0.903235 -0.384495
+ 2.24e+10Hz 0.902522 -0.386079
+ 2.25e+10Hz 0.901806 -0.387663
+ 2.26e+10Hz 0.901089 -0.389244
+ 2.27e+10Hz 0.900369 -0.390824
+ 2.28e+10Hz 0.899647 -0.392402
+ 2.29e+10Hz 0.898924 -0.393979
+ 2.3e+10Hz 0.898198 -0.395554
+ 2.31e+10Hz 0.89747 -0.397128
+ 2.32e+10Hz 0.89674 -0.3987
+ 2.33e+10Hz 0.896008 -0.40027
+ 2.34e+10Hz 0.895274 -0.401839
+ 2.35e+10Hz 0.894538 -0.403407
+ 2.36e+10Hz 0.8938 -0.404973
+ 2.37e+10Hz 0.89306 -0.406538
+ 2.38e+10Hz 0.892318 -0.408102
+ 2.39e+10Hz 0.891573 -0.409664
+ 2.4e+10Hz 0.890827 -0.411225
+ 2.41e+10Hz 0.890079 -0.412785
+ 2.42e+10Hz 0.889329 -0.414343
+ 2.43e+10Hz 0.888577 -0.4159
+ 2.44e+10Hz 0.887823 -0.417456
+ 2.45e+10Hz 0.887066 -0.419011
+ 2.46e+10Hz 0.886308 -0.420565
+ 2.47e+10Hz 0.885548 -0.422117
+ 2.48e+10Hz 0.884785 -0.423669
+ 2.49e+10Hz 0.884021 -0.425219
+ 2.5e+10Hz 0.883254 -0.426768
+ 2.51e+10Hz 0.882486 -0.428316
+ 2.52e+10Hz 0.881715 -0.429864
+ 2.53e+10Hz 0.880942 -0.43141
+ 2.54e+10Hz 0.880167 -0.432955
+ 2.55e+10Hz 0.87939 -0.434499
+ 2.56e+10Hz 0.87861 -0.436043
+ 2.57e+10Hz 0.877829 -0.437585
+ 2.58e+10Hz 0.877045 -0.439126
+ 2.59e+10Hz 0.876259 -0.440667
+ 2.6e+10Hz 0.875471 -0.442207
+ 2.61e+10Hz 0.87468 -0.443745
+ 2.62e+10Hz 0.873887 -0.445283
+ 2.63e+10Hz 0.873092 -0.44682
+ 2.64e+10Hz 0.872295 -0.448357
+ 2.65e+10Hz 0.871495 -0.449892
+ 2.66e+10Hz 0.870693 -0.451427
+ 2.67e+10Hz 0.869888 -0.45296
+ 2.68e+10Hz 0.869081 -0.454493
+ 2.69e+10Hz 0.868271 -0.456025
+ 2.7e+10Hz 0.867459 -0.457557
+ 2.71e+10Hz 0.866645 -0.459087
+ 2.72e+10Hz 0.865827 -0.460617
+ 2.73e+10Hz 0.865008 -0.462146
+ 2.74e+10Hz 0.864185 -0.463674
+ 2.75e+10Hz 0.86336 -0.465201
+ 2.76e+10Hz 0.862533 -0.466727
+ 2.77e+10Hz 0.861703 -0.468253
+ 2.78e+10Hz 0.86087 -0.469778
+ 2.79e+10Hz 0.860034 -0.471302
+ 2.8e+10Hz 0.859196 -0.472825
+ 2.81e+10Hz 0.858354 -0.474347
+ 2.82e+10Hz 0.85751 -0.475868
+ 2.83e+10Hz 0.856663 -0.477389
+ 2.84e+10Hz 0.855814 -0.478908
+ 2.85e+10Hz 0.854961 -0.480427
+ 2.86e+10Hz 0.854106 -0.481944
+ 2.87e+10Hz 0.853247 -0.483461
+ 2.88e+10Hz 0.852386 -0.484977
+ 2.89e+10Hz 0.851522 -0.486492
+ 2.9e+10Hz 0.850654 -0.488006
+ 2.91e+10Hz 0.849784 -0.489519
+ 2.92e+10Hz 0.848911 -0.49103
+ 2.93e+10Hz 0.848035 -0.492541
+ 2.94e+10Hz 0.847155 -0.494051
+ 2.95e+10Hz 0.846273 -0.495559
+ 2.96e+10Hz 0.845387 -0.497067
+ 2.97e+10Hz 0.844498 -0.498573
+ 2.98e+10Hz 0.843606 -0.500078
+ 2.99e+10Hz 0.842711 -0.501582
+ 3e+10Hz 0.841813 -0.503085
+ 3.01e+10Hz 0.840912 -0.504586
+ 3.02e+10Hz 0.840008 -0.506086
+ 3.03e+10Hz 0.8391 -0.507585
+ 3.04e+10Hz 0.838189 -0.509082
+ 3.05e+10Hz 0.837275 -0.510578
+ 3.06e+10Hz 0.836358 -0.512073
+ 3.07e+10Hz 0.835437 -0.513566
+ 3.08e+10Hz 0.834513 -0.515058
+ 3.09e+10Hz 0.833587 -0.516548
+ 3.1e+10Hz 0.832656 -0.518037
+ 3.11e+10Hz 0.831723 -0.519524
+ 3.12e+10Hz 0.830786 -0.521009
+ 3.13e+10Hz 0.829847 -0.522493
+ 3.14e+10Hz 0.828903 -0.523975
+ 3.15e+10Hz 0.827957 -0.525456
+ 3.16e+10Hz 0.827008 -0.526935
+ 3.17e+10Hz 0.826055 -0.528412
+ 3.18e+10Hz 0.825099 -0.529887
+ 3.19e+10Hz 0.82414 -0.531361
+ 3.2e+10Hz 0.823177 -0.532833
+ 3.21e+10Hz 0.822212 -0.534302
+ 3.22e+10Hz 0.821243 -0.53577
+ 3.23e+10Hz 0.820271 -0.537236
+ 3.24e+10Hz 0.819296 -0.5387
+ 3.25e+10Hz 0.818318 -0.540162
+ 3.26e+10Hz 0.817337 -0.541622
+ 3.27e+10Hz 0.816353 -0.54308
+ 3.28e+10Hz 0.815365 -0.544536
+ 3.29e+10Hz 0.814375 -0.54599
+ 3.3e+10Hz 0.813381 -0.547442
+ 3.31e+10Hz 0.812385 -0.548892
+ 3.32e+10Hz 0.811385 -0.550339
+ 3.33e+10Hz 0.810382 -0.551784
+ 3.34e+10Hz 0.809377 -0.553227
+ 3.35e+10Hz 0.808368 -0.554668
+ 3.36e+10Hz 0.807357 -0.556107
+ 3.37e+10Hz 0.806343 -0.557543
+ 3.38e+10Hz 0.805325 -0.558977
+ 3.39e+10Hz 0.804305 -0.560408
+ 3.4e+10Hz 0.803282 -0.561838
+ 3.41e+10Hz 0.802257 -0.563265
+ 3.42e+10Hz 0.801228 -0.564689
+ 3.43e+10Hz 0.800197 -0.566112
+ 3.44e+10Hz 0.799163 -0.567531
+ 3.45e+10Hz 0.798126 -0.568949
+ 3.46e+10Hz 0.797087 -0.570364
+ 3.47e+10Hz 0.796045 -0.571777
+ 3.48e+10Hz 0.795 -0.573187
+ 3.49e+10Hz 0.793953 -0.574594
+ 3.5e+10Hz 0.792903 -0.576
+ 3.51e+10Hz 0.791851 -0.577403
+ 3.52e+10Hz 0.790796 -0.578803
+ 3.53e+10Hz 0.789738 -0.580201
+ 3.54e+10Hz 0.788679 -0.581596
+ 3.55e+10Hz 0.787616 -0.582989
+ 3.56e+10Hz 0.786552 -0.58438
+ 3.57e+10Hz 0.785485 -0.585768
+ 3.58e+10Hz 0.784415 -0.587153
+ 3.59e+10Hz 0.783344 -0.588536
+ 3.6e+10Hz 0.78227 -0.589917
+ 3.61e+10Hz 0.781194 -0.591295
+ 3.62e+10Hz 0.780115 -0.592671
+ 3.63e+10Hz 0.779035 -0.594044
+ 3.64e+10Hz 0.777952 -0.595415
+ 3.65e+10Hz 0.776867 -0.596783
+ 3.66e+10Hz 0.77578 -0.598149
+ 3.67e+10Hz 0.77469 -0.599512
+ 3.68e+10Hz 0.773599 -0.600873
+ 3.69e+10Hz 0.772506 -0.602232
+ 3.7e+10Hz 0.77141 -0.603588
+ 3.71e+10Hz 0.770313 -0.604942
+ 3.72e+10Hz 0.769213 -0.606294
+ 3.73e+10Hz 0.768112 -0.607643
+ 3.74e+10Hz 0.767008 -0.60899
+ 3.75e+10Hz 0.765903 -0.610334
+ 3.76e+10Hz 0.764795 -0.611676
+ 3.77e+10Hz 0.763686 -0.613016
+ 3.78e+10Hz 0.762575 -0.614354
+ 3.79e+10Hz 0.761462 -0.615689
+ 3.8e+10Hz 0.760347 -0.617022
+ 3.81e+10Hz 0.75923 -0.618353
+ 3.82e+10Hz 0.758111 -0.619682
+ 3.83e+10Hz 0.756991 -0.621008
+ 3.84e+10Hz 0.755869 -0.622332
+ 3.85e+10Hz 0.754744 -0.623654
+ 3.86e+10Hz 0.753619 -0.624974
+ 3.87e+10Hz 0.752491 -0.626292
+ 3.88e+10Hz 0.751361 -0.627608
+ 3.89e+10Hz 0.75023 -0.628921
+ 3.9e+10Hz 0.749097 -0.630233
+ 3.91e+10Hz 0.747962 -0.631542
+ 3.92e+10Hz 0.746825 -0.63285
+ 3.93e+10Hz 0.745687 -0.634155
+ 3.94e+10Hz 0.744546 -0.635458
+ 3.95e+10Hz 0.743404 -0.63676
+ 3.96e+10Hz 0.74226 -0.638059
+ 3.97e+10Hz 0.741115 -0.639357
+ 3.98e+10Hz 0.739968 -0.640652
+ 3.99e+10Hz 0.738818 -0.641946
+ 4e+10Hz 0.737667 -0.643238
+ 4.01e+10Hz 0.736515 -0.644528
+ 4.02e+10Hz 0.73536 -0.645816
+ 4.03e+10Hz 0.734204 -0.647102
+ 4.04e+10Hz 0.733046 -0.648387
+ 4.05e+10Hz 0.731886 -0.649669
+ 4.06e+10Hz 0.730724 -0.65095
+ 4.07e+10Hz 0.72956 -0.652229
+ 4.08e+10Hz 0.728395 -0.653506
+ 4.09e+10Hz 0.727227 -0.654782
+ 4.1e+10Hz 0.726058 -0.656055
+ 4.11e+10Hz 0.724887 -0.657327
+ 4.12e+10Hz 0.723714 -0.658597
+ 4.13e+10Hz 0.722539 -0.659866
+ 4.14e+10Hz 0.721362 -0.661133
+ 4.15e+10Hz 0.720183 -0.662398
+ 4.16e+10Hz 0.719003 -0.663661
+ 4.17e+10Hz 0.71782 -0.664923
+ 4.18e+10Hz 0.716635 -0.666183
+ 4.19e+10Hz 0.715449 -0.667442
+ 4.2e+10Hz 0.71426 -0.668698
+ 4.21e+10Hz 0.713069 -0.669953
+ 4.22e+10Hz 0.711876 -0.671207
+ 4.23e+10Hz 0.710682 -0.672458
+ 4.24e+10Hz 0.709485 -0.673708
+ 4.25e+10Hz 0.708286 -0.674957
+ 4.26e+10Hz 0.707085 -0.676204
+ 4.27e+10Hz 0.705881 -0.677449
+ 4.28e+10Hz 0.704676 -0.678692
+ 4.29e+10Hz 0.703468 -0.679934
+ 4.3e+10Hz 0.702259 -0.681174
+ 4.31e+10Hz 0.701047 -0.682412
+ 4.32e+10Hz 0.699833 -0.683649
+ 4.33e+10Hz 0.698616 -0.684884
+ 4.34e+10Hz 0.697398 -0.686117
+ 4.35e+10Hz 0.696177 -0.687349
+ 4.36e+10Hz 0.694954 -0.688579
+ 4.37e+10Hz 0.693728 -0.689807
+ 4.38e+10Hz 0.6925 -0.691033
+ 4.39e+10Hz 0.69127 -0.692258
+ 4.4e+10Hz 0.690038 -0.693481
+ 4.41e+10Hz 0.688803 -0.694702
+ 4.42e+10Hz 0.687566 -0.695922
+ 4.43e+10Hz 0.686326 -0.697139
+ 4.44e+10Hz 0.685084 -0.698355
+ 4.45e+10Hz 0.68384 -0.699569
+ 4.46e+10Hz 0.682593 -0.700781
+ 4.47e+10Hz 0.681344 -0.701991
+ 4.48e+10Hz 0.680092 -0.7032
+ 4.49e+10Hz 0.678838 -0.704406
+ 4.5e+10Hz 0.677582 -0.705611
+ 4.51e+10Hz 0.676322 -0.706814
+ 4.52e+10Hz 0.675061 -0.708014
+ 4.53e+10Hz 0.673797 -0.709213
+ 4.54e+10Hz 0.67253 -0.71041
+ 4.55e+10Hz 0.671261 -0.711605
+ 4.56e+10Hz 0.66999 -0.712798
+ 4.57e+10Hz 0.668716 -0.713988
+ 4.58e+10Hz 0.667439 -0.715177
+ 4.59e+10Hz 0.66616 -0.716363
+ 4.6e+10Hz 0.664878 -0.717548
+ 4.61e+10Hz 0.663594 -0.71873
+ 4.62e+10Hz 0.662307 -0.71991
+ 4.63e+10Hz 0.661018 -0.721088
+ 4.64e+10Hz 0.659726 -0.722264
+ 4.65e+10Hz 0.658432 -0.723437
+ 4.66e+10Hz 0.657135 -0.724609
+ 4.67e+10Hz 0.655836 -0.725778
+ 4.68e+10Hz 0.654534 -0.726944
+ 4.69e+10Hz 0.65323 -0.728109
+ 4.7e+10Hz 0.651923 -0.729271
+ 4.71e+10Hz 0.650613 -0.730431
+ 4.72e+10Hz 0.649302 -0.731588
+ 4.73e+10Hz 0.647987 -0.732743
+ 4.74e+10Hz 0.64667 -0.733895
+ 4.75e+10Hz 0.645351 -0.735045
+ 4.76e+10Hz 0.644029 -0.736193
+ 4.77e+10Hz 0.642705 -0.737338
+ 4.78e+10Hz 0.641378 -0.73848
+ 4.79e+10Hz 0.640049 -0.73962
+ 4.8e+10Hz 0.638717 -0.740758
+ 4.81e+10Hz 0.637383 -0.741893
+ 4.82e+10Hz 0.636047 -0.743025
+ 4.83e+10Hz 0.634708 -0.744155
+ 4.84e+10Hz 0.633367 -0.745282
+ 4.85e+10Hz 0.632023 -0.746406
+ 4.86e+10Hz 0.630678 -0.747528
+ 4.87e+10Hz 0.629329 -0.748647
+ 4.88e+10Hz 0.627979 -0.749763
+ 4.89e+10Hz 0.626626 -0.750877
+ 4.9e+10Hz 0.625271 -0.751988
+ 4.91e+10Hz 0.623914 -0.753096
+ 4.92e+10Hz 0.622554 -0.754201
+ 4.93e+10Hz 0.621193 -0.755304
+ 4.94e+10Hz 0.619829 -0.756403
+ 4.95e+10Hz 0.618463 -0.7575
+ 4.96e+10Hz 0.617095 -0.758595
+ 4.97e+10Hz 0.615724 -0.759686
+ 4.98e+10Hz 0.614352 -0.760775
+ 4.99e+10Hz 0.612977 -0.76186
+ 5e+10Hz 0.6116 -0.762943
+ 5.01e+10Hz 0.610222 -0.764023
+ 5.02e+10Hz 0.608841 -0.7651
+ 5.03e+10Hz 0.607458 -0.766174
+ 5.04e+10Hz 0.606074 -0.767246
+ 5.05e+10Hz 0.604687 -0.768314
+ 5.06e+10Hz 0.603298 -0.76938
+ 5.07e+10Hz 0.601908 -0.770443
+ 5.08e+10Hz 0.600515 -0.771503
+ 5.09e+10Hz 0.599121 -0.772559
+ 5.1e+10Hz 0.597725 -0.773613
+ 5.11e+10Hz 0.596327 -0.774665
+ 5.12e+10Hz 0.594927 -0.775713
+ 5.13e+10Hz 0.593526 -0.776758
+ 5.14e+10Hz 0.592122 -0.777801
+ 5.15e+10Hz 0.590717 -0.77884
+ 5.16e+10Hz 0.58931 -0.779877
+ 5.17e+10Hz 0.587902 -0.780911
+ 5.18e+10Hz 0.586492 -0.781942
+ 5.19e+10Hz 0.58508 -0.78297
+ 5.2e+10Hz 0.583666 -0.783995
+ 5.21e+10Hz 0.582251 -0.785017
+ 5.22e+10Hz 0.580834 -0.786036
+ 5.23e+10Hz 0.579416 -0.787053
+ 5.24e+10Hz 0.577996 -0.788067
+ 5.25e+10Hz 0.576574 -0.789077
+ 5.26e+10Hz 0.575151 -0.790085
+ 5.27e+10Hz 0.573726 -0.791091
+ 5.28e+10Hz 0.5723 -0.792093
+ 5.29e+10Hz 0.570872 -0.793093
+ 5.3e+10Hz 0.569443 -0.794089
+ 5.31e+10Hz 0.568013 -0.795084
+ 5.32e+10Hz 0.566581 -0.796075
+ 5.33e+10Hz 0.565147 -0.797063
+ 5.34e+10Hz 0.563712 -0.798049
+ 5.35e+10Hz 0.562276 -0.799032
+ 5.36e+10Hz 0.560838 -0.800012
+ 5.37e+10Hz 0.559399 -0.80099
+ 5.38e+10Hz 0.557958 -0.801965
+ 5.39e+10Hz 0.556516 -0.802937
+ 5.4e+10Hz 0.555072 -0.803906
+ 5.41e+10Hz 0.553628 -0.804873
+ 5.42e+10Hz 0.552181 -0.805837
+ 5.43e+10Hz 0.550734 -0.806799
+ 5.44e+10Hz 0.549285 -0.807758
+ 5.45e+10Hz 0.547835 -0.808714
+ 5.46e+10Hz 0.546383 -0.809668
+ 5.47e+10Hz 0.54493 -0.810619
+ 5.48e+10Hz 0.543476 -0.811567
+ 5.49e+10Hz 0.54202 -0.812513
+ 5.5e+10Hz 0.540563 -0.813457
+ 5.51e+10Hz 0.539105 -0.814397
+ 5.52e+10Hz 0.537645 -0.815336
+ 5.53e+10Hz 0.536184 -0.816272
+ 5.54e+10Hz 0.534722 -0.817205
+ 5.55e+10Hz 0.533258 -0.818136
+ 5.56e+10Hz 0.531793 -0.819064
+ 5.57e+10Hz 0.530327 -0.81999
+ 5.58e+10Hz 0.528859 -0.820913
+ 5.59e+10Hz 0.52739 -0.821834
+ 5.6e+10Hz 0.52592 -0.822753
+ 5.61e+10Hz 0.524448 -0.823669
+ 5.62e+10Hz 0.522975 -0.824582
+ 5.63e+10Hz 0.5215 -0.825494
+ 5.64e+10Hz 0.520024 -0.826402
+ 5.65e+10Hz 0.518547 -0.827309
+ 5.66e+10Hz 0.517068 -0.828213
+ 5.67e+10Hz 0.515588 -0.829115
+ 5.68e+10Hz 0.514106 -0.830014
+ 5.69e+10Hz 0.512623 -0.830911
+ 5.7e+10Hz 0.511139 -0.831805
+ 5.71e+10Hz 0.509653 -0.832697
+ 5.72e+10Hz 0.508166 -0.833587
+ 5.73e+10Hz 0.506677 -0.834475
+ 5.74e+10Hz 0.505187 -0.83536
+ 5.75e+10Hz 0.503695 -0.836242
+ 5.76e+10Hz 0.502202 -0.837123
+ 5.77e+10Hz 0.500707 -0.838001
+ 5.78e+10Hz 0.499211 -0.838876
+ 5.79e+10Hz 0.497713 -0.83975
+ 5.8e+10Hz 0.496214 -0.840621
+ 5.81e+10Hz 0.494713 -0.841489
+ 5.82e+10Hz 0.493211 -0.842356
+ 5.83e+10Hz 0.491707 -0.843219
+ 5.84e+10Hz 0.490201 -0.844081
+ 5.85e+10Hz 0.488694 -0.84494
+ 5.86e+10Hz 0.487186 -0.845797
+ 5.87e+10Hz 0.485675 -0.846651
+ 5.88e+10Hz 0.484163 -0.847503
+ 5.89e+10Hz 0.48265 -0.848353
+ 5.9e+10Hz 0.481135 -0.8492
+ 5.91e+10Hz 0.479618 -0.850045
+ 5.92e+10Hz 0.4781 -0.850887
+ 5.93e+10Hz 0.476579 -0.851727
+ 5.94e+10Hz 0.475058 -0.852565
+ 5.95e+10Hz 0.473534 -0.8534
+ 5.96e+10Hz 0.472009 -0.854232
+ 5.97e+10Hz 0.470482 -0.855062
+ 5.98e+10Hz 0.468954 -0.85589
+ 5.99e+10Hz 0.467423 -0.856715
+ 6e+10Hz 0.465891 -0.857538
+ 6.01e+10Hz 0.464358 -0.858358
+ 6.02e+10Hz 0.462822 -0.859176
+ 6.03e+10Hz 0.461285 -0.859991
+ 6.04e+10Hz 0.459746 -0.860803
+ 6.05e+10Hz 0.458205 -0.861613
+ 6.06e+10Hz 0.456663 -0.862421
+ 6.07e+10Hz 0.455119 -0.863225
+ 6.08e+10Hz 0.453573 -0.864028
+ 6.09e+10Hz 0.452025 -0.864827
+ 6.1e+10Hz 0.450475 -0.865624
+ 6.11e+10Hz 0.448924 -0.866418
+ 6.12e+10Hz 0.447371 -0.86721
+ 6.13e+10Hz 0.445816 -0.867999
+ 6.14e+10Hz 0.44426 -0.868785
+ 6.15e+10Hz 0.442702 -0.869568
+ 6.16e+10Hz 0.441141 -0.870349
+ 6.17e+10Hz 0.43958 -0.871127
+ 6.18e+10Hz 0.438016 -0.871902
+ 6.19e+10Hz 0.436451 -0.872674
+ 6.2e+10Hz 0.434883 -0.873443
+ 6.21e+10Hz 0.433315 -0.87421
+ 6.22e+10Hz 0.431744 -0.874974
+ 6.23e+10Hz 0.430172 -0.875734
+ 6.24e+10Hz 0.428597 -0.876492
+ 6.25e+10Hz 0.427022 -0.877247
+ 6.26e+10Hz 0.425444 -0.878
+ 6.27e+10Hz 0.423865 -0.878749
+ 6.28e+10Hz 0.422284 -0.879495
+ 6.29e+10Hz 0.420701 -0.880238
+ 6.3e+10Hz 0.419117 -0.880978
+ 6.31e+10Hz 0.417531 -0.881716
+ 6.32e+10Hz 0.415943 -0.88245
+ 6.33e+10Hz 0.414354 -0.883181
+ 6.34e+10Hz 0.412763 -0.883909
+ 6.35e+10Hz 0.41117 -0.884634
+ 6.36e+10Hz 0.409576 -0.885356
+ 6.37e+10Hz 0.40798 -0.886075
+ 6.38e+10Hz 0.406382 -0.88679
+ 6.39e+10Hz 0.404783 -0.887503
+ 6.4e+10Hz 0.403183 -0.888212
+ 6.41e+10Hz 0.401581 -0.888918
+ 6.42e+10Hz 0.399977 -0.889621
+ 6.43e+10Hz 0.398372 -0.890321
+ 6.44e+10Hz 0.396765 -0.891018
+ 6.45e+10Hz 0.395157 -0.891711
+ 6.46e+10Hz 0.393547 -0.892401
+ 6.47e+10Hz 0.391936 -0.893088
+ 6.48e+10Hz 0.390324 -0.893772
+ 6.49e+10Hz 0.38871 -0.894452
+ 6.5e+10Hz 0.387094 -0.895129
+ 6.51e+10Hz 0.385477 -0.895803
+ 6.52e+10Hz 0.383859 -0.896473
+ 6.53e+10Hz 0.38224 -0.89714
+ 6.54e+10Hz 0.380619 -0.897804
+ 6.55e+10Hz 0.378997 -0.898465
+ 6.56e+10Hz 0.377374 -0.899122
+ 6.57e+10Hz 0.375749 -0.899776
+ 6.58e+10Hz 0.374123 -0.900427
+ 6.59e+10Hz 0.372496 -0.901074
+ 6.6e+10Hz 0.370868 -0.901718
+ 6.61e+10Hz 0.369238 -0.902358
+ 6.62e+10Hz 0.367608 -0.902996
+ 6.63e+10Hz 0.365976 -0.90363
+ 6.64e+10Hz 0.364343 -0.90426
+ 6.65e+10Hz 0.362709 -0.904887
+ 6.66e+10Hz 0.361074 -0.905511
+ 6.67e+10Hz 0.359437 -0.906131
+ 6.68e+10Hz 0.3578 -0.906748
+ 6.69e+10Hz 0.356162 -0.907362
+ 6.7e+10Hz 0.354522 -0.907973
+ 6.71e+10Hz 0.352882 -0.90858
+ 6.72e+10Hz 0.351241 -0.909183
+ 6.73e+10Hz 0.349599 -0.909783
+ 6.74e+10Hz 0.347955 -0.91038
+ 6.75e+10Hz 0.346311 -0.910974
+ 6.76e+10Hz 0.344666 -0.911564
+ 6.77e+10Hz 0.34302 -0.912151
+ 6.78e+10Hz 0.341373 -0.912735
+ 6.79e+10Hz 0.339726 -0.913315
+ 6.8e+10Hz 0.338077 -0.913892
+ 6.81e+10Hz 0.336428 -0.914466
+ 6.82e+10Hz 0.334778 -0.915036
+ 6.83e+10Hz 0.333127 -0.915603
+ 6.84e+10Hz 0.331475 -0.916167
+ 6.85e+10Hz 0.329823 -0.916727
+ 6.86e+10Hz 0.32817 -0.917284
+ 6.87e+10Hz 0.326516 -0.917838
+ 6.88e+10Hz 0.324861 -0.918389
+ 6.89e+10Hz 0.323206 -0.918936
+ 6.9e+10Hz 0.32155 -0.91948
+ 6.91e+10Hz 0.319893 -0.920021
+ 6.92e+10Hz 0.318236 -0.920559
+ 6.93e+10Hz 0.316578 -0.921093
+ 6.94e+10Hz 0.314919 -0.921625
+ 6.95e+10Hz 0.31326 -0.922153
+ 6.96e+10Hz 0.3116 -0.922678
+ 6.97e+10Hz 0.309939 -0.923199
+ 6.98e+10Hz 0.308278 -0.923718
+ 6.99e+10Hz 0.306616 -0.924233
+ 7e+10Hz 0.304954 -0.924745
+ 7.01e+10Hz 0.303291 -0.925255
+ 7.02e+10Hz 0.301627 -0.92576
+ 7.03e+10Hz 0.299963 -0.926263
+ 7.04e+10Hz 0.298298 -0.926763
+ 7.05e+10Hz 0.296633 -0.92726
+ 7.06e+10Hz 0.294967 -0.927753
+ 7.07e+10Hz 0.2933 -0.928244
+ 7.08e+10Hz 0.291634 -0.928731
+ 7.09e+10Hz 0.289966 -0.929215
+ 7.1e+10Hz 0.288298 -0.929697
+ 7.11e+10Hz 0.286629 -0.930175
+ 7.12e+10Hz 0.28496 -0.93065
+ 7.13e+10Hz 0.28329 -0.931122
+ 7.14e+10Hz 0.28162 -0.931592
+ 7.15e+10Hz 0.279949 -0.932058
+ 7.16e+10Hz 0.278278 -0.932521
+ 7.17e+10Hz 0.276606 -0.932981
+ 7.18e+10Hz 0.274934 -0.933438
+ 7.19e+10Hz 0.273261 -0.933892
+ 7.2e+10Hz 0.271587 -0.934344
+ 7.21e+10Hz 0.269913 -0.934792
+ 7.22e+10Hz 0.268239 -0.935237
+ 7.23e+10Hz 0.266564 -0.93568
+ 7.24e+10Hz 0.264888 -0.936119
+ 7.25e+10Hz 0.263212 -0.936556
+ 7.26e+10Hz 0.261535 -0.936989
+ 7.27e+10Hz 0.259858 -0.93742
+ 7.28e+10Hz 0.25818 -0.937848
+ 7.29e+10Hz 0.256502 -0.938272
+ 7.3e+10Hz 0.254823 -0.938694
+ 7.31e+10Hz 0.253143 -0.939113
+ 7.32e+10Hz 0.251463 -0.939529
+ 7.33e+10Hz 0.249782 -0.939942
+ 7.34e+10Hz 0.248101 -0.940353
+ 7.35e+10Hz 0.246419 -0.94076
+ 7.36e+10Hz 0.244737 -0.941164
+ 7.37e+10Hz 0.243054 -0.941566
+ 7.38e+10Hz 0.24137 -0.941964
+ 7.39e+10Hz 0.239686 -0.94236
+ 7.4e+10Hz 0.238001 -0.942753
+ 7.41e+10Hz 0.236315 -0.943143
+ 7.42e+10Hz 0.234629 -0.94353
+ 7.43e+10Hz 0.232943 -0.943914
+ 7.44e+10Hz 0.231255 -0.944295
+ 7.45e+10Hz 0.229568 -0.944673
+ 7.46e+10Hz 0.227879 -0.945048
+ 7.47e+10Hz 0.22619 -0.94542
+ 7.48e+10Hz 0.2245 -0.94579
+ 7.49e+10Hz 0.22281 -0.946156
+ 7.5e+10Hz 0.221119 -0.94652
+ 7.51e+10Hz 0.219427 -0.94688
+ 7.52e+10Hz 0.217735 -0.947238
+ 7.53e+10Hz 0.216042 -0.947592
+ 7.54e+10Hz 0.214348 -0.947944
+ 7.55e+10Hz 0.212654 -0.948293
+ 7.56e+10Hz 0.210959 -0.948638
+ 7.57e+10Hz 0.209263 -0.948981
+ 7.58e+10Hz 0.207567 -0.949321
+ 7.59e+10Hz 0.20587 -0.949657
+ 7.6e+10Hz 0.204172 -0.949991
+ 7.61e+10Hz 0.202474 -0.950322
+ 7.62e+10Hz 0.200775 -0.950649
+ 7.63e+10Hz 0.199076 -0.950974
+ 7.64e+10Hz 0.197376 -0.951295
+ 7.65e+10Hz 0.195675 -0.951614
+ 7.66e+10Hz 0.193973 -0.951929
+ 7.67e+10Hz 0.192271 -0.952241
+ 7.68e+10Hz 0.190569 -0.952551
+ 7.69e+10Hz 0.188865 -0.952857
+ 7.7e+10Hz 0.187161 -0.95316
+ 7.71e+10Hz 0.185457 -0.95346
+ 7.72e+10Hz 0.183751 -0.953756
+ 7.73e+10Hz 0.182045 -0.95405
+ 7.74e+10Hz 0.180339 -0.95434
+ 7.75e+10Hz 0.178632 -0.954627
+ 7.76e+10Hz 0.176924 -0.954911
+ 7.77e+10Hz 0.175216 -0.955192
+ 7.78e+10Hz 0.173507 -0.95547
+ 7.79e+10Hz 0.171797 -0.955744
+ 7.8e+10Hz 0.170087 -0.956016
+ 7.81e+10Hz 0.168377 -0.956284
+ 7.82e+10Hz 0.166665 -0.956548
+ 7.83e+10Hz 0.164954 -0.95681
+ 7.84e+10Hz 0.163241 -0.957068
+ 7.85e+10Hz 0.161529 -0.957323
+ 7.86e+10Hz 0.159815 -0.957574
+ 7.87e+10Hz 0.158101 -0.957823
+ 7.88e+10Hz 0.156387 -0.958068
+ 7.89e+10Hz 0.154672 -0.958309
+ 7.9e+10Hz 0.152957 -0.958548
+ 7.91e+10Hz 0.151241 -0.958783
+ 7.92e+10Hz 0.149525 -0.959014
+ 7.93e+10Hz 0.147808 -0.959243
+ 7.94e+10Hz 0.146091 -0.959468
+ 7.95e+10Hz 0.144374 -0.959689
+ 7.96e+10Hz 0.142656 -0.959907
+ 7.97e+10Hz 0.140938 -0.960122
+ 7.98e+10Hz 0.139219 -0.960334
+ 7.99e+10Hz 0.1375 -0.960542
+ 8e+10Hz 0.135781 -0.960746
+ 8.01e+10Hz 0.134062 -0.960947
+ 8.02e+10Hz 0.132342 -0.961145
+ 8.03e+10Hz 0.130622 -0.96134
+ 8.04e+10Hz 0.128901 -0.96153
+ 8.05e+10Hz 0.127181 -0.961718
+ 8.06e+10Hz 0.12546 -0.961902
+ 8.07e+10Hz 0.123739 -0.962082
+ 8.08e+10Hz 0.122017 -0.962259
+ 8.09e+10Hz 0.120296 -0.962433
+ 8.1e+10Hz 0.118574 -0.962603
+ 8.11e+10Hz 0.116852 -0.96277
+ 8.12e+10Hz 0.11513 -0.962933
+ 8.13e+10Hz 0.113408 -0.963093
+ 8.14e+10Hz 0.111686 -0.963249
+ 8.15e+10Hz 0.109964 -0.963402
+ 8.16e+10Hz 0.108242 -0.963552
+ 8.17e+10Hz 0.10652 -0.963698
+ 8.18e+10Hz 0.104797 -0.96384
+ 8.19e+10Hz 0.103075 -0.963979
+ 8.2e+10Hz 0.101353 -0.964115
+ 8.21e+10Hz 0.0996305 -0.964247
+ 8.22e+10Hz 0.0979083 -0.964375
+ 8.23e+10Hz 0.0961862 -0.9645
+ 8.24e+10Hz 0.0944642 -0.964622
+ 8.25e+10Hz 0.0927423 -0.96474
+ 8.26e+10Hz 0.0910205 -0.964855
+ 8.27e+10Hz 0.0892989 -0.964966
+ 8.28e+10Hz 0.0875775 -0.965074
+ 8.29e+10Hz 0.0858562 -0.965179
+ 8.3e+10Hz 0.0841352 -0.96528
+ 8.31e+10Hz 0.0824143 -0.965377
+ 8.32e+10Hz 0.0806937 -0.965472
+ 8.33e+10Hz 0.0789734 -0.965563
+ 8.34e+10Hz 0.0772533 -0.96565
+ 8.35e+10Hz 0.0755335 -0.965734
+ 8.36e+10Hz 0.073814 -0.965815
+ 8.37e+10Hz 0.0720948 -0.965892
+ 8.38e+10Hz 0.0703759 -0.965966
+ 8.39e+10Hz 0.0686575 -0.966036
+ 8.4e+10Hz 0.0669393 -0.966103
+ 8.41e+10Hz 0.0652216 -0.966167
+ 8.42e+10Hz 0.0635042 -0.966228
+ 8.43e+10Hz 0.0617873 -0.966285
+ 8.44e+10Hz 0.0600707 -0.966339
+ 8.45e+10Hz 0.0583546 -0.966389
+ 8.46e+10Hz 0.056639 -0.966437
+ 8.47e+10Hz 0.0549238 -0.966481
+ 8.48e+10Hz 0.0532091 -0.966522
+ 8.49e+10Hz 0.0514949 -0.966559
+ 8.5e+10Hz 0.0497812 -0.966593
+ 8.51e+10Hz 0.048068 -0.966624
+ 8.52e+10Hz 0.0463553 -0.966652
+ 8.53e+10Hz 0.0446431 -0.966677
+ 8.54e+10Hz 0.0429315 -0.966698
+ 8.55e+10Hz 0.0412205 -0.966716
+ 8.56e+10Hz 0.03951 -0.966731
+ 8.57e+10Hz 0.0378001 -0.966743
+ 8.58e+10Hz 0.0360907 -0.966752
+ 8.59e+10Hz 0.034382 -0.966758
+ 8.6e+10Hz 0.0326738 -0.96676
+ 8.61e+10Hz 0.0309663 -0.96676
+ 8.62e+10Hz 0.0292594 -0.966756
+ 8.63e+10Hz 0.0275531 -0.966749
+ 8.64e+10Hz 0.0258474 -0.966739
+ 8.65e+10Hz 0.0241424 -0.966727
+ 8.66e+10Hz 0.022438 -0.966711
+ 8.67e+10Hz 0.0207343 -0.966692
+ 8.68e+10Hz 0.0190312 -0.96667
+ 8.69e+10Hz 0.0173288 -0.966645
+ 8.7e+10Hz 0.015627 -0.966617
+ 8.71e+10Hz 0.0139259 -0.966586
+ 8.72e+10Hz 0.0122255 -0.966552
+ 8.73e+10Hz 0.0105258 -0.966515
+ 8.74e+10Hz 0.00882669 -0.966476
+ 8.75e+10Hz 0.0071283 -0.966433
+ 8.76e+10Hz 0.0054306 -0.966388
+ 8.77e+10Hz 0.00373359 -0.966339
+ 8.78e+10Hz 0.00203726 -0.966288
+ 8.79e+10Hz 0.00034163 -0.966233
+ 8.8e+10Hz -0.00135331 -0.966176
+ 8.81e+10Hz -0.00304755 -0.966116
+ 8.82e+10Hz -0.0047411 -0.966054
+ 8.83e+10Hz -0.00643395 -0.965988
+ 8.84e+10Hz -0.00812611 -0.96592
+ 8.85e+10Hz -0.00981757 -0.965848
+ 8.86e+10Hz -0.0115083 -0.965774
+ 8.87e+10Hz -0.0131984 -0.965698
+ 8.88e+10Hz -0.0148877 -0.965618
+ 8.89e+10Hz -0.0165764 -0.965536
+ 8.9e+10Hz -0.0182644 -0.965451
+ 8.91e+10Hz -0.0199517 -0.965363
+ 8.92e+10Hz -0.0216382 -0.965272
+ 8.93e+10Hz -0.0233241 -0.965179
+ 8.94e+10Hz -0.0250093 -0.965083
+ 8.95e+10Hz -0.0266938 -0.964984
+ 8.96e+10Hz -0.0283776 -0.964883
+ 8.97e+10Hz -0.0300607 -0.964778
+ 8.98e+10Hz -0.0317432 -0.964672
+ 8.99e+10Hz -0.0334249 -0.964562
+ 9e+10Hz -0.035106 -0.96445
+ 9.01e+10Hz -0.0367864 -0.964335
+ 9.02e+10Hz -0.0384661 -0.964217
+ 9.03e+10Hz -0.0401451 -0.964097
+ 9.04e+10Hz -0.0418235 -0.963975
+ 9.05e+10Hz -0.0435011 -0.963849
+ 9.06e+10Hz -0.0451782 -0.963721
+ 9.07e+10Hz -0.0468545 -0.96359
+ 9.08e+10Hz -0.0485302 -0.963457
+ 9.09e+10Hz -0.0502052 -0.963321
+ 9.1e+10Hz -0.0518795 -0.963183
+ 9.11e+10Hz -0.0535532 -0.963041
+ 9.12e+10Hz -0.0552262 -0.962898
+ 9.13e+10Hz -0.0568986 -0.962751
+ 9.14e+10Hz -0.0585703 -0.962602
+ 9.15e+10Hz -0.0602414 -0.962451
+ 9.16e+10Hz -0.0619118 -0.962297
+ 9.17e+10Hz -0.0635815 -0.96214
+ 9.18e+10Hz -0.0652506 -0.961981
+ 9.19e+10Hz -0.0669191 -0.961819
+ 9.2e+10Hz -0.0685869 -0.961655
+ 9.21e+10Hz -0.0702541 -0.961488
+ 9.22e+10Hz -0.0719206 -0.961318
+ 9.23e+10Hz -0.0735865 -0.961146
+ 9.24e+10Hz -0.0752518 -0.960971
+ 9.25e+10Hz -0.0769164 -0.960794
+ 9.26e+10Hz -0.0785804 -0.960615
+ 9.27e+10Hz -0.0802437 -0.960432
+ 9.28e+10Hz -0.0819064 -0.960247
+ 9.29e+10Hz -0.0835685 -0.96006
+ 9.3e+10Hz -0.0852299 -0.95987
+ 9.31e+10Hz -0.0868907 -0.959678
+ 9.32e+10Hz -0.0885509 -0.959483
+ 9.33e+10Hz -0.0902104 -0.959285
+ 9.34e+10Hz -0.0918693 -0.959085
+ 9.35e+10Hz -0.0935276 -0.958883
+ 9.36e+10Hz -0.0951853 -0.958678
+ 9.37e+10Hz -0.0968423 -0.95847
+ 9.38e+10Hz -0.0984986 -0.95826
+ 9.39e+10Hz -0.100154 -0.958047
+ 9.4e+10Hz -0.10181 -0.957832
+ 9.41e+10Hz -0.103464 -0.957614
+ 9.42e+10Hz -0.105118 -0.957394
+ 9.43e+10Hz -0.106771 -0.957172
+ 9.44e+10Hz -0.108424 -0.956946
+ 9.45e+10Hz -0.110076 -0.956719
+ 9.46e+10Hz -0.111727 -0.956488
+ 9.47e+10Hz -0.113377 -0.956256
+ 9.48e+10Hz -0.115028 -0.95602
+ 9.49e+10Hz -0.116677 -0.955783
+ 9.5e+10Hz -0.118326 -0.955542
+ 9.51e+10Hz -0.119974 -0.9553
+ 9.52e+10Hz -0.121621 -0.955055
+ 9.53e+10Hz -0.123268 -0.954807
+ 9.54e+10Hz -0.124914 -0.954557
+ 9.55e+10Hz -0.12656 -0.954304
+ 9.56e+10Hz -0.128205 -0.954049
+ 9.57e+10Hz -0.129849 -0.953791
+ 9.58e+10Hz -0.131492 -0.953531
+ 9.59e+10Hz -0.133135 -0.953269
+ 9.6e+10Hz -0.134777 -0.953004
+ 9.61e+10Hz -0.136419 -0.952736
+ 9.62e+10Hz -0.13806 -0.952466
+ 9.63e+10Hz -0.1397 -0.952194
+ 9.64e+10Hz -0.14134 -0.951919
+ 9.65e+10Hz -0.142979 -0.951642
+ 9.66e+10Hz -0.144617 -0.951362
+ 9.67e+10Hz -0.146255 -0.95108
+ 9.68e+10Hz -0.147892 -0.950795
+ 9.69e+10Hz -0.149528 -0.950508
+ 9.7e+10Hz -0.151164 -0.950219
+ 9.71e+10Hz -0.152799 -0.949927
+ 9.72e+10Hz -0.154433 -0.949633
+ 9.73e+10Hz -0.156067 -0.949336
+ 9.74e+10Hz -0.1577 -0.949037
+ 9.75e+10Hz -0.159332 -0.948735
+ 9.76e+10Hz -0.160964 -0.948431
+ 9.77e+10Hz -0.162595 -0.948125
+ 9.78e+10Hz -0.164225 -0.947816
+ 9.79e+10Hz -0.165855 -0.947505
+ 9.8e+10Hz -0.167484 -0.947191
+ 9.81e+10Hz -0.169112 -0.946875
+ 9.82e+10Hz -0.17074 -0.946557
+ 9.83e+10Hz -0.172367 -0.946236
+ 9.84e+10Hz -0.173993 -0.945913
+ 9.85e+10Hz -0.175619 -0.945588
+ 9.86e+10Hz -0.177244 -0.94526
+ 9.87e+10Hz -0.178868 -0.94493
+ 9.88e+10Hz -0.180492 -0.944598
+ 9.89e+10Hz -0.182115 -0.944263
+ 9.9e+10Hz -0.183737 -0.943926
+ 9.91e+10Hz -0.185359 -0.943586
+ 9.92e+10Hz -0.18698 -0.943244
+ 9.93e+10Hz -0.1886 -0.9429
+ 9.94e+10Hz -0.19022 -0.942554
+ 9.95e+10Hz -0.191839 -0.942205
+ 9.96e+10Hz -0.193458 -0.941854
+ 9.97e+10Hz -0.195076 -0.941501
+ 9.98e+10Hz -0.196693 -0.941145
+ 9.99e+10Hz -0.19831 -0.940787
+ 1e+11Hz -0.199926 -0.940427
+ 1.001e+11Hz -0.201541 -0.940064
+ 1.002e+11Hz -0.203156 -0.939699
+ 1.003e+11Hz -0.20477 -0.939332
+ 1.004e+11Hz -0.206384 -0.938962
+ 1.005e+11Hz -0.207997 -0.938591
+ 1.006e+11Hz -0.209609 -0.938217
+ 1.007e+11Hz -0.211221 -0.93784
+ 1.008e+11Hz -0.212832 -0.937462
+ 1.009e+11Hz -0.214443 -0.937081
+ 1.01e+11Hz -0.216053 -0.936698
+ 1.011e+11Hz -0.217662 -0.936312
+ 1.012e+11Hz -0.219271 -0.935925
+ 1.013e+11Hz -0.22088 -0.935535
+ 1.014e+11Hz -0.222488 -0.935143
+ 1.015e+11Hz -0.224095 -0.934748
+ 1.016e+11Hz -0.225702 -0.934351
+ 1.017e+11Hz -0.227308 -0.933952
+ 1.018e+11Hz -0.228914 -0.933551
+ 1.019e+11Hz -0.230519 -0.933148
+ 1.02e+11Hz -0.232124 -0.932742
+ 1.021e+11Hz -0.233728 -0.932334
+ 1.022e+11Hz -0.235332 -0.931924
+ 1.023e+11Hz -0.236935 -0.931511
+ 1.024e+11Hz -0.238538 -0.931096
+ 1.025e+11Hz -0.24014 -0.930679
+ 1.026e+11Hz -0.241742 -0.93026
+ 1.027e+11Hz -0.243343 -0.929838
+ 1.028e+11Hz -0.244944 -0.929414
+ 1.029e+11Hz -0.246545 -0.928988
+ 1.03e+11Hz -0.248145 -0.928559
+ 1.031e+11Hz -0.249744 -0.928128
+ 1.032e+11Hz -0.251343 -0.927695
+ 1.033e+11Hz -0.252942 -0.92726
+ 1.034e+11Hz -0.254541 -0.926822
+ 1.035e+11Hz -0.256138 -0.926382
+ 1.036e+11Hz -0.257736 -0.925939
+ 1.037e+11Hz -0.259333 -0.925495
+ 1.038e+11Hz -0.26093 -0.925048
+ 1.039e+11Hz -0.262526 -0.924598
+ 1.04e+11Hz -0.264122 -0.924146
+ 1.041e+11Hz -0.265718 -0.923692
+ 1.042e+11Hz -0.267313 -0.923236
+ 1.043e+11Hz -0.268908 -0.922777
+ 1.044e+11Hz -0.270503 -0.922316
+ 1.045e+11Hz -0.272097 -0.921852
+ 1.046e+11Hz -0.273691 -0.921386
+ 1.047e+11Hz -0.275285 -0.920918
+ 1.048e+11Hz -0.276878 -0.920447
+ 1.049e+11Hz -0.278471 -0.919974
+ 1.05e+11Hz -0.280064 -0.919498
+ 1.051e+11Hz -0.281656 -0.91902
+ 1.052e+11Hz -0.283248 -0.918539
+ 1.053e+11Hz -0.28484 -0.918056
+ 1.054e+11Hz -0.286431 -0.917571
+ 1.055e+11Hz -0.288022 -0.917083
+ 1.056e+11Hz -0.289613 -0.916592
+ 1.057e+11Hz -0.291203 -0.916099
+ 1.058e+11Hz -0.292793 -0.915604
+ 1.059e+11Hz -0.294383 -0.915106
+ 1.06e+11Hz -0.295973 -0.914605
+ 1.061e+11Hz -0.297562 -0.914102
+ 1.062e+11Hz -0.299151 -0.913596
+ 1.063e+11Hz -0.30074 -0.913088
+ 1.064e+11Hz -0.302328 -0.912577
+ 1.065e+11Hz -0.303916 -0.912063
+ 1.066e+11Hz -0.305504 -0.911547
+ 1.067e+11Hz -0.307091 -0.911028
+ 1.068e+11Hz -0.308678 -0.910507
+ 1.069e+11Hz -0.310265 -0.909983
+ 1.07e+11Hz -0.311852 -0.909456
+ 1.071e+11Hz -0.313438 -0.908926
+ 1.072e+11Hz -0.315024 -0.908394
+ 1.073e+11Hz -0.31661 -0.907859
+ 1.074e+11Hz -0.318195 -0.907321
+ 1.075e+11Hz -0.31978 -0.906781
+ 1.076e+11Hz -0.321364 -0.906238
+ 1.077e+11Hz -0.322948 -0.905692
+ 1.078e+11Hz -0.324532 -0.905143
+ 1.079e+11Hz -0.326116 -0.904591
+ 1.08e+11Hz -0.327699 -0.904037
+ 1.081e+11Hz -0.329282 -0.90348
+ 1.082e+11Hz -0.330864 -0.90292
+ 1.083e+11Hz -0.332446 -0.902357
+ 1.084e+11Hz -0.334028 -0.901791
+ 1.085e+11Hz -0.335609 -0.901222
+ 1.086e+11Hz -0.33719 -0.900651
+ 1.087e+11Hz -0.33877 -0.900076
+ 1.088e+11Hz -0.34035 -0.899499
+ 1.089e+11Hz -0.34193 -0.898919
+ 1.09e+11Hz -0.343509 -0.898335
+ 1.091e+11Hz -0.345087 -0.897749
+ 1.092e+11Hz -0.346665 -0.89716
+ 1.093e+11Hz -0.348243 -0.896568
+ 1.094e+11Hz -0.34982 -0.895972
+ 1.095e+11Hz -0.351396 -0.895374
+ 1.096e+11Hz -0.352972 -0.894773
+ 1.097e+11Hz -0.354548 -0.894169
+ 1.098e+11Hz -0.356123 -0.893561
+ 1.099e+11Hz -0.357697 -0.892951
+ 1.1e+11Hz -0.359271 -0.892338
+ 1.101e+11Hz -0.360844 -0.891721
+ 1.102e+11Hz -0.362416 -0.891102
+ 1.103e+11Hz -0.363988 -0.890479
+ 1.104e+11Hz -0.365559 -0.889854
+ 1.105e+11Hz -0.36713 -0.889225
+ 1.106e+11Hz -0.368699 -0.888593
+ 1.107e+11Hz -0.370268 -0.887958
+ 1.108e+11Hz -0.371837 -0.88732
+ 1.109e+11Hz -0.373404 -0.886679
+ 1.11e+11Hz -0.374971 -0.886034
+ 1.111e+11Hz -0.376537 -0.885387
+ 1.112e+11Hz -0.378103 -0.884736
+ 1.113e+11Hz -0.379667 -0.884082
+ 1.114e+11Hz -0.381231 -0.883425
+ 1.115e+11Hz -0.382794 -0.882765
+ 1.116e+11Hz -0.384356 -0.882102
+ 1.117e+11Hz -0.385917 -0.881436
+ 1.118e+11Hz -0.387477 -0.880766
+ 1.119e+11Hz -0.389036 -0.880093
+ 1.12e+11Hz -0.390594 -0.879418
+ 1.121e+11Hz -0.392152 -0.878739
+ 1.122e+11Hz -0.393708 -0.878056
+ 1.123e+11Hz -0.395264 -0.877371
+ 1.124e+11Hz -0.396818 -0.876682
+ 1.125e+11Hz -0.398371 -0.875991
+ 1.126e+11Hz -0.399924 -0.875296
+ 1.127e+11Hz -0.401475 -0.874598
+ 1.128e+11Hz -0.403025 -0.873897
+ 1.129e+11Hz -0.404574 -0.873192
+ 1.13e+11Hz -0.406122 -0.872485
+ 1.131e+11Hz -0.407669 -0.871774
+ 1.132e+11Hz -0.409215 -0.87106
+ 1.133e+11Hz -0.410759 -0.870343
+ 1.134e+11Hz -0.412302 -0.869623
+ 1.135e+11Hz -0.413845 -0.8689
+ 1.136e+11Hz -0.415385 -0.868174
+ 1.137e+11Hz -0.416925 -0.867444
+ 1.138e+11Hz -0.418463 -0.866711
+ 1.139e+11Hz -0.420001 -0.865976
+ 1.14e+11Hz -0.421536 -0.865237
+ 1.141e+11Hz -0.423071 -0.864495
+ 1.142e+11Hz -0.424604 -0.86375
+ 1.143e+11Hz -0.426136 -0.863002
+ 1.144e+11Hz -0.427666 -0.862251
+ 1.145e+11Hz -0.429195 -0.861496
+ 1.146e+11Hz -0.430723 -0.860739
+ 1.147e+11Hz -0.432249 -0.859979
+ 1.148e+11Hz -0.433774 -0.859215
+ 1.149e+11Hz -0.435298 -0.858449
+ 1.15e+11Hz -0.43682 -0.857679
+ 1.151e+11Hz -0.438341 -0.856907
+ 1.152e+11Hz -0.43986 -0.856131
+ 1.153e+11Hz -0.441377 -0.855352
+ 1.154e+11Hz -0.442893 -0.854571
+ 1.155e+11Hz -0.444408 -0.853786
+ 1.156e+11Hz -0.445921 -0.852999
+ 1.157e+11Hz -0.447433 -0.852209
+ 1.158e+11Hz -0.448943 -0.851415
+ 1.159e+11Hz -0.450451 -0.850619
+ 1.16e+11Hz -0.451958 -0.84982
+ 1.161e+11Hz -0.453464 -0.849018
+ 1.162e+11Hz -0.454967 -0.848213
+ 1.163e+11Hz -0.45647 -0.847405
+ 1.164e+11Hz -0.45797 -0.846594
+ 1.165e+11Hz -0.459469 -0.84578
+ 1.166e+11Hz -0.460967 -0.844964
+ 1.167e+11Hz -0.462462 -0.844144
+ 1.168e+11Hz -0.463957 -0.843322
+ 1.169e+11Hz -0.465449 -0.842497
+ 1.17e+11Hz -0.46694 -0.841669
+ 1.171e+11Hz -0.468429 -0.840839
+ 1.172e+11Hz -0.469917 -0.840005
+ 1.173e+11Hz -0.471402 -0.839169
+ 1.174e+11Hz -0.472887 -0.83833
+ 1.175e+11Hz -0.474369 -0.837488
+ 1.176e+11Hz -0.47585 -0.836644
+ 1.177e+11Hz -0.477329 -0.835797
+ 1.178e+11Hz -0.478807 -0.834947
+ 1.179e+11Hz -0.480282 -0.834094
+ 1.18e+11Hz -0.481757 -0.833239
+ 1.181e+11Hz -0.483229 -0.832381
+ 1.182e+11Hz -0.4847 -0.83152
+ 1.183e+11Hz -0.486169 -0.830657
+ 1.184e+11Hz -0.487636 -0.829791
+ 1.185e+11Hz -0.489101 -0.828923
+ 1.186e+11Hz -0.490565 -0.828051
+ 1.187e+11Hz -0.492027 -0.827177
+ 1.188e+11Hz -0.493488 -0.826301
+ 1.189e+11Hz -0.494947 -0.825422
+ 1.19e+11Hz -0.496404 -0.82454
+ 1.191e+11Hz -0.497859 -0.823656
+ 1.192e+11Hz -0.499312 -0.822769
+ 1.193e+11Hz -0.500764 -0.82188
+ 1.194e+11Hz -0.502214 -0.820988
+ 1.195e+11Hz -0.503663 -0.820093
+ 1.196e+11Hz -0.50511 -0.819196
+ 1.197e+11Hz -0.506554 -0.818296
+ 1.198e+11Hz -0.507998 -0.817394
+ 1.199e+11Hz -0.509439 -0.81649
+ 1.2e+11Hz -0.510879 -0.815582
+ 1.201e+11Hz -0.512317 -0.814673
+ 1.202e+11Hz -0.513754 -0.81376
+ 1.203e+11Hz -0.515188 -0.812846
+ 1.204e+11Hz -0.516621 -0.811928
+ 1.205e+11Hz -0.518052 -0.811009
+ 1.206e+11Hz -0.519482 -0.810086
+ 1.207e+11Hz -0.52091 -0.809162
+ 1.208e+11Hz -0.522336 -0.808235
+ 1.209e+11Hz -0.52376 -0.807305
+ 1.21e+11Hz -0.525183 -0.806373
+ 1.211e+11Hz -0.526604 -0.805438
+ 1.212e+11Hz -0.528023 -0.804501
+ 1.213e+11Hz -0.52944 -0.803562
+ 1.214e+11Hz -0.530856 -0.80262
+ 1.215e+11Hz -0.53227 -0.801675
+ 1.216e+11Hz -0.533683 -0.800728
+ 1.217e+11Hz -0.535093 -0.799779
+ 1.218e+11Hz -0.536502 -0.798827
+ 1.219e+11Hz -0.53791 -0.797873
+ 1.22e+11Hz -0.539315 -0.796917
+ 1.221e+11Hz -0.540719 -0.795958
+ 1.222e+11Hz -0.542121 -0.794996
+ 1.223e+11Hz -0.543522 -0.794032
+ 1.224e+11Hz -0.54492 -0.793066
+ 1.225e+11Hz -0.546317 -0.792097
+ 1.226e+11Hz -0.547713 -0.791125
+ 1.227e+11Hz -0.549106 -0.790152
+ 1.228e+11Hz -0.550498 -0.789176
+ 1.229e+11Hz -0.551888 -0.788197
+ 1.23e+11Hz -0.553277 -0.787216
+ 1.231e+11Hz -0.554664 -0.786233
+ 1.232e+11Hz -0.556049 -0.785247
+ 1.233e+11Hz -0.557432 -0.784258
+ 1.234e+11Hz -0.558813 -0.783267
+ 1.235e+11Hz -0.560193 -0.782274
+ 1.236e+11Hz -0.561571 -0.781279
+ 1.237e+11Hz -0.562948 -0.78028
+ 1.238e+11Hz -0.564322 -0.77928
+ 1.239e+11Hz -0.565695 -0.778277
+ 1.24e+11Hz -0.567066 -0.777271
+ 1.241e+11Hz -0.568436 -0.776264
+ 1.242e+11Hz -0.569803 -0.775253
+ 1.243e+11Hz -0.571169 -0.77424
+ 1.244e+11Hz -0.572533 -0.773225
+ 1.245e+11Hz -0.573896 -0.772208
+ 1.246e+11Hz -0.575256 -0.771187
+ 1.247e+11Hz -0.576615 -0.770165
+ 1.248e+11Hz -0.577972 -0.76914
+ 1.249e+11Hz -0.579327 -0.768112
+ 1.25e+11Hz -0.580681 -0.767082
+ 1.251e+11Hz -0.582032 -0.76605
+ 1.252e+11Hz -0.583382 -0.765015
+ 1.253e+11Hz -0.58473 -0.763978
+ 1.254e+11Hz -0.586076 -0.762938
+ 1.255e+11Hz -0.587421 -0.761896
+ 1.256e+11Hz -0.588763 -0.760851
+ 1.257e+11Hz -0.590104 -0.759804
+ 1.258e+11Hz -0.591443 -0.758754
+ 1.259e+11Hz -0.59278 -0.757702
+ 1.26e+11Hz -0.594115 -0.756648
+ 1.261e+11Hz -0.595448 -0.755591
+ 1.262e+11Hz -0.596779 -0.754531
+ 1.263e+11Hz -0.598109 -0.753469
+ 1.264e+11Hz -0.599436 -0.752405
+ 1.265e+11Hz -0.600762 -0.751338
+ 1.266e+11Hz -0.602086 -0.750269
+ 1.267e+11Hz -0.603407 -0.749197
+ 1.268e+11Hz -0.604727 -0.748123
+ 1.269e+11Hz -0.606045 -0.747047
+ 1.27e+11Hz -0.607361 -0.745968
+ 1.271e+11Hz -0.608675 -0.744886
+ 1.272e+11Hz -0.609987 -0.743802
+ 1.273e+11Hz -0.611297 -0.742716
+ 1.274e+11Hz -0.612605 -0.741627
+ 1.275e+11Hz -0.613911 -0.740536
+ 1.276e+11Hz -0.615215 -0.739442
+ 1.277e+11Hz -0.616517 -0.738346
+ 1.278e+11Hz -0.617817 -0.737248
+ 1.279e+11Hz -0.619115 -0.736147
+ 1.28e+11Hz -0.62041 -0.735044
+ 1.281e+11Hz -0.621704 -0.733938
+ 1.282e+11Hz -0.622996 -0.73283
+ 1.283e+11Hz -0.624285 -0.73172
+ 1.284e+11Hz -0.625573 -0.730607
+ 1.285e+11Hz -0.626858 -0.729492
+ 1.286e+11Hz -0.628141 -0.728375
+ 1.287e+11Hz -0.629422 -0.727255
+ 1.288e+11Hz -0.630701 -0.726133
+ 1.289e+11Hz -0.631978 -0.725008
+ 1.29e+11Hz -0.633253 -0.723881
+ 1.291e+11Hz -0.634525 -0.722752
+ 1.292e+11Hz -0.635795 -0.721621
+ 1.293e+11Hz -0.637064 -0.720487
+ 1.294e+11Hz -0.63833 -0.719351
+ 1.295e+11Hz -0.639593 -0.718212
+ 1.296e+11Hz -0.640855 -0.717072
+ 1.297e+11Hz -0.642114 -0.715929
+ 1.298e+11Hz -0.643371 -0.714783
+ 1.299e+11Hz -0.644626 -0.713636
+ 1.3e+11Hz -0.645879 -0.712486
+ 1.301e+11Hz -0.647129 -0.711334
+ 1.302e+11Hz -0.648377 -0.71018
+ 1.303e+11Hz -0.649623 -0.709024
+ 1.304e+11Hz -0.650866 -0.707865
+ 1.305e+11Hz -0.652108 -0.706704
+ 1.306e+11Hz -0.653347 -0.705541
+ 1.307e+11Hz -0.654583 -0.704376
+ 1.308e+11Hz -0.655818 -0.703209
+ 1.309e+11Hz -0.65705 -0.70204
+ 1.31e+11Hz -0.65828 -0.700868
+ 1.311e+11Hz -0.659507 -0.699695
+ 1.312e+11Hz -0.660732 -0.698519
+ 1.313e+11Hz -0.661955 -0.697341
+ 1.314e+11Hz -0.663176 -0.696161
+ 1.315e+11Hz -0.664394 -0.694979
+ 1.316e+11Hz -0.66561 -0.693795
+ 1.317e+11Hz -0.666823 -0.692609
+ 1.318e+11Hz -0.668034 -0.691421
+ 1.319e+11Hz -0.669243 -0.690231
+ 1.32e+11Hz -0.670449 -0.689039
+ 1.321e+11Hz -0.671654 -0.687844
+ 1.322e+11Hz -0.672855 -0.686648
+ 1.323e+11Hz -0.674055 -0.68545
+ 1.324e+11Hz -0.675252 -0.68425
+ 1.325e+11Hz -0.676447 -0.683048
+ 1.326e+11Hz -0.677639 -0.681844
+ 1.327e+11Hz -0.678829 -0.680639
+ 1.328e+11Hz -0.680017 -0.679431
+ 1.329e+11Hz -0.681202 -0.678221
+ 1.33e+11Hz -0.682385 -0.67701
+ 1.331e+11Hz -0.683566 -0.675796
+ 1.332e+11Hz -0.684744 -0.674581
+ 1.333e+11Hz -0.68592 -0.673364
+ 1.334e+11Hz -0.687093 -0.672145
+ 1.335e+11Hz -0.688264 -0.670925
+ 1.336e+11Hz -0.689433 -0.669702
+ 1.337e+11Hz -0.6906 -0.668478
+ 1.338e+11Hz -0.691764 -0.667252
+ 1.339e+11Hz -0.692926 -0.666024
+ 1.34e+11Hz -0.694085 -0.664794
+ 1.341e+11Hz -0.695243 -0.663563
+ 1.342e+11Hz -0.696398 -0.66233
+ 1.343e+11Hz -0.69755 -0.661095
+ 1.344e+11Hz -0.6987 -0.659858
+ 1.345e+11Hz -0.699848 -0.65862
+ 1.346e+11Hz -0.700994 -0.65738
+ 1.347e+11Hz -0.702137 -0.656138
+ 1.348e+11Hz -0.703278 -0.654895
+ 1.349e+11Hz -0.704417 -0.65365
+ 1.35e+11Hz -0.705554 -0.652403
+ 1.351e+11Hz -0.706688 -0.651155
+ 1.352e+11Hz -0.70782 -0.649905
+ 1.353e+11Hz -0.70895 -0.648653
+ 1.354e+11Hz -0.710077 -0.6474
+ 1.355e+11Hz -0.711202 -0.646145
+ 1.356e+11Hz -0.712325 -0.644888
+ 1.357e+11Hz -0.713446 -0.64363
+ 1.358e+11Hz -0.714564 -0.642371
+ 1.359e+11Hz -0.715681 -0.641109
+ 1.36e+11Hz -0.716795 -0.639846
+ 1.361e+11Hz -0.717907 -0.638582
+ 1.362e+11Hz -0.719016 -0.637316
+ 1.363e+11Hz -0.720124 -0.636048
+ 1.364e+11Hz -0.721229 -0.634779
+ 1.365e+11Hz -0.722332 -0.633508
+ 1.366e+11Hz -0.723433 -0.632235
+ 1.367e+11Hz -0.724532 -0.630962
+ 1.368e+11Hz -0.725628 -0.629686
+ 1.369e+11Hz -0.726723 -0.628409
+ 1.37e+11Hz -0.727815 -0.62713
+ 1.371e+11Hz -0.728905 -0.62585
+ 1.372e+11Hz -0.729994 -0.624569
+ 1.373e+11Hz -0.731079 -0.623285
+ 1.374e+11Hz -0.732163 -0.622
+ 1.375e+11Hz -0.733245 -0.620714
+ 1.376e+11Hz -0.734325 -0.619426
+ 1.377e+11Hz -0.735402 -0.618137
+ 1.378e+11Hz -0.736478 -0.616846
+ 1.379e+11Hz -0.737551 -0.615553
+ 1.38e+11Hz -0.738623 -0.614259
+ 1.381e+11Hz -0.739692 -0.612964
+ 1.382e+11Hz -0.740759 -0.611667
+ 1.383e+11Hz -0.741825 -0.610368
+ 1.384e+11Hz -0.742888 -0.609068
+ 1.385e+11Hz -0.743949 -0.607766
+ 1.386e+11Hz -0.745008 -0.606463
+ 1.387e+11Hz -0.746065 -0.605158
+ 1.388e+11Hz -0.74712 -0.603851
+ 1.389e+11Hz -0.748174 -0.602543
+ 1.39e+11Hz -0.749225 -0.601234
+ 1.391e+11Hz -0.750274 -0.599923
+ 1.392e+11Hz -0.751321 -0.59861
+ 1.393e+11Hz -0.752366 -0.597296
+ 1.394e+11Hz -0.753409 -0.59598
+ 1.395e+11Hz -0.754451 -0.594663
+ 1.396e+11Hz -0.75549 -0.593344
+ 1.397e+11Hz -0.756527 -0.592023
+ 1.398e+11Hz -0.757562 -0.590701
+ 1.399e+11Hz -0.758596 -0.589377
+ 1.4e+11Hz -0.759627 -0.588052
+ 1.401e+11Hz -0.760657 -0.586725
+ 1.402e+11Hz -0.761684 -0.585396
+ 1.403e+11Hz -0.76271 -0.584066
+ 1.404e+11Hz -0.763733 -0.582735
+ 1.405e+11Hz -0.764755 -0.581401
+ 1.406e+11Hz -0.765775 -0.580066
+ 1.407e+11Hz -0.766792 -0.578729
+ 1.408e+11Hz -0.767808 -0.577391
+ 1.409e+11Hz -0.768822 -0.576051
+ 1.41e+11Hz -0.769834 -0.574709
+ 1.411e+11Hz -0.770844 -0.573366
+ 1.412e+11Hz -0.771852 -0.572021
+ 1.413e+11Hz -0.772858 -0.570674
+ 1.414e+11Hz -0.773863 -0.569326
+ 1.415e+11Hz -0.774865 -0.567976
+ 1.416e+11Hz -0.775865 -0.566624
+ 1.417e+11Hz -0.776864 -0.565271
+ 1.418e+11Hz -0.77786 -0.563916
+ 1.419e+11Hz -0.778855 -0.562559
+ 1.42e+11Hz -0.779848 -0.561201
+ 1.421e+11Hz -0.780838 -0.55984
+ 1.422e+11Hz -0.781827 -0.558478
+ 1.423e+11Hz -0.782814 -0.557115
+ 1.424e+11Hz -0.783799 -0.555749
+ 1.425e+11Hz -0.784782 -0.554382
+ 1.426e+11Hz -0.785762 -0.553013
+ 1.427e+11Hz -0.786741 -0.551642
+ 1.428e+11Hz -0.787718 -0.550269
+ 1.429e+11Hz -0.788694 -0.548895
+ 1.43e+11Hz -0.789667 -0.547519
+ 1.431e+11Hz -0.790638 -0.546141
+ 1.432e+11Hz -0.791607 -0.544762
+ 1.433e+11Hz -0.792574 -0.54338
+ 1.434e+11Hz -0.793539 -0.541997
+ 1.435e+11Hz -0.794502 -0.540612
+ 1.436e+11Hz -0.795463 -0.539225
+ 1.437e+11Hz -0.796423 -0.537836
+ 1.438e+11Hz -0.79738 -0.536446
+ 1.439e+11Hz -0.798335 -0.535053
+ 1.44e+11Hz -0.799288 -0.533659
+ 1.441e+11Hz -0.800239 -0.532263
+ 1.442e+11Hz -0.801188 -0.530865
+ 1.443e+11Hz -0.802135 -0.529465
+ 1.444e+11Hz -0.80308 -0.528064
+ 1.445e+11Hz -0.804023 -0.52666
+ 1.446e+11Hz -0.804964 -0.525255
+ 1.447e+11Hz -0.805903 -0.523848
+ 1.448e+11Hz -0.806839 -0.522439
+ 1.449e+11Hz -0.807774 -0.521028
+ 1.45e+11Hz -0.808706 -0.519615
+ 1.451e+11Hz -0.809637 -0.5182
+ 1.452e+11Hz -0.810565 -0.516784
+ 1.453e+11Hz -0.811491 -0.515365
+ 1.454e+11Hz -0.812415 -0.513945
+ 1.455e+11Hz -0.813337 -0.512522
+ 1.456e+11Hz -0.814257 -0.511098
+ 1.457e+11Hz -0.815175 -0.509672
+ 1.458e+11Hz -0.81609 -0.508244
+ 1.459e+11Hz -0.817003 -0.506814
+ 1.46e+11Hz -0.817914 -0.505383
+ 1.461e+11Hz -0.818823 -0.503949
+ 1.462e+11Hz -0.81973 -0.502514
+ 1.463e+11Hz -0.820635 -0.501076
+ 1.464e+11Hz -0.821537 -0.499637
+ 1.465e+11Hz -0.822437 -0.498195
+ 1.466e+11Hz -0.823335 -0.496752
+ 1.467e+11Hz -0.824231 -0.495307
+ 1.468e+11Hz -0.825124 -0.49386
+ 1.469e+11Hz -0.826015 -0.492411
+ 1.47e+11Hz -0.826904 -0.49096
+ 1.471e+11Hz -0.827791 -0.489507
+ 1.472e+11Hz -0.828675 -0.488052
+ 1.473e+11Hz -0.829557 -0.486596
+ 1.474e+11Hz -0.830437 -0.485137
+ 1.475e+11Hz -0.831314 -0.483677
+ 1.476e+11Hz -0.83219 -0.482214
+ 1.477e+11Hz -0.833062 -0.48075
+ 1.478e+11Hz -0.833933 -0.479284
+ 1.479e+11Hz -0.834801 -0.477816
+ 1.48e+11Hz -0.835667 -0.476346
+ 1.481e+11Hz -0.83653 -0.474874
+ 1.482e+11Hz -0.837391 -0.4734
+ 1.483e+11Hz -0.83825 -0.471924
+ 1.484e+11Hz -0.839106 -0.470446
+ 1.485e+11Hz -0.83996 -0.468967
+ 1.486e+11Hz -0.840811 -0.467485
+ 1.487e+11Hz -0.84166 -0.466002
+ 1.488e+11Hz -0.842507 -0.464516
+ 1.489e+11Hz -0.843351 -0.463029
+ 1.49e+11Hz -0.844193 -0.46154
+ 1.491e+11Hz -0.845032 -0.460049
+ 1.492e+11Hz -0.845869 -0.458556
+ 1.493e+11Hz -0.846703 -0.457061
+ 1.494e+11Hz -0.847535 -0.455564
+ 1.495e+11Hz -0.848364 -0.454065
+ 1.496e+11Hz -0.849191 -0.452565
+ 1.497e+11Hz -0.850015 -0.451062
+ 1.498e+11Hz -0.850837 -0.449558
+ 1.499e+11Hz -0.851656 -0.448052
+ 1.5e+11Hz -0.852473 -0.446544
+ 1.501e+11Hz -0.853287 -0.445034
+ 1.502e+11Hz -0.854099 -0.443522
+ 1.503e+11Hz -0.854908 -0.442008
+ 1.504e+11Hz -0.855715 -0.440492
+ 1.505e+11Hz -0.856518 -0.438975
+ 1.506e+11Hz -0.85732 -0.437456
+ 1.507e+11Hz -0.858118 -0.435934
+ 1.508e+11Hz -0.858915 -0.434411
+ 1.509e+11Hz -0.859708 -0.432886
+ 1.51e+11Hz -0.860499 -0.431359
+ 1.511e+11Hz -0.861287 -0.429831
+ 1.512e+11Hz -0.862073 -0.4283
+ 1.513e+11Hz -0.862856 -0.426768
+ 1.514e+11Hz -0.863636 -0.425234
+ 1.515e+11Hz -0.864413 -0.423698
+ 1.516e+11Hz -0.865188 -0.42216
+ 1.517e+11Hz -0.865961 -0.42062
+ 1.518e+11Hz -0.86673 -0.419079
+ 1.519e+11Hz -0.867497 -0.417535
+ 1.52e+11Hz -0.868261 -0.41599
+ 1.521e+11Hz -0.869022 -0.414443
+ 1.522e+11Hz -0.869781 -0.412894
+ 1.523e+11Hz -0.870537 -0.411344
+ 1.524e+11Hz -0.87129 -0.409791
+ 1.525e+11Hz -0.87204 -0.408237
+ 1.526e+11Hz -0.872788 -0.406681
+ 1.527e+11Hz -0.873532 -0.405123
+ 1.528e+11Hz -0.874274 -0.403563
+ 1.529e+11Hz -0.875013 -0.402002
+ 1.53e+11Hz -0.87575 -0.400439
+ 1.531e+11Hz -0.876483 -0.398874
+ 1.532e+11Hz -0.877214 -0.397307
+ 1.533e+11Hz -0.877942 -0.395739
+ 1.534e+11Hz -0.878667 -0.394168
+ 1.535e+11Hz -0.879389 -0.392596
+ 1.536e+11Hz -0.880108 -0.391022
+ 1.537e+11Hz -0.880824 -0.389447
+ 1.538e+11Hz -0.881538 -0.38787
+ 1.539e+11Hz -0.882248 -0.386291
+ 1.54e+11Hz -0.882956 -0.38471
+ 1.541e+11Hz -0.883661 -0.383127
+ 1.542e+11Hz -0.884362 -0.381543
+ 1.543e+11Hz -0.885061 -0.379957
+ 1.544e+11Hz -0.885757 -0.378369
+ 1.545e+11Hz -0.88645 -0.37678
+ 1.546e+11Hz -0.88714 -0.375189
+ 1.547e+11Hz -0.887827 -0.373596
+ 1.548e+11Hz -0.888511 -0.372002
+ 1.549e+11Hz -0.889192 -0.370406
+ 1.55e+11Hz -0.88987 -0.368808
+ 1.551e+11Hz -0.890544 -0.367208
+ 1.552e+11Hz -0.891216 -0.365607
+ 1.553e+11Hz -0.891885 -0.364004
+ 1.554e+11Hz -0.892551 -0.3624
+ 1.555e+11Hz -0.893213 -0.360794
+ 1.556e+11Hz -0.893873 -0.359186
+ 1.557e+11Hz -0.894529 -0.357577
+ 1.558e+11Hz -0.895183 -0.355966
+ 1.559e+11Hz -0.895833 -0.354353
+ 1.56e+11Hz -0.89648 -0.352739
+ 1.561e+11Hz -0.897124 -0.351123
+ 1.562e+11Hz -0.897765 -0.349506
+ 1.563e+11Hz -0.898403 -0.347887
+ 1.564e+11Hz -0.899037 -0.346267
+ 1.565e+11Hz -0.899669 -0.344645
+ 1.566e+11Hz -0.900297 -0.343021
+ 1.567e+11Hz -0.900922 -0.341396
+ 1.568e+11Hz -0.901543 -0.339769
+ 1.569e+11Hz -0.902162 -0.338141
+ 1.57e+11Hz -0.902777 -0.336511
+ 1.571e+11Hz -0.903389 -0.33488
+ 1.572e+11Hz -0.903998 -0.333247
+ 1.573e+11Hz -0.904604 -0.331613
+ 1.574e+11Hz -0.905206 -0.329978
+ 1.575e+11Hz -0.905805 -0.328341
+ 1.576e+11Hz -0.906401 -0.326702
+ 1.577e+11Hz -0.906993 -0.325062
+ 1.578e+11Hz -0.907582 -0.323421
+ 1.579e+11Hz -0.908168 -0.321778
+ 1.58e+11Hz -0.90875 -0.320134
+ 1.581e+11Hz -0.90933 -0.318488
+ 1.582e+11Hz -0.909905 -0.316841
+ 1.583e+11Hz -0.910478 -0.315193
+ 1.584e+11Hz -0.911047 -0.313543
+ 1.585e+11Hz -0.911613 -0.311892
+ 1.586e+11Hz -0.912175 -0.31024
+ 1.587e+11Hz -0.912734 -0.308586
+ 1.588e+11Hz -0.913289 -0.306931
+ 1.589e+11Hz -0.913841 -0.305275
+ 1.59e+11Hz -0.91439 -0.303618
+ 1.591e+11Hz -0.914935 -0.301959
+ 1.592e+11Hz -0.915477 -0.300299
+ 1.593e+11Hz -0.916016 -0.298638
+ 1.594e+11Hz -0.916551 -0.296975
+ 1.595e+11Hz -0.917082 -0.295312
+ 1.596e+11Hz -0.91761 -0.293647
+ 1.597e+11Hz -0.918135 -0.291981
+ 1.598e+11Hz -0.918656 -0.290314
+ 1.599e+11Hz -0.919173 -0.288645
+ 1.6e+11Hz -0.919688 -0.286976
+ 1.601e+11Hz -0.920198 -0.285305
+ 1.602e+11Hz -0.920705 -0.283634
+ 1.603e+11Hz -0.921209 -0.281961
+ 1.604e+11Hz -0.921709 -0.280287
+ 1.605e+11Hz -0.922206 -0.278613
+ 1.606e+11Hz -0.922699 -0.276937
+ 1.607e+11Hz -0.923189 -0.27526
+ 1.608e+11Hz -0.923675 -0.273582
+ 1.609e+11Hz -0.924157 -0.271903
+ 1.61e+11Hz -0.924636 -0.270223
+ 1.611e+11Hz -0.925112 -0.268543
+ 1.612e+11Hz -0.925584 -0.266861
+ 1.613e+11Hz -0.926052 -0.265178
+ 1.614e+11Hz -0.926517 -0.263495
+ 1.615e+11Hz -0.926979 -0.26181
+ 1.616e+11Hz -0.927436 -0.260125
+ 1.617e+11Hz -0.927891 -0.258439
+ 1.618e+11Hz -0.928341 -0.256752
+ 1.619e+11Hz -0.928788 -0.255064
+ 1.62e+11Hz -0.929232 -0.253376
+ 1.621e+11Hz -0.929672 -0.251686
+ 1.622e+11Hz -0.930109 -0.249996
+ 1.623e+11Hz -0.930542 -0.248305
+ 1.624e+11Hz -0.930971 -0.246613
+ 1.625e+11Hz -0.931397 -0.244921
+ 1.626e+11Hz -0.931819 -0.243228
+ 1.627e+11Hz -0.932238 -0.241534
+ 1.628e+11Hz -0.932653 -0.23984
+ 1.629e+11Hz -0.933065 -0.238145
+ 1.63e+11Hz -0.933473 -0.236449
+ 1.631e+11Hz -0.933877 -0.234752
+ 1.632e+11Hz -0.934278 -0.233055
+ 1.633e+11Hz -0.934676 -0.231358
+ 1.634e+11Hz -0.93507 -0.229659
+ 1.635e+11Hz -0.93546 -0.22796
+ 1.636e+11Hz -0.935847 -0.226261
+ 1.637e+11Hz -0.93623 -0.224561
+ 1.638e+11Hz -0.93661 -0.222861
+ 1.639e+11Hz -0.936986 -0.22116
+ 1.64e+11Hz -0.937359 -0.219458
+ 1.641e+11Hz -0.937728 -0.217756
+ 1.642e+11Hz -0.938094 -0.216054
+ 1.643e+11Hz -0.938456 -0.214351
+ 1.644e+11Hz -0.938815 -0.212648
+ 1.645e+11Hz -0.93917 -0.210944
+ 1.646e+11Hz -0.939522 -0.20924
+ 1.647e+11Hz -0.93987 -0.207535
+ 1.648e+11Hz -0.940215 -0.20583
+ 1.649e+11Hz -0.940557 -0.204125
+ 1.65e+11Hz -0.940894 -0.202419
+ 1.651e+11Hz -0.941229 -0.200713
+ 1.652e+11Hz -0.94156 -0.199006
+ 1.653e+11Hz -0.941887 -0.1973
+ 1.654e+11Hz -0.942211 -0.195593
+ 1.655e+11Hz -0.942532 -0.193885
+ 1.656e+11Hz -0.942849 -0.192177
+ 1.657e+11Hz -0.943163 -0.190469
+ 1.658e+11Hz -0.943473 -0.188761
+ 1.659e+11Hz -0.94378 -0.187053
+ 1.66e+11Hz -0.944084 -0.185344
+ 1.661e+11Hz -0.944384 -0.183635
+ 1.662e+11Hz -0.94468 -0.181925
+ 1.663e+11Hz -0.944974 -0.180216
+ 1.664e+11Hz -0.945264 -0.178506
+ 1.665e+11Hz -0.94555 -0.176796
+ 1.666e+11Hz -0.945834 -0.175086
+ 1.667e+11Hz -0.946113 -0.173376
+ 1.668e+11Hz -0.94639 -0.171665
+ 1.669e+11Hz -0.946663 -0.169954
+ 1.67e+11Hz -0.946933 -0.168244
+ 1.671e+11Hz -0.947199 -0.166532
+ 1.672e+11Hz -0.947463 -0.164821
+ 1.673e+11Hz -0.947722 -0.16311
+ 1.674e+11Hz -0.947979 -0.161398
+ 1.675e+11Hz -0.948232 -0.159687
+ 1.676e+11Hz -0.948482 -0.157975
+ 1.677e+11Hz -0.948729 -0.156263
+ 1.678e+11Hz -0.948972 -0.154551
+ 1.679e+11Hz -0.949212 -0.152839
+ 1.68e+11Hz -0.949449 -0.151127
+ 1.681e+11Hz -0.949683 -0.149414
+ 1.682e+11Hz -0.949913 -0.147702
+ 1.683e+11Hz -0.95014 -0.145989
+ 1.684e+11Hz -0.950364 -0.144277
+ 1.685e+11Hz -0.950584 -0.142564
+ 1.686e+11Hz -0.950802 -0.140851
+ 1.687e+11Hz -0.951016 -0.139138
+ 1.688e+11Hz -0.951227 -0.137425
+ 1.689e+11Hz -0.951434 -0.135712
+ 1.69e+11Hz -0.951639 -0.133999
+ 1.691e+11Hz -0.95184 -0.132286
+ 1.692e+11Hz -0.952038 -0.130573
+ 1.693e+11Hz -0.952233 -0.12886
+ 1.694e+11Hz -0.952424 -0.127147
+ 1.695e+11Hz -0.952613 -0.125433
+ 1.696e+11Hz -0.952798 -0.12372
+ 1.697e+11Hz -0.95298 -0.122007
+ 1.698e+11Hz -0.953159 -0.120293
+ 1.699e+11Hz -0.953335 -0.11858
+ 1.7e+11Hz -0.953507 -0.116866
+ 1.701e+11Hz -0.953677 -0.115153
+ 1.702e+11Hz -0.953843 -0.113439
+ 1.703e+11Hz -0.954006 -0.111726
+ 1.704e+11Hz -0.954166 -0.110012
+ 1.705e+11Hz -0.954323 -0.108299
+ 1.706e+11Hz -0.954476 -0.106585
+ 1.707e+11Hz -0.954627 -0.104871
+ 1.708e+11Hz -0.954774 -0.103158
+ 1.709e+11Hz -0.954918 -0.101444
+ 1.71e+11Hz -0.955059 -0.0997304
+ 1.711e+11Hz -0.955197 -0.0980167
+ 1.712e+11Hz -0.955332 -0.0963031
+ 1.713e+11Hz -0.955463 -0.0945894
+ 1.714e+11Hz -0.955592 -0.0928758
+ 1.715e+11Hz -0.955717 -0.0911621
+ 1.716e+11Hz -0.955839 -0.0894485
+ 1.717e+11Hz -0.955958 -0.0877349
+ 1.718e+11Hz -0.956074 -0.0860213
+ 1.719e+11Hz -0.956187 -0.0843077
+ 1.72e+11Hz -0.956297 -0.0825942
+ 1.721e+11Hz -0.956403 -0.0808806
+ 1.722e+11Hz -0.956506 -0.0791671
+ 1.723e+11Hz -0.956607 -0.0774537
+ 1.724e+11Hz -0.956704 -0.0757402
+ 1.725e+11Hz -0.956798 -0.0740268
+ 1.726e+11Hz -0.956888 -0.0723134
+ 1.727e+11Hz -0.956976 -0.0706001
+ 1.728e+11Hz -0.957061 -0.0688868
+ 1.729e+11Hz -0.957142 -0.0671736
+ 1.73e+11Hz -0.95722 -0.0654604
+ 1.731e+11Hz -0.957295 -0.0637473
+ 1.732e+11Hz -0.957367 -0.0620342
+ 1.733e+11Hz -0.957436 -0.0603212
+ 1.734e+11Hz -0.957502 -0.0586083
+ 1.735e+11Hz -0.957564 -0.0568954
+ 1.736e+11Hz -0.957623 -0.0551826
+ 1.737e+11Hz -0.95768 -0.0534699
+ 1.738e+11Hz -0.957733 -0.0517573
+ 1.739e+11Hz -0.957783 -0.0500448
+ 1.74e+11Hz -0.957829 -0.0483324
+ 1.741e+11Hz -0.957873 -0.0466201
+ 1.742e+11Hz -0.957913 -0.0449079
+ 1.743e+11Hz -0.95795 -0.0431958
+ 1.744e+11Hz -0.957985 -0.0414839
+ 1.745e+11Hz -0.958015 -0.039772
+ 1.746e+11Hz -0.958043 -0.0380603
+ 1.747e+11Hz -0.958068 -0.0363488
+ 1.748e+11Hz -0.958089 -0.0346373
+ 1.749e+11Hz -0.958107 -0.0329261
+ 1.75e+11Hz -0.958122 -0.031215
+ 1.751e+11Hz -0.958134 -0.029504
+ 1.752e+11Hz -0.958143 -0.0277932
+ 1.753e+11Hz -0.958148 -0.0260826
+ 1.754e+11Hz -0.958151 -0.0243722
+ 1.755e+11Hz -0.95815 -0.022662
+ 1.756e+11Hz -0.958146 -0.020952
+ 1.757e+11Hz -0.958139 -0.0192422
+ 1.758e+11Hz -0.958128 -0.0175326
+ 1.759e+11Hz -0.958114 -0.0158233
+ 1.76e+11Hz -0.958098 -0.0141142
+ 1.761e+11Hz -0.958078 -0.0124053
+ 1.762e+11Hz -0.958054 -0.0106967
+ 1.763e+11Hz -0.958028 -0.00898832
+ 1.764e+11Hz -0.957998 -0.00728022
+ 1.765e+11Hz -0.957965 -0.0055724
+ 1.766e+11Hz -0.957929 -0.00386487
+ 1.767e+11Hz -0.95789 -0.00215764
+ 1.768e+11Hz -0.957848 -0.00045071
+ 1.769e+11Hz -0.957802 0.00125591
+ 1.77e+11Hz -0.957753 0.0029622
+ 1.771e+11Hz -0.957701 0.00466815
+ 1.772e+11Hz -0.957646 0.00637377
+ 1.773e+11Hz -0.957587 0.00807903
+ 1.774e+11Hz -0.957526 0.00978393
+ 1.775e+11Hz -0.957461 0.0114885
+ 1.776e+11Hz -0.957393 0.0131926
+ 1.777e+11Hz -0.957322 0.0148964
+ 1.778e+11Hz -0.957247 0.0165997
+ 1.779e+11Hz -0.957169 0.0183026
+ 1.78e+11Hz -0.957089 0.0200052
+ 1.781e+11Hz -0.957004 0.0217072
+ 1.782e+11Hz -0.956917 0.0234089
+ 1.783e+11Hz -0.956827 0.0251101
+ 1.784e+11Hz -0.956733 0.0268108
+ 1.785e+11Hz -0.956636 0.028511
+ 1.786e+11Hz -0.956536 0.0302108
+ 1.787e+11Hz -0.956433 0.0319101
+ 1.788e+11Hz -0.956326 0.0336088
+ 1.789e+11Hz -0.956217 0.0353071
+ 1.79e+11Hz -0.956104 0.0370048
+ 1.791e+11Hz -0.955988 0.038702
+ 1.792e+11Hz -0.955869 0.0403986
+ 1.793e+11Hz -0.955747 0.0420947
+ 1.794e+11Hz -0.955621 0.0437902
+ 1.795e+11Hz -0.955493 0.0454851
+ 1.796e+11Hz -0.955361 0.0471795
+ 1.797e+11Hz -0.955226 0.0488732
+ 1.798e+11Hz -0.955088 0.0505664
+ 1.799e+11Hz -0.954947 0.0522589
+ 1.8e+11Hz -0.954802 0.0539508
+ 1.801e+11Hz -0.954655 0.055642
+ 1.802e+11Hz -0.954504 0.0573326
+ 1.803e+11Hz -0.95435 0.0590226
+ 1.804e+11Hz -0.954193 0.0607119
+ 1.805e+11Hz -0.954033 0.0624005
+ 1.806e+11Hz -0.95387 0.0640884
+ 1.807e+11Hz -0.953704 0.0657756
+ 1.808e+11Hz -0.953534 0.0674621
+ 1.809e+11Hz -0.953362 0.0691479
+ 1.81e+11Hz -0.953186 0.070833
+ 1.811e+11Hz -0.953008 0.0725173
+ 1.812e+11Hz -0.952826 0.0742009
+ 1.813e+11Hz -0.952641 0.0758837
+ 1.814e+11Hz -0.952453 0.0775658
+ 1.815e+11Hz -0.952262 0.0792471
+ 1.816e+11Hz -0.952068 0.0809276
+ 1.817e+11Hz -0.951871 0.0826073
+ 1.818e+11Hz -0.951671 0.0842863
+ 1.819e+11Hz -0.951468 0.0859644
+ 1.82e+11Hz -0.951262 0.0876417
+ 1.821e+11Hz -0.951053 0.0893182
+ 1.822e+11Hz -0.95084 0.0909938
+ 1.823e+11Hz -0.950625 0.0926687
+ 1.824e+11Hz -0.950407 0.0943426
+ 1.825e+11Hz -0.950186 0.0960158
+ 1.826e+11Hz -0.949961 0.097688
+ 1.827e+11Hz -0.949734 0.0993594
+ 1.828e+11Hz -0.949504 0.10103
+ 1.829e+11Hz -0.949271 0.1027
+ 1.83e+11Hz -0.949035 0.104368
+ 1.831e+11Hz -0.948796 0.106036
+ 1.832e+11Hz -0.948553 0.107703
+ 1.833e+11Hz -0.948308 0.109369
+ 1.834e+11Hz -0.948061 0.111034
+ 1.835e+11Hz -0.94781 0.112698
+ 1.836e+11Hz -0.947556 0.114362
+ 1.837e+11Hz -0.947299 0.116024
+ 1.838e+11Hz -0.94704 0.117685
+ 1.839e+11Hz -0.946777 0.119346
+ 1.84e+11Hz -0.946512 0.121005
+ 1.841e+11Hz -0.946244 0.122663
+ 1.842e+11Hz -0.945972 0.124321
+ 1.843e+11Hz -0.945698 0.125977
+ 1.844e+11Hz -0.945422 0.127633
+ 1.845e+11Hz -0.945142 0.129288
+ 1.846e+11Hz -0.944859 0.130941
+ 1.847e+11Hz -0.944574 0.132594
+ 1.848e+11Hz -0.944286 0.134245
+ 1.849e+11Hz -0.943995 0.135896
+ 1.85e+11Hz -0.943701 0.137545
+ 1.851e+11Hz -0.943404 0.139194
+ 1.852e+11Hz -0.943105 0.140841
+ 1.853e+11Hz -0.942802 0.142488
+ 1.854e+11Hz -0.942497 0.144133
+ 1.855e+11Hz -0.942189 0.145777
+ 1.856e+11Hz -0.941879 0.147421
+ 1.857e+11Hz -0.941565 0.149063
+ 1.858e+11Hz -0.941249 0.150704
+ 1.859e+11Hz -0.940931 0.152344
+ 1.86e+11Hz -0.940609 0.153983
+ 1.861e+11Hz -0.940285 0.155621
+ 1.862e+11Hz -0.939958 0.157258
+ 1.863e+11Hz -0.939628 0.158894
+ 1.864e+11Hz -0.939295 0.160529
+ 1.865e+11Hz -0.93896 0.162162
+ 1.866e+11Hz -0.938622 0.163795
+ 1.867e+11Hz -0.938282 0.165426
+ 1.868e+11Hz -0.937938 0.167056
+ 1.869e+11Hz -0.937593 0.168686
+ 1.87e+11Hz -0.937244 0.170314
+ 1.871e+11Hz -0.936893 0.171941
+ 1.872e+11Hz -0.936539 0.173567
+ 1.873e+11Hz -0.936182 0.175191
+ 1.874e+11Hz -0.935823 0.176815
+ 1.875e+11Hz -0.935462 0.178437
+ 1.876e+11Hz -0.935097 0.180059
+ 1.877e+11Hz -0.93473 0.181679
+ 1.878e+11Hz -0.934361 0.183298
+ 1.879e+11Hz -0.933989 0.184916
+ 1.88e+11Hz -0.933614 0.186532
+ 1.881e+11Hz -0.933237 0.188148
+ 1.882e+11Hz -0.932857 0.189762
+ 1.883e+11Hz -0.932474 0.191375
+ 1.884e+11Hz -0.932089 0.192987
+ 1.885e+11Hz -0.931702 0.194598
+ 1.886e+11Hz -0.931312 0.196208
+ 1.887e+11Hz -0.930919 0.197816
+ 1.888e+11Hz -0.930524 0.199424
+ 1.889e+11Hz -0.930127 0.20103
+ 1.89e+11Hz -0.929727 0.202635
+ 1.891e+11Hz -0.929324 0.204238
+ 1.892e+11Hz -0.928919 0.205841
+ 1.893e+11Hz -0.928512 0.207442
+ 1.894e+11Hz -0.928102 0.209042
+ 1.895e+11Hz -0.927689 0.210641
+ 1.896e+11Hz -0.927274 0.212239
+ 1.897e+11Hz -0.926857 0.213835
+ 1.898e+11Hz -0.926438 0.21543
+ 1.899e+11Hz -0.926016 0.217024
+ 1.9e+11Hz -0.925591 0.218617
+ 1.901e+11Hz -0.925164 0.220209
+ 1.902e+11Hz -0.924735 0.221799
+ 1.903e+11Hz -0.924303 0.223388
+ 1.904e+11Hz -0.92387 0.224976
+ 1.905e+11Hz -0.923433 0.226562
+ 1.906e+11Hz -0.922995 0.228148
+ 1.907e+11Hz -0.922554 0.229732
+ 1.908e+11Hz -0.92211 0.231315
+ 1.909e+11Hz -0.921665 0.232896
+ 1.91e+11Hz -0.921217 0.234477
+ 1.911e+11Hz -0.920767 0.236056
+ 1.912e+11Hz -0.920315 0.237634
+ 1.913e+11Hz -0.91986 0.23921
+ 1.914e+11Hz -0.919403 0.240786
+ 1.915e+11Hz -0.918944 0.24236
+ 1.916e+11Hz -0.918483 0.243933
+ 1.917e+11Hz -0.918019 0.245504
+ 1.918e+11Hz -0.917553 0.247075
+ 1.919e+11Hz -0.917085 0.248644
+ 1.92e+11Hz -0.916615 0.250212
+ 1.921e+11Hz -0.916143 0.251779
+ 1.922e+11Hz -0.915669 0.253344
+ 1.923e+11Hz -0.915192 0.254908
+ 1.924e+11Hz -0.914713 0.256471
+ 1.925e+11Hz -0.914233 0.258033
+ 1.926e+11Hz -0.91375 0.259593
+ 1.927e+11Hz -0.913265 0.261153
+ 1.928e+11Hz -0.912778 0.262711
+ 1.929e+11Hz -0.912289 0.264267
+ 1.93e+11Hz -0.911797 0.265823
+ 1.931e+11Hz -0.911304 0.267377
+ 1.932e+11Hz -0.910809 0.26893
+ 1.933e+11Hz -0.910312 0.270482
+ 1.934e+11Hz -0.909813 0.272033
+ 1.935e+11Hz -0.909311 0.273583
+ 1.936e+11Hz -0.908808 0.275131
+ 1.937e+11Hz -0.908303 0.276678
+ 1.938e+11Hz -0.907796 0.278224
+ 1.939e+11Hz -0.907287 0.279769
+ 1.94e+11Hz -0.906776 0.281313
+ 1.941e+11Hz -0.906263 0.282855
+ 1.942e+11Hz -0.905748 0.284396
+ 1.943e+11Hz -0.905231 0.285937
+ 1.944e+11Hz -0.904712 0.287476
+ 1.945e+11Hz -0.904192 0.289014
+ 1.946e+11Hz -0.90367 0.29055
+ 1.947e+11Hz -0.903145 0.292086
+ 1.948e+11Hz -0.902619 0.293621
+ 1.949e+11Hz -0.902091 0.295154
+ 1.95e+11Hz -0.901562 0.296687
+ 1.951e+11Hz -0.90103 0.298218
+ 1.952e+11Hz -0.900497 0.299749
+ 1.953e+11Hz -0.899962 0.301278
+ 1.954e+11Hz -0.899425 0.302806
+ 1.955e+11Hz -0.898886 0.304333
+ 1.956e+11Hz -0.898346 0.30586
+ 1.957e+11Hz -0.897804 0.307385
+ 1.958e+11Hz -0.89726 0.308909
+ 1.959e+11Hz -0.896714 0.310432
+ 1.96e+11Hz -0.896167 0.311955
+ 1.961e+11Hz -0.895617 0.313476
+ 1.962e+11Hz -0.895067 0.314997
+ 1.963e+11Hz -0.894514 0.316516
+ 1.964e+11Hz -0.89396 0.318035
+ 1.965e+11Hz -0.893404 0.319553
+ 1.966e+11Hz -0.892846 0.32107
+ 1.967e+11Hz -0.892287 0.322586
+ 1.968e+11Hz -0.891726 0.324101
+ 1.969e+11Hz -0.891163 0.325615
+ 1.97e+11Hz -0.890599 0.327129
+ 1.971e+11Hz -0.890033 0.328642
+ 1.972e+11Hz -0.889465 0.330154
+ 1.973e+11Hz -0.888896 0.331665
+ 1.974e+11Hz -0.888324 0.333176
+ 1.975e+11Hz -0.887752 0.334686
+ 1.976e+11Hz -0.887177 0.336195
+ 1.977e+11Hz -0.886601 0.337704
+ 1.978e+11Hz -0.886024 0.339211
+ 1.979e+11Hz -0.885444 0.340719
+ 1.98e+11Hz -0.884863 0.342225
+ 1.981e+11Hz -0.88428 0.343731
+ 1.982e+11Hz -0.883696 0.345237
+ 1.983e+11Hz -0.88311 0.346741
+ 1.984e+11Hz -0.882522 0.348246
+ 1.985e+11Hz -0.881933 0.34975
+ 1.986e+11Hz -0.881342 0.351253
+ 1.987e+11Hz -0.880749 0.352755
+ 1.988e+11Hz -0.880154 0.354258
+ 1.989e+11Hz -0.879558 0.35576
+ 1.99e+11Hz -0.87896 0.357261
+ 1.991e+11Hz -0.878361 0.358762
+ 1.992e+11Hz -0.877759 0.360262
+ 1.993e+11Hz -0.877156 0.361763
+ 1.994e+11Hz -0.876551 0.363262
+ 1.995e+11Hz -0.875945 0.364762
+ 1.996e+11Hz -0.875336 0.366261
+ 1.997e+11Hz -0.874726 0.36776
+ 1.998e+11Hz -0.874114 0.369258
+ 1.999e+11Hz -0.8735 0.370756
+ 2e+11Hz -0.872885 0.372254
+ 2.001e+11Hz -0.872267 0.373752
+ 2.002e+11Hz -0.871648 0.37525
+ 2.003e+11Hz -0.871027 0.376747
+ 2.004e+11Hz -0.870404 0.378244
+ 2.005e+11Hz -0.869779 0.379741
+ 2.006e+11Hz -0.869152 0.381238
+ 2.007e+11Hz -0.868524 0.382734
+ 2.008e+11Hz -0.867893 0.384231
+ 2.009e+11Hz -0.86726 0.385727
+ 2.01e+11Hz -0.866626 0.387223
+ 2.011e+11Hz -0.865989 0.388719
+ 2.012e+11Hz -0.86535 0.390215
+ 2.013e+11Hz -0.86471 0.391711
+ 2.014e+11Hz -0.864067 0.393207
+ 2.015e+11Hz -0.863422 0.394703
+ 2.016e+11Hz -0.862775 0.396198
+ 2.017e+11Hz -0.862126 0.397694
+ 2.018e+11Hz -0.861475 0.39919
+ 2.019e+11Hz -0.860822 0.400686
+ 2.02e+11Hz -0.860166 0.402181
+ 2.021e+11Hz -0.859508 0.403677
+ 2.022e+11Hz -0.858848 0.405173
+ 2.023e+11Hz -0.858186 0.406668
+ 2.024e+11Hz -0.857522 0.408164
+ 2.025e+11Hz -0.856855 0.40966
+ 2.026e+11Hz -0.856185 0.411156
+ 2.027e+11Hz -0.855514 0.412652
+ 2.028e+11Hz -0.85484 0.414148
+ 2.029e+11Hz -0.854163 0.415644
+ 2.03e+11Hz -0.853485 0.41714
+ 2.031e+11Hz -0.852803 0.418636
+ 2.032e+11Hz -0.852119 0.420132
+ 2.033e+11Hz -0.851433 0.421628
+ 2.034e+11Hz -0.850744 0.423124
+ 2.035e+11Hz -0.850053 0.42462
+ 2.036e+11Hz -0.849358 0.426116
+ 2.037e+11Hz -0.848662 0.427613
+ 2.038e+11Hz -0.847962 0.429109
+ 2.039e+11Hz -0.84726 0.430606
+ 2.04e+11Hz -0.846555 0.432102
+ 2.041e+11Hz -0.845847 0.433598
+ 2.042e+11Hz -0.845137 0.435095
+ 2.043e+11Hz -0.844424 0.436591
+ 2.044e+11Hz -0.843708 0.438088
+ 2.045e+11Hz -0.842989 0.439584
+ 2.046e+11Hz -0.842267 0.44108
+ 2.047e+11Hz -0.841542 0.442577
+ 2.048e+11Hz -0.840815 0.444073
+ 2.049e+11Hz -0.840084 0.445569
+ 2.05e+11Hz -0.83935 0.447065
+ 2.051e+11Hz -0.838614 0.448561
+ 2.052e+11Hz -0.837874 0.450057
+ 2.053e+11Hz -0.837131 0.451553
+ 2.054e+11Hz -0.836385 0.453049
+ 2.055e+11Hz -0.835636 0.454545
+ 2.056e+11Hz -0.834884 0.45604
+ 2.057e+11Hz -0.834129 0.457535
+ 2.058e+11Hz -0.83337 0.45903
+ 2.059e+11Hz -0.832608 0.460525
+ 2.06e+11Hz -0.831843 0.462019
+ 2.061e+11Hz -0.831075 0.463514
+ 2.062e+11Hz -0.830303 0.465008
+ 2.063e+11Hz -0.829528 0.466501
+ 2.064e+11Hz -0.82875 0.467995
+ 2.065e+11Hz -0.827968 0.469488
+ 2.066e+11Hz -0.827183 0.47098
+ 2.067e+11Hz -0.826394 0.472472
+ 2.068e+11Hz -0.825602 0.473964
+ 2.069e+11Hz -0.824807 0.475456
+ 2.07e+11Hz -0.824008 0.476946
+ 2.071e+11Hz -0.823206 0.478437
+ 2.072e+11Hz -0.8224 0.479926
+ 2.073e+11Hz -0.821591 0.481416
+ 2.074e+11Hz -0.820778 0.482904
+ 2.075e+11Hz -0.819961 0.484392
+ 2.076e+11Hz -0.819141 0.48588
+ 2.077e+11Hz -0.818318 0.487366
+ 2.078e+11Hz -0.81749 0.488852
+ 2.079e+11Hz -0.81666 0.490337
+ 2.08e+11Hz -0.815825 0.491822
+ 2.081e+11Hz -0.814987 0.493306
+ 2.082e+11Hz -0.814146 0.494788
+ 2.083e+11Hz -0.8133 0.49627
+ 2.084e+11Hz -0.812451 0.497751
+ 2.085e+11Hz -0.811599 0.499231
+ 2.086e+11Hz -0.810742 0.500711
+ 2.087e+11Hz -0.809882 0.502189
+ 2.088e+11Hz -0.809019 0.503666
+ 2.089e+11Hz -0.808151 0.505142
+ 2.09e+11Hz -0.80728 0.506617
+ 2.091e+11Hz -0.806405 0.508091
+ 2.092e+11Hz -0.805527 0.509564
+ 2.093e+11Hz -0.804645 0.511035
+ 2.094e+11Hz -0.803759 0.512505
+ 2.095e+11Hz -0.802869 0.513974
+ 2.096e+11Hz -0.801976 0.515442
+ 2.097e+11Hz -0.801079 0.516909
+ 2.098e+11Hz -0.800178 0.518374
+ 2.099e+11Hz -0.799274 0.519837
+ 2.1e+11Hz -0.798365 0.5213
+ 2.101e+11Hz -0.797454 0.522761
+ 2.102e+11Hz -0.796538 0.52422
+ 2.103e+11Hz -0.795619 0.525678
+ 2.104e+11Hz -0.794696 0.527134
+ 2.105e+11Hz -0.79377 0.528589
+ 2.106e+11Hz -0.792839 0.530042
+ 2.107e+11Hz -0.791905 0.531493
+ 2.108e+11Hz -0.790968 0.532943
+ 2.109e+11Hz -0.790027 0.534391
+ 2.11e+11Hz -0.789082 0.535838
+ 2.111e+11Hz -0.788134 0.537282
+ 2.112e+11Hz -0.787182 0.538725
+ 2.113e+11Hz -0.786226 0.540166
+ 2.114e+11Hz -0.785267 0.541605
+ 2.115e+11Hz -0.784304 0.543043
+ 2.116e+11Hz -0.783338 0.544478
+ 2.117e+11Hz -0.782368 0.545912
+ 2.118e+11Hz -0.781395 0.547343
+ 2.119e+11Hz -0.780418 0.548773
+ 2.12e+11Hz -0.779438 0.5502
+ 2.121e+11Hz -0.778454 0.551626
+ 2.122e+11Hz -0.777467 0.553049
+ 2.123e+11Hz -0.776476 0.554471
+ 2.124e+11Hz -0.775482 0.55589
+ 2.125e+11Hz -0.774484 0.557307
+ 2.126e+11Hz -0.773484 0.558722
+ 2.127e+11Hz -0.772479 0.560135
+ 2.128e+11Hz -0.771472 0.561545
+ 2.129e+11Hz -0.770461 0.562954
+ 2.13e+11Hz -0.769446 0.56436
+ 2.131e+11Hz -0.768429 0.565764
+ 2.132e+11Hz -0.767408 0.567166
+ 2.133e+11Hz -0.766384 0.568565
+ 2.134e+11Hz -0.765357 0.569962
+ 2.135e+11Hz -0.764326 0.571357
+ 2.136e+11Hz -0.763293 0.57275
+ 2.137e+11Hz -0.762256 0.57414
+ 2.138e+11Hz -0.761216 0.575528
+ 2.139e+11Hz -0.760173 0.576913
+ 2.14e+11Hz -0.759127 0.578296
+ 2.141e+11Hz -0.758078 0.579677
+ 2.142e+11Hz -0.757025 0.581055
+ 2.143e+11Hz -0.75597 0.58243
+ 2.144e+11Hz -0.754912 0.583804
+ 2.145e+11Hz -0.753851 0.585175
+ 2.146e+11Hz -0.752786 0.586543
+ 2.147e+11Hz -0.751719 0.587909
+ 2.148e+11Hz -0.750649 0.589272
+ 2.149e+11Hz -0.749576 0.590633
+ 2.15e+11Hz -0.7485 0.591992
+ 2.151e+11Hz -0.747421 0.593348
+ 2.152e+11Hz -0.74634 0.594701
+ 2.153e+11Hz -0.745255 0.596052
+ 2.154e+11Hz -0.744168 0.597401
+ 2.155e+11Hz -0.743078 0.598746
+ 2.156e+11Hz -0.741985 0.60009
+ 2.157e+11Hz -0.74089 0.601431
+ 2.158e+11Hz -0.739792 0.602769
+ 2.159e+11Hz -0.738691 0.604105
+ 2.16e+11Hz -0.737587 0.605438
+ 2.161e+11Hz -0.736481 0.606769
+ 2.162e+11Hz -0.735372 0.608097
+ 2.163e+11Hz -0.734261 0.609422
+ 2.164e+11Hz -0.733147 0.610745
+ 2.165e+11Hz -0.73203 0.612066
+ 2.166e+11Hz -0.730911 0.613384
+ 2.167e+11Hz -0.729789 0.614699
+ 2.168e+11Hz -0.728665 0.616012
+ 2.169e+11Hz -0.727538 0.617322
+ 2.17e+11Hz -0.726409 0.61863
+ 2.171e+11Hz -0.725277 0.619935
+ 2.172e+11Hz -0.724142 0.621238
+ 2.173e+11Hz -0.723006 0.622538
+ 2.174e+11Hz -0.721866 0.623836
+ 2.175e+11Hz -0.720725 0.625131
+ 2.176e+11Hz -0.719581 0.626424
+ 2.177e+11Hz -0.718434 0.627714
+ 2.178e+11Hz -0.717285 0.629001
+ 2.179e+11Hz -0.716134 0.630286
+ 2.18e+11Hz -0.714981 0.631569
+ 2.181e+11Hz -0.713825 0.632848
+ 2.182e+11Hz -0.712666 0.634126
+ 2.183e+11Hz -0.711506 0.635401
+ 2.184e+11Hz -0.710343 0.636673
+ 2.185e+11Hz -0.709177 0.637943
+ 2.186e+11Hz -0.70801 0.639211
+ 2.187e+11Hz -0.70684 0.640475
+ 2.188e+11Hz -0.705667 0.641738
+ 2.189e+11Hz -0.704493 0.642998
+ 2.19e+11Hz -0.703316 0.644255
+ 2.191e+11Hz -0.702137 0.64551
+ 2.192e+11Hz -0.700956 0.646763
+ 2.193e+11Hz -0.699772 0.648012
+ 2.194e+11Hz -0.698586 0.64926
+ 2.195e+11Hz -0.697398 0.650505
+ 2.196e+11Hz -0.696207 0.651747
+ 2.197e+11Hz -0.695015 0.652988
+ 2.198e+11Hz -0.69382 0.654225
+ 2.199e+11Hz -0.692623 0.65546
+ 2.2e+11Hz -0.691423 0.656693
+ 2.201e+11Hz -0.690222 0.657923
+ 2.202e+11Hz -0.689018 0.659151
+ 2.203e+11Hz -0.687812 0.660376
+ 2.204e+11Hz -0.686604 0.661599
+ 2.205e+11Hz -0.685393 0.662819
+ 2.206e+11Hz -0.684181 0.664037
+ 2.207e+11Hz -0.682966 0.665252
+ 2.208e+11Hz -0.681749 0.666465
+ 2.209e+11Hz -0.680529 0.667676
+ 2.21e+11Hz -0.679308 0.668884
+ 2.211e+11Hz -0.678084 0.670089
+ 2.212e+11Hz -0.676858 0.671292
+ 2.213e+11Hz -0.67563 0.672492
+ 2.214e+11Hz -0.674399 0.673691
+ 2.215e+11Hz -0.673167 0.674886
+ 2.216e+11Hz -0.671932 0.676079
+ 2.217e+11Hz -0.670695 0.67727
+ 2.218e+11Hz -0.669456 0.678458
+ 2.219e+11Hz -0.668215 0.679643
+ 2.22e+11Hz -0.666971 0.680826
+ 2.221e+11Hz -0.665725 0.682007
+ 2.222e+11Hz -0.664477 0.683185
+ 2.223e+11Hz -0.663227 0.68436
+ 2.224e+11Hz -0.661975 0.685533
+ 2.225e+11Hz -0.66072 0.686704
+ 2.226e+11Hz -0.659463 0.687871
+ 2.227e+11Hz -0.658204 0.689037
+ 2.228e+11Hz -0.656943 0.690199
+ 2.229e+11Hz -0.65568 0.691359
+ 2.23e+11Hz -0.654414 0.692517
+ 2.231e+11Hz -0.653147 0.693672
+ 2.232e+11Hz -0.651877 0.694824
+ 2.233e+11Hz -0.650605 0.695974
+ 2.234e+11Hz -0.64933 0.697121
+ 2.235e+11Hz -0.648054 0.698266
+ 2.236e+11Hz -0.646775 0.699407
+ 2.237e+11Hz -0.645495 0.700546
+ 2.238e+11Hz -0.644212 0.701683
+ 2.239e+11Hz -0.642927 0.702817
+ 2.24e+11Hz -0.64164 0.703948
+ 2.241e+11Hz -0.64035 0.705076
+ 2.242e+11Hz -0.639059 0.706202
+ 2.243e+11Hz -0.637765 0.707325
+ 2.244e+11Hz -0.636469 0.708445
+ 2.245e+11Hz -0.635172 0.709563
+ 2.246e+11Hz -0.633872 0.710678
+ 2.247e+11Hz -0.632569 0.71179
+ 2.248e+11Hz -0.631265 0.712899
+ 2.249e+11Hz -0.629959 0.714005
+ 2.25e+11Hz -0.628651 0.715109
+ 2.251e+11Hz -0.62734 0.716209
+ 2.252e+11Hz -0.626028 0.717307
+ 2.253e+11Hz -0.624713 0.718402
+ 2.254e+11Hz -0.623397 0.719494
+ 2.255e+11Hz -0.622078 0.720584
+ 2.256e+11Hz -0.620757 0.72167
+ 2.257e+11Hz -0.619435 0.722754
+ 2.258e+11Hz -0.61811 0.723834
+ 2.259e+11Hz -0.616784 0.724912
+ 2.26e+11Hz -0.615455 0.725987
+ 2.261e+11Hz -0.614125 0.727058
+ 2.262e+11Hz -0.612792 0.728127
+ 2.263e+11Hz -0.611458 0.729193
+ 2.264e+11Hz -0.610122 0.730256
+ 2.265e+11Hz -0.608783 0.731315
+ 2.266e+11Hz -0.607443 0.732372
+ 2.267e+11Hz -0.606102 0.733426
+ 2.268e+11Hz -0.604758 0.734477
+ 2.269e+11Hz -0.603412 0.735524
+ 2.27e+11Hz -0.602065 0.736569
+ 2.271e+11Hz -0.600716 0.737611
+ 2.272e+11Hz -0.599365 0.738649
+ 2.273e+11Hz -0.598012 0.739684
+ 2.274e+11Hz -0.596658 0.740717
+ 2.275e+11Hz -0.595302 0.741746
+ 2.276e+11Hz -0.593944 0.742772
+ 2.277e+11Hz -0.592584 0.743795
+ 2.278e+11Hz -0.591223 0.744815
+ 2.279e+11Hz -0.589861 0.745831
+ 2.28e+11Hz -0.588496 0.746845
+ 2.281e+11Hz -0.58713 0.747855
+ 2.282e+11Hz -0.585763 0.748863
+ 2.283e+11Hz -0.584394 0.749867
+ 2.284e+11Hz -0.583023 0.750868
+ 2.285e+11Hz -0.581651 0.751865
+ 2.286e+11Hz -0.580278 0.75286
+ 2.287e+11Hz -0.578903 0.753851
+ 2.288e+11Hz -0.577526 0.75484
+ 2.289e+11Hz -0.576149 0.755825
+ 2.29e+11Hz -0.574769 0.756807
+ 2.291e+11Hz -0.573389 0.757785
+ 2.292e+11Hz -0.572007 0.758761
+ 2.293e+11Hz -0.570624 0.759733
+ 2.294e+11Hz -0.569239 0.760702
+ 2.295e+11Hz -0.567854 0.761668
+ 2.296e+11Hz -0.566467 0.762631
+ 2.297e+11Hz -0.565079 0.763591
+ 2.298e+11Hz -0.563689 0.764547
+ 2.299e+11Hz -0.562299 0.7655
+ 2.3e+11Hz -0.560907 0.76645
+ 2.301e+11Hz -0.559514 0.767397
+ 2.302e+11Hz -0.558121 0.768341
+ 2.303e+11Hz -0.556726 0.769282
+ 2.304e+11Hz -0.55533 0.770219
+ 2.305e+11Hz -0.553933 0.771154
+ 2.306e+11Hz -0.552535 0.772085
+ 2.307e+11Hz -0.551136 0.773013
+ 2.308e+11Hz -0.549736 0.773938
+ 2.309e+11Hz -0.548335 0.77486
+ 2.31e+11Hz -0.546933 0.775779
+ 2.311e+11Hz -0.545531 0.776695
+ 2.312e+11Hz -0.544127 0.777608
+ 2.313e+11Hz -0.542723 0.778517
+ 2.314e+11Hz -0.541318 0.779424
+ 2.315e+11Hz -0.539912 0.780328
+ 2.316e+11Hz -0.538505 0.781228
+ 2.317e+11Hz -0.537098 0.782126
+ 2.318e+11Hz -0.53569 0.78302
+ 2.319e+11Hz -0.534281 0.783912
+ 2.32e+11Hz -0.532871 0.784801
+ 2.321e+11Hz -0.531461 0.785686
+ 2.322e+11Hz -0.53005 0.786569
+ 2.323e+11Hz -0.528638 0.787449
+ 2.324e+11Hz -0.527226 0.788326
+ 2.325e+11Hz -0.525813 0.789201
+ 2.326e+11Hz -0.5244 0.790072
+ 2.327e+11Hz -0.522986 0.79094
+ 2.328e+11Hz -0.521572 0.791806
+ 2.329e+11Hz -0.520156 0.792669
+ 2.33e+11Hz -0.518741 0.793529
+ 2.331e+11Hz -0.517325 0.794386
+ 2.332e+11Hz -0.515908 0.795241
+ 2.333e+11Hz -0.514491 0.796093
+ 2.334e+11Hz -0.513073 0.796942
+ 2.335e+11Hz -0.511655 0.797789
+ 2.336e+11Hz -0.510237 0.798633
+ 2.337e+11Hz -0.508818 0.799474
+ 2.338e+11Hz -0.507398 0.800313
+ 2.339e+11Hz -0.505978 0.801149
+ 2.34e+11Hz -0.504558 0.801982
+ 2.341e+11Hz -0.503137 0.802813
+ 2.342e+11Hz -0.501716 0.803642
+ 2.343e+11Hz -0.500295 0.804468
+ 2.344e+11Hz -0.498873 0.805291
+ 2.345e+11Hz -0.49745 0.806112
+ 2.346e+11Hz -0.496028 0.806931
+ 2.347e+11Hz -0.494605 0.807747
+ 2.348e+11Hz -0.493181 0.808561
+ 2.349e+11Hz -0.491757 0.809372
+ 2.35e+11Hz -0.490333 0.810181
+ 2.351e+11Hz -0.488909 0.810988
+ 2.352e+11Hz -0.487484 0.811793
+ 2.353e+11Hz -0.486058 0.812595
+ 2.354e+11Hz -0.484633 0.813395
+ 2.355e+11Hz -0.483207 0.814192
+ 2.356e+11Hz -0.48178 0.814988
+ 2.357e+11Hz -0.480353 0.815781
+ 2.358e+11Hz -0.478926 0.816572
+ 2.359e+11Hz -0.477498 0.817361
+ 2.36e+11Hz -0.47607 0.818148
+ 2.361e+11Hz -0.474642 0.818933
+ 2.362e+11Hz -0.473213 0.819716
+ 2.363e+11Hz -0.471784 0.820496
+ 2.364e+11Hz -0.470355 0.821275
+ 2.365e+11Hz -0.468925 0.822051
+ 2.366e+11Hz -0.467494 0.822826
+ 2.367e+11Hz -0.466063 0.823598
+ 2.368e+11Hz -0.464632 0.824369
+ 2.369e+11Hz -0.4632 0.825138
+ 2.37e+11Hz -0.461768 0.825904
+ 2.371e+11Hz -0.460335 0.826669
+ 2.372e+11Hz -0.458902 0.827432
+ 2.373e+11Hz -0.457469 0.828193
+ 2.374e+11Hz -0.456034 0.828952
+ 2.375e+11Hz -0.4546 0.829709
+ 2.376e+11Hz -0.453165 0.830465
+ 2.377e+11Hz -0.451729 0.831218
+ 2.378e+11Hz -0.450293 0.83197
+ 2.379e+11Hz -0.448856 0.83272
+ 2.38e+11Hz -0.447419 0.833468
+ 2.381e+11Hz -0.445981 0.834215
+ 2.382e+11Hz -0.444542 0.83496
+ 2.383e+11Hz -0.443103 0.835703
+ 2.384e+11Hz -0.441663 0.836444
+ 2.385e+11Hz -0.440223 0.837184
+ 2.386e+11Hz -0.438782 0.837921
+ 2.387e+11Hz -0.43734 0.838658
+ 2.388e+11Hz -0.435897 0.839392
+ 2.389e+11Hz -0.434454 0.840125
+ 2.39e+11Hz -0.43301 0.840856
+ 2.391e+11Hz -0.431566 0.841585
+ 2.392e+11Hz -0.43012 0.842313
+ 2.393e+11Hz -0.428674 0.843039
+ 2.394e+11Hz -0.427227 0.843764
+ 2.395e+11Hz -0.42578 0.844487
+ 2.396e+11Hz -0.424331 0.845208
+ 2.397e+11Hz -0.422882 0.845928
+ 2.398e+11Hz -0.421432 0.846646
+ 2.399e+11Hz -0.419981 0.847362
+ 2.4e+11Hz -0.418529 0.848077
+ 2.401e+11Hz -0.417076 0.84879
+ 2.402e+11Hz -0.415623 0.849502
+ 2.403e+11Hz -0.414168 0.850212
+ 2.404e+11Hz -0.412712 0.85092
+ 2.405e+11Hz -0.411256 0.851627
+ 2.406e+11Hz -0.409798 0.852333
+ 2.407e+11Hz -0.40834 0.853036
+ 2.408e+11Hz -0.40688 0.853738
+ 2.409e+11Hz -0.40542 0.854439
+ 2.41e+11Hz -0.403959 0.855138
+ 2.411e+11Hz -0.402496 0.855835
+ 2.412e+11Hz -0.401032 0.856531
+ 2.413e+11Hz -0.399568 0.857225
+ 2.414e+11Hz -0.398102 0.857917
+ 2.415e+11Hz -0.396635 0.858608
+ 2.416e+11Hz -0.395167 0.859298
+ 2.417e+11Hz -0.393698 0.859985
+ 2.418e+11Hz -0.392227 0.860671
+ 2.419e+11Hz -0.390756 0.861356
+ 2.42e+11Hz -0.389283 0.862039
+ 2.421e+11Hz -0.387809 0.86272
+ 2.422e+11Hz -0.386334 0.8634
+ 2.423e+11Hz -0.384858 0.864078
+ 2.424e+11Hz -0.38338 0.864754
+ 2.425e+11Hz -0.381901 0.865429
+ 2.426e+11Hz -0.380421 0.866102
+ 2.427e+11Hz -0.37894 0.866773
+ 2.428e+11Hz -0.377457 0.867443
+ 2.429e+11Hz -0.375973 0.868111
+ 2.43e+11Hz -0.374488 0.868777
+ 2.431e+11Hz -0.373002 0.869442
+ 2.432e+11Hz -0.371514 0.870105
+ 2.433e+11Hz -0.370024 0.870767
+ 2.434e+11Hz -0.368534 0.871426
+ 2.435e+11Hz -0.367042 0.872084
+ 2.436e+11Hz -0.365548 0.87274
+ 2.437e+11Hz -0.364054 0.873395
+ 2.438e+11Hz -0.362558 0.874048
+ 2.439e+11Hz -0.36106 0.874699
+ 2.44e+11Hz -0.359561 0.875348
+ 2.441e+11Hz -0.35806 0.875995
+ 2.442e+11Hz -0.356559 0.876641
+ 2.443e+11Hz -0.355055 0.877285
+ 2.444e+11Hz -0.35355 0.877927
+ 2.445e+11Hz -0.352044 0.878568
+ 2.446e+11Hz -0.350536 0.879206
+ 2.447e+11Hz -0.349027 0.879843
+ 2.448e+11Hz -0.347517 0.880478
+ 2.449e+11Hz -0.346004 0.881111
+ 2.45e+11Hz -0.344491 0.881742
+ 2.451e+11Hz -0.342975 0.882371
+ 2.452e+11Hz -0.341459 0.882999
+ 2.453e+11Hz -0.33994 0.883624
+ 2.454e+11Hz -0.33842 0.884248
+ 2.455e+11Hz -0.336899 0.88487
+ 2.456e+11Hz -0.335376 0.88549
+ 2.457e+11Hz -0.333852 0.886108
+ 2.458e+11Hz -0.332326 0.886724
+ 2.459e+11Hz -0.330798 0.887338
+ 2.46e+11Hz -0.329269 0.887951
+ 2.461e+11Hz -0.327738 0.888561
+ 2.462e+11Hz -0.326205 0.889169
+ 2.463e+11Hz -0.324671 0.889776
+ 2.464e+11Hz -0.323136 0.89038
+ 2.465e+11Hz -0.321599 0.890982
+ 2.466e+11Hz -0.32006 0.891583
+ 2.467e+11Hz -0.318519 0.892181
+ 2.468e+11Hz -0.316977 0.892777
+ 2.469e+11Hz -0.315434 0.893372
+ 2.47e+11Hz -0.313888 0.893964
+ 2.471e+11Hz -0.312341 0.894554
+ 2.472e+11Hz -0.310793 0.895142
+ 2.473e+11Hz -0.309242 0.895728
+ 2.474e+11Hz -0.30769 0.896312
+ 2.475e+11Hz -0.306137 0.896894
+ 2.476e+11Hz -0.304581 0.897474
+ 2.477e+11Hz -0.303024 0.898051
+ 2.478e+11Hz -0.301466 0.898627
+ 2.479e+11Hz -0.299905 0.8992
+ 2.48e+11Hz -0.298343 0.899771
+ 2.481e+11Hz -0.296779 0.900341
+ 2.482e+11Hz -0.295214 0.900907
+ 2.483e+11Hz -0.293647 0.901472
+ 2.484e+11Hz -0.292078 0.902035
+ 2.485e+11Hz -0.290507 0.902595
+ 2.486e+11Hz -0.288935 0.903153
+ 2.487e+11Hz -0.287361 0.903709
+ 2.488e+11Hz -0.285785 0.904262
+ 2.489e+11Hz -0.284208 0.904814
+ 2.49e+11Hz -0.282628 0.905363
+ 2.491e+11Hz -0.281047 0.90591
+ 2.492e+11Hz -0.279465 0.906454
+ 2.493e+11Hz -0.27788 0.906996
+ 2.494e+11Hz -0.276294 0.907536
+ 2.495e+11Hz -0.274706 0.908074
+ 2.496e+11Hz -0.273116 0.908609
+ 2.497e+11Hz -0.271524 0.909142
+ 2.498e+11Hz -0.269931 0.909672
+ 2.499e+11Hz -0.268336 0.9102
+ 2.5e+11Hz -0.266739 0.910726
+ 2.501e+11Hz -0.26514 0.911249
+ 2.502e+11Hz -0.26354 0.91177
+ 2.503e+11Hz -0.261937 0.912289
+ 2.504e+11Hz -0.260333 0.912805
+ 2.505e+11Hz -0.258727 0.913318
+ 2.506e+11Hz -0.257119 0.913829
+ 2.507e+11Hz -0.25551 0.914338
+ 2.508e+11Hz -0.253898 0.914844
+ 2.509e+11Hz -0.252285 0.915347
+ 2.51e+11Hz -0.25067 0.915848
+ 2.511e+11Hz -0.249053 0.916346
+ 2.512e+11Hz -0.247434 0.916842
+ 2.513e+11Hz -0.245814 0.917335
+ 2.514e+11Hz -0.244191 0.917826
+ 2.515e+11Hz -0.242567 0.918314
+ 2.516e+11Hz -0.240941 0.918799
+ 2.517e+11Hz -0.239313 0.919282
+ 2.518e+11Hz -0.237683 0.919762
+ 2.519e+11Hz -0.236051 0.920239
+ 2.52e+11Hz -0.234418 0.920714
+ 2.521e+11Hz -0.232782 0.921185
+ 2.522e+11Hz -0.231145 0.921654
+ 2.523e+11Hz -0.229506 0.922121
+ 2.524e+11Hz -0.227864 0.922584
+ 2.525e+11Hz -0.226222 0.923045
+ 2.526e+11Hz -0.224577 0.923502
+ 2.527e+11Hz -0.22293 0.923957
+ 2.528e+11Hz -0.221282 0.924409
+ 2.529e+11Hz -0.219631 0.924859
+ 2.53e+11Hz -0.217979 0.925305
+ 2.531e+11Hz -0.216325 0.925748
+ 2.532e+11Hz -0.214669 0.926188
+ 2.533e+11Hz -0.213011 0.926626
+ 2.534e+11Hz -0.211351 0.92706
+ 2.535e+11Hz -0.20969 0.927491
+ 2.536e+11Hz -0.208026 0.92792
+ 2.537e+11Hz -0.206361 0.928345
+ 2.538e+11Hz -0.204694 0.928767
+ 2.539e+11Hz -0.203025 0.929186
+ 2.54e+11Hz -0.201354 0.929602
+ 2.541e+11Hz -0.199682 0.930014
+ 2.542e+11Hz -0.198007 0.930424
+ 2.543e+11Hz -0.196331 0.93083
+ 2.544e+11Hz -0.194653 0.931233
+ 2.545e+11Hz -0.192973 0.931633
+ 2.546e+11Hz -0.191291 0.932029
+ 2.547e+11Hz -0.189608 0.932422
+ 2.548e+11Hz -0.187923 0.932812
+ 2.549e+11Hz -0.186235 0.933199
+ 2.55e+11Hz -0.184547 0.933582
+ 2.551e+11Hz -0.182856 0.933961
+ 2.552e+11Hz -0.181164 0.934338
+ 2.553e+11Hz -0.17947 0.93471
+ 2.554e+11Hz -0.177774 0.93508
+ 2.555e+11Hz -0.176077 0.935445
+ 2.556e+11Hz -0.174378 0.935808
+ 2.557e+11Hz -0.172677 0.936166
+ 2.558e+11Hz -0.170974 0.936522
+ 2.559e+11Hz -0.16927 0.936873
+ 2.56e+11Hz -0.167564 0.937221
+ 2.561e+11Hz -0.165857 0.937565
+ 2.562e+11Hz -0.164148 0.937906
+ 2.563e+11Hz -0.162437 0.938243
+ 2.564e+11Hz -0.160725 0.938576
+ 2.565e+11Hz -0.159011 0.938906
+ 2.566e+11Hz -0.157296 0.939231
+ 2.567e+11Hz -0.155579 0.939553
+ 2.568e+11Hz -0.153861 0.939872
+ 2.569e+11Hz -0.152141 0.940186
+ 2.57e+11Hz -0.15042 0.940496
+ 2.571e+11Hz -0.148697 0.940803
+ 2.572e+11Hz -0.146973 0.941106
+ 2.573e+11Hz -0.145248 0.941405
+ 2.574e+11Hz -0.143521 0.9417
+ 2.575e+11Hz -0.141793 0.941991
+ 2.576e+11Hz -0.140063 0.942278
+ 2.577e+11Hz -0.138333 0.942561
+ 2.578e+11Hz -0.136601 0.94284
+ 2.579e+11Hz -0.134867 0.943115
+ 2.58e+11Hz -0.133133 0.943385
+ 2.581e+11Hz -0.131397 0.943652
+ 2.582e+11Hz -0.12966 0.943915
+ 2.583e+11Hz -0.127922 0.944174
+ 2.584e+11Hz -0.126183 0.944429
+ 2.585e+11Hz -0.124442 0.944679
+ 2.586e+11Hz -0.122701 0.944925
+ 2.587e+11Hz -0.120959 0.945168
+ 2.588e+11Hz -0.119215 0.945406
+ 2.589e+11Hz -0.117471 0.94564
+ 2.59e+11Hz -0.115725 0.945869
+ 2.591e+11Hz -0.113979 0.946095
+ 2.592e+11Hz -0.112232 0.946316
+ 2.593e+11Hz -0.110484 0.946533
+ 2.594e+11Hz -0.108735 0.946746
+ 2.595e+11Hz -0.106985 0.946955
+ 2.596e+11Hz -0.105235 0.947159
+ 2.597e+11Hz -0.103484 0.947359
+ 2.598e+11Hz -0.101732 0.947555
+ 2.599e+11Hz -0.0999791 0.947746
+ 2.6e+11Hz -0.0982258 0.947934
+ 2.601e+11Hz -0.0964719 0.948116
+ 2.602e+11Hz -0.0947175 0.948295
+ 2.603e+11Hz -0.0929624 0.94847
+ 2.604e+11Hz -0.0912069 0.94864
+ 2.605e+11Hz -0.0894508 0.948805
+ 2.606e+11Hz -0.0876943 0.948967
+ 2.607e+11Hz -0.0859373 0.949124
+ 2.608e+11Hz -0.08418 0.949277
+ 2.609e+11Hz -0.0824222 0.949425
+ 2.61e+11Hz -0.0806641 0.94957
+ 2.611e+11Hz -0.0789058 0.94971
+ 2.612e+11Hz -0.0771471 0.949845
+ 2.613e+11Hz -0.0753882 0.949976
+ 2.614e+11Hz -0.073629 0.950103
+ 2.615e+11Hz -0.0718697 0.950226
+ 2.616e+11Hz -0.0701102 0.950345
+ 2.617e+11Hz -0.0683506 0.950459
+ 2.618e+11Hz -0.0665909 0.950568
+ 2.619e+11Hz -0.0648312 0.950674
+ 2.62e+11Hz -0.0630714 0.950775
+ 2.621e+11Hz -0.0613115 0.950872
+ 2.622e+11Hz -0.0595517 0.950965
+ 2.623e+11Hz -0.057792 0.951053
+ 2.624e+11Hz -0.0560323 0.951138
+ 2.625e+11Hz -0.0542728 0.951218
+ 2.626e+11Hz -0.0525133 0.951293
+ 2.627e+11Hz -0.050754 0.951365
+ 2.628e+11Hz -0.048995 0.951432
+ 2.629e+11Hz -0.0472361 0.951495
+ 2.63e+11Hz -0.0454774 0.951554
+ 2.631e+11Hz -0.0437191 0.951609
+ 2.632e+11Hz -0.041961 0.95166
+ 2.633e+11Hz -0.0402032 0.951706
+ 2.634e+11Hz -0.0384458 0.951749
+ 2.635e+11Hz -0.0366887 0.951787
+ 2.636e+11Hz -0.034932 0.951821
+ 2.637e+11Hz -0.0331757 0.951851
+ 2.638e+11Hz -0.0314199 0.951877
+ 2.639e+11Hz -0.0296645 0.951898
+ 2.64e+11Hz -0.0279096 0.951916
+ 2.641e+11Hz -0.0261552 0.95193
+ 2.642e+11Hz -0.0244013 0.95194
+ 2.643e+11Hz -0.0226479 0.951945
+ 2.644e+11Hz -0.0208951 0.951947
+ 2.645e+11Hz -0.0191429 0.951945
+ 2.646e+11Hz -0.0173912 0.951939
+ 2.647e+11Hz -0.0156402 0.951928
+ 2.648e+11Hz -0.0138898 0.951914
+ 2.649e+11Hz -0.01214 0.951896
+ 2.65e+11Hz -0.0103909 0.951874
+ 2.651e+11Hz -0.0086425 0.951849
+ 2.652e+11Hz -0.00689477 0.951819
+ 2.653e+11Hz -0.00514776 0.951785
+ 2.654e+11Hz -0.00340146 0.951748
+ 2.655e+11Hz -0.00165591 0.951707
+ 2.656e+11Hz 8.89001e-05 0.951662
+ 2.657e+11Hz 0.00183294 0.951613
+ 2.658e+11Hz 0.00357621 0.951561
+ 2.659e+11Hz 0.00531869 0.951504
+ 2.66e+11Hz 0.00706037 0.951445
+ 2.661e+11Hz 0.00880125 0.951381
+ 2.662e+11Hz 0.0105413 0.951313
+ 2.663e+11Hz 0.0122805 0.951242
+ 2.664e+11Hz 0.0140189 0.951168
+ 2.665e+11Hz 0.0157564 0.951089
+ 2.666e+11Hz 0.0174931 0.951007
+ 2.667e+11Hz 0.0192289 0.950922
+ 2.668e+11Hz 0.0209638 0.950833
+ 2.669e+11Hz 0.0226979 0.95074
+ 2.67e+11Hz 0.024431 0.950643
+ 2.671e+11Hz 0.0261633 0.950544
+ 2.672e+11Hz 0.0278947 0.95044
+ 2.673e+11Hz 0.0296251 0.950333
+ 2.674e+11Hz 0.0313546 0.950223
+ 2.675e+11Hz 0.0330832 0.950109
+ 2.676e+11Hz 0.0348109 0.949991
+ 2.677e+11Hz 0.0365377 0.94987
+ 2.678e+11Hz 0.0382635 0.949746
+ 2.679e+11Hz 0.0399883 0.949618
+ 2.68e+11Hz 0.0417123 0.949487
+ 2.681e+11Hz 0.0434352 0.949352
+ 2.682e+11Hz 0.0451572 0.949214
+ 2.683e+11Hz 0.0468783 0.949072
+ 2.684e+11Hz 0.0485984 0.948927
+ 2.685e+11Hz 0.0503175 0.948779
+ 2.686e+11Hz 0.0520357 0.948627
+ 2.687e+11Hz 0.0537528 0.948472
+ 2.688e+11Hz 0.055469 0.948314
+ 2.689e+11Hz 0.0571842 0.948152
+ 2.69e+11Hz 0.0588985 0.947987
+ 2.691e+11Hz 0.0606117 0.947819
+ 2.692e+11Hz 0.062324 0.947647
+ 2.693e+11Hz 0.0640352 0.947472
+ 2.694e+11Hz 0.0657455 0.947294
+ 2.695e+11Hz 0.0674548 0.947113
+ 2.696e+11Hz 0.069163 0.946928
+ 2.697e+11Hz 0.0708703 0.94674
+ 2.698e+11Hz 0.0725765 0.946549
+ 2.699e+11Hz 0.0742817 0.946354
+ 2.7e+11Hz 0.0759859 0.946156
+ 2.701e+11Hz 0.0776891 0.945955
+ 2.702e+11Hz 0.0793913 0.945751
+ 2.703e+11Hz 0.0810924 0.945543
+ 2.704e+11Hz 0.0827925 0.945332
+ 2.705e+11Hz 0.0844915 0.945118
+ 2.706e+11Hz 0.0861895 0.944901
+ 2.707e+11Hz 0.0878865 0.944681
+ 2.708e+11Hz 0.0895824 0.944457
+ 2.709e+11Hz 0.0912772 0.94423
+ 2.71e+11Hz 0.092971 0.944
+ 2.711e+11Hz 0.0946637 0.943767
+ 2.712e+11Hz 0.0963553 0.943531
+ 2.713e+11Hz 0.0980458 0.943291
+ 2.714e+11Hz 0.0997353 0.943049
+ 2.715e+11Hz 0.101424 0.942803
+ 2.716e+11Hz 0.103111 0.942553
+ 2.717e+11Hz 0.104797 0.942301
+ 2.718e+11Hz 0.106482 0.942046
+ 2.719e+11Hz 0.108166 0.941787
+ 2.72e+11Hz 0.109849 0.941525
+ 2.721e+11Hz 0.11153 0.941261
+ 2.722e+11Hz 0.113211 0.940993
+ 2.723e+11Hz 0.11489 0.940721
+ 2.724e+11Hz 0.116568 0.940447
+ 2.725e+11Hz 0.118245 0.94017
+ 2.726e+11Hz 0.119921 0.939889
+ 2.727e+11Hz 0.121596 0.939605
+ 2.728e+11Hz 0.123269 0.939318
+ 2.729e+11Hz 0.124941 0.939028
+ 2.73e+11Hz 0.126612 0.938735
+ 2.731e+11Hz 0.128282 0.938439
+ 2.732e+11Hz 0.12995 0.93814
+ 2.733e+11Hz 0.131617 0.937838
+ 2.734e+11Hz 0.133283 0.937532
+ 2.735e+11Hz 0.134948 0.937224
+ 2.736e+11Hz 0.136611 0.936912
+ 2.737e+11Hz 0.138273 0.936597
+ 2.738e+11Hz 0.139934 0.93628
+ 2.739e+11Hz 0.141593 0.935959
+ 2.74e+11Hz 0.143251 0.935635
+ 2.741e+11Hz 0.144908 0.935308
+ 2.742e+11Hz 0.146563 0.934978
+ 2.743e+11Hz 0.148217 0.934646
+ 2.744e+11Hz 0.149869 0.93431
+ 2.745e+11Hz 0.15152 0.933971
+ 2.746e+11Hz 0.15317 0.933629
+ 2.747e+11Hz 0.154818 0.933284
+ 2.748e+11Hz 0.156465 0.932936
+ 2.749e+11Hz 0.15811 0.932586
+ 2.75e+11Hz 0.159754 0.932232
+ 2.751e+11Hz 0.161396 0.931875
+ 2.752e+11Hz 0.163037 0.931516
+ 2.753e+11Hz 0.164676 0.931153
+ 2.754e+11Hz 0.166313 0.930788
+ 2.755e+11Hz 0.16795 0.93042
+ 2.756e+11Hz 0.169584 0.930049
+ 2.757e+11Hz 0.171217 0.929675
+ 2.758e+11Hz 0.172848 0.929298
+ 2.759e+11Hz 0.174478 0.928918
+ 2.76e+11Hz 0.176106 0.928536
+ 2.761e+11Hz 0.177733 0.928151
+ 2.762e+11Hz 0.179358 0.927763
+ 2.763e+11Hz 0.180981 0.927373
+ 2.764e+11Hz 0.182603 0.926979
+ 2.765e+11Hz 0.184223 0.926583
+ 2.766e+11Hz 0.185841 0.926184
+ 2.767e+11Hz 0.187457 0.925783
+ 2.768e+11Hz 0.189072 0.925379
+ 2.769e+11Hz 0.190685 0.924973
+ 2.77e+11Hz 0.192297 0.924563
+ 2.771e+11Hz 0.193906 0.924152
+ 2.772e+11Hz 0.195514 0.923737
+ 2.773e+11Hz 0.19712 0.92332
+ 2.774e+11Hz 0.198725 0.922901
+ 2.775e+11Hz 0.200327 0.922479
+ 2.776e+11Hz 0.201928 0.922055
+ 2.777e+11Hz 0.203527 0.921628
+ 2.778e+11Hz 0.205125 0.921199
+ 2.779e+11Hz 0.20672 0.920767
+ 2.78e+11Hz 0.208314 0.920333
+ 2.781e+11Hz 0.209906 0.919897
+ 2.782e+11Hz 0.211496 0.919459
+ 2.783e+11Hz 0.213084 0.919018
+ 2.784e+11Hz 0.214671 0.918575
+ 2.785e+11Hz 0.216256 0.918129
+ 2.786e+11Hz 0.217839 0.917682
+ 2.787e+11Hz 0.21942 0.917232
+ 2.788e+11Hz 0.220999 0.916781
+ 2.789e+11Hz 0.222577 0.916327
+ 2.79e+11Hz 0.224153 0.915871
+ 2.791e+11Hz 0.225727 0.915412
+ 2.792e+11Hz 0.227299 0.914952
+ 2.793e+11Hz 0.228869 0.91449
+ 2.794e+11Hz 0.230438 0.914026
+ 2.795e+11Hz 0.232005 0.91356
+ 2.796e+11Hz 0.23357 0.913092
+ 2.797e+11Hz 0.235134 0.912622
+ 2.798e+11Hz 0.236695 0.91215
+ 2.799e+11Hz 0.238255 0.911677
+ 2.8e+11Hz 0.239813 0.911201
+ 2.801e+11Hz 0.24137 0.910724
+ 2.802e+11Hz 0.242925 0.910245
+ 2.803e+11Hz 0.244478 0.909764
+ 2.804e+11Hz 0.246029 0.909282
+ 2.805e+11Hz 0.247579 0.908798
+ 2.806e+11Hz 0.249127 0.908312
+ 2.807e+11Hz 0.250674 0.907824
+ 2.808e+11Hz 0.252219 0.907335
+ 2.809e+11Hz 0.253762 0.906844
+ 2.81e+11Hz 0.255304 0.906352
+ 2.811e+11Hz 0.256845 0.905858
+ 2.812e+11Hz 0.258383 0.905363
+ 2.813e+11Hz 0.259921 0.904866
+ 2.814e+11Hz 0.261456 0.904368
+ 2.815e+11Hz 0.262991 0.903868
+ 2.816e+11Hz 0.264524 0.903367
+ 2.817e+11Hz 0.266055 0.902864
+ 2.818e+11Hz 0.267585 0.90236
+ 2.819e+11Hz 0.269114 0.901855
+ 2.82e+11Hz 0.270641 0.901348
+ 2.821e+11Hz 0.272167 0.90084
+ 2.822e+11Hz 0.273692 0.900331
+ 2.823e+11Hz 0.275215 0.89982
+ 2.824e+11Hz 0.276738 0.899308
+ 2.825e+11Hz 0.278259 0.898795
+ 2.826e+11Hz 0.279779 0.89828
+ 2.827e+11Hz 0.281297 0.897764
+ 2.828e+11Hz 0.282815 0.897247
+ 2.829e+11Hz 0.284332 0.896729
+ 2.83e+11Hz 0.285847 0.896209
+ 2.831e+11Hz 0.287361 0.895688
+ 2.832e+11Hz 0.288875 0.895166
+ 2.833e+11Hz 0.290387 0.894643
+ 2.834e+11Hz 0.291899 0.894118
+ 2.835e+11Hz 0.29341 0.893593
+ 2.836e+11Hz 0.29492 0.893066
+ 2.837e+11Hz 0.296429 0.892538
+ 2.838e+11Hz 0.297937 0.892009
+ 2.839e+11Hz 0.299444 0.891478
+ 2.84e+11Hz 0.300951 0.890947
+ 2.841e+11Hz 0.302457 0.890414
+ 2.842e+11Hz 0.303962 0.88988
+ 2.843e+11Hz 0.305467 0.889345
+ 2.844e+11Hz 0.306971 0.888808
+ 2.845e+11Hz 0.308474 0.888271
+ 2.846e+11Hz 0.309977 0.887732
+ 2.847e+11Hz 0.31148 0.887192
+ 2.848e+11Hz 0.312982 0.886651
+ 2.849e+11Hz 0.314483 0.886108
+ 2.85e+11Hz 0.315984 0.885564
+ 2.851e+11Hz 0.317485 0.885019
+ 2.852e+11Hz 0.318985 0.884473
+ 2.853e+11Hz 0.320485 0.883926
+ 2.854e+11Hz 0.321985 0.883377
+ 2.855e+11Hz 0.323485 0.882827
+ 2.856e+11Hz 0.324984 0.882275
+ 2.857e+11Hz 0.326483 0.881722
+ 2.858e+11Hz 0.327982 0.881168
+ 2.859e+11Hz 0.329481 0.880613
+ 2.86e+11Hz 0.330979 0.880056
+ 2.861e+11Hz 0.332478 0.879497
+ 2.862e+11Hz 0.333976 0.878937
+ 2.863e+11Hz 0.335475 0.878376
+ 2.864e+11Hz 0.336973 0.877813
+ 2.865e+11Hz 0.338472 0.877249
+ 2.866e+11Hz 0.33997 0.876683
+ 2.867e+11Hz 0.341469 0.876116
+ 2.868e+11Hz 0.342967 0.875546
+ 2.869e+11Hz 0.344466 0.874976
+ 2.87e+11Hz 0.345965 0.874404
+ 2.871e+11Hz 0.347464 0.873829
+ 2.872e+11Hz 0.348963 0.873254
+ 2.873e+11Hz 0.350463 0.872676
+ 2.874e+11Hz 0.351962 0.872097
+ 2.875e+11Hz 0.353462 0.871516
+ 2.876e+11Hz 0.354962 0.870933
+ 2.877e+11Hz 0.356462 0.870349
+ 2.878e+11Hz 0.357963 0.869762
+ 2.879e+11Hz 0.359463 0.869173
+ 2.88e+11Hz 0.360965 0.868583
+ 2.881e+11Hz 0.362466 0.86799
+ 2.882e+11Hz 0.363968 0.867396
+ 2.883e+11Hz 0.36547 0.866799
+ 2.884e+11Hz 0.366972 0.8662
+ 2.885e+11Hz 0.368474 0.8656
+ 2.886e+11Hz 0.369977 0.864997
+ 2.887e+11Hz 0.371481 0.864391
+ 2.888e+11Hz 0.372984 0.863784
+ 2.889e+11Hz 0.374488 0.863174
+ 2.89e+11Hz 0.375993 0.862562
+ 2.891e+11Hz 0.377497 0.861948
+ 2.892e+11Hz 0.379002 0.861331
+ 2.893e+11Hz 0.380507 0.860711
+ 2.894e+11Hz 0.382013 0.86009
+ 2.895e+11Hz 0.383519 0.859466
+ 2.896e+11Hz 0.385025 0.858839
+ 2.897e+11Hz 0.386532 0.85821
+ 2.898e+11Hz 0.388039 0.857578
+ 2.899e+11Hz 0.389546 0.856943
+ 2.9e+11Hz 0.391054 0.856306
+ 2.901e+11Hz 0.392561 0.855666
+ 2.902e+11Hz 0.394069 0.855023
+ 2.903e+11Hz 0.395578 0.854378
+ 2.904e+11Hz 0.397086 0.85373
+ 2.905e+11Hz 0.398595 0.853079
+ 2.906e+11Hz 0.400104 0.852425
+ 2.907e+11Hz 0.401613 0.851768
+ 2.908e+11Hz 0.403123 0.851108
+ 2.909e+11Hz 0.404632 0.850445
+ 2.91e+11Hz 0.406142 0.849779
+ 2.911e+11Hz 0.407652 0.849111
+ 2.912e+11Hz 0.409162 0.848439
+ 2.913e+11Hz 0.410672 0.847764
+ 2.914e+11Hz 0.412182 0.847086
+ 2.915e+11Hz 0.413692 0.846405
+ 2.916e+11Hz 0.415202 0.84572
+ 2.917e+11Hz 0.416712 0.845033
+ 2.918e+11Hz 0.418222 0.844342
+ 2.919e+11Hz 0.419732 0.843648
+ 2.92e+11Hz 0.421242 0.842951
+ 2.921e+11Hz 0.422752 0.84225
+ 2.922e+11Hz 0.424261 0.841546
+ 2.923e+11Hz 0.425771 0.840839
+ 2.924e+11Hz 0.42728 0.840128
+ 2.925e+11Hz 0.428789 0.839414
+ 2.926e+11Hz 0.430298 0.838697
+ 2.927e+11Hz 0.431807 0.837976
+ 2.928e+11Hz 0.433315 0.837252
+ 2.929e+11Hz 0.434823 0.836524
+ 2.93e+11Hz 0.43633 0.835793
+ 2.931e+11Hz 0.437837 0.835059
+ 2.932e+11Hz 0.439344 0.834321
+ 2.933e+11Hz 0.44085 0.833579
+ 2.934e+11Hz 0.442356 0.832834
+ 2.935e+11Hz 0.443861 0.832085
+ 2.936e+11Hz 0.445365 0.831333
+ 2.937e+11Hz 0.446869 0.830577
+ 2.938e+11Hz 0.448373 0.829818
+ 2.939e+11Hz 0.449875 0.829055
+ 2.94e+11Hz 0.451377 0.828289
+ 2.941e+11Hz 0.452878 0.827519
+ 2.942e+11Hz 0.454379 0.826745
+ 2.943e+11Hz 0.455879 0.825968
+ 2.944e+11Hz 0.457377 0.825187
+ 2.945e+11Hz 0.458875 0.824403
+ 2.946e+11Hz 0.460373 0.823615
+ 2.947e+11Hz 0.461869 0.822824
+ 2.948e+11Hz 0.463364 0.822028
+ 2.949e+11Hz 0.464858 0.82123
+ 2.95e+11Hz 0.466351 0.820427
+ 2.951e+11Hz 0.467844 0.819622
+ 2.952e+11Hz 0.469335 0.818812
+ 2.953e+11Hz 0.470825 0.817999
+ 2.954e+11Hz 0.472314 0.817183
+ 2.955e+11Hz 0.473801 0.816362
+ 2.956e+11Hz 0.475288 0.815539
+ 2.957e+11Hz 0.476773 0.814711
+ 2.958e+11Hz 0.478257 0.813881
+ 2.959e+11Hz 0.47974 0.813046
+ 2.96e+11Hz 0.481222 0.812208
+ 2.961e+11Hz 0.482702 0.811367
+ 2.962e+11Hz 0.484181 0.810522
+ 2.963e+11Hz 0.485658 0.809674
+ 2.964e+11Hz 0.487134 0.808822
+ 2.965e+11Hz 0.488609 0.807966
+ 2.966e+11Hz 0.490082 0.807107
+ 2.967e+11Hz 0.491553 0.806245
+ 2.968e+11Hz 0.493024 0.805379
+ 2.969e+11Hz 0.494492 0.80451
+ 2.97e+11Hz 0.495959 0.803637
+ 2.971e+11Hz 0.497425 0.802761
+ 2.972e+11Hz 0.498889 0.801882
+ 2.973e+11Hz 0.500351 0.800999
+ 2.974e+11Hz 0.501812 0.800113
+ 2.975e+11Hz 0.503271 0.799223
+ 2.976e+11Hz 0.504728 0.798331
+ 2.977e+11Hz 0.506184 0.797434
+ 2.978e+11Hz 0.507638 0.796535
+ 2.979e+11Hz 0.50909 0.795632
+ 2.98e+11Hz 0.510541 0.794726
+ 2.981e+11Hz 0.51199 0.793817
+ 2.982e+11Hz 0.513437 0.792904
+ 2.983e+11Hz 0.514882 0.791989
+ 2.984e+11Hz 0.516326 0.79107
+ 2.985e+11Hz 0.517768 0.790148
+ 2.986e+11Hz 0.519208 0.789222
+ 2.987e+11Hz 0.520646 0.788294
+ 2.988e+11Hz 0.522082 0.787362
+ 2.989e+11Hz 0.523516 0.786427
+ 2.99e+11Hz 0.524949 0.785489
+ 2.991e+11Hz 0.52638 0.784548
+ 2.992e+11Hz 0.527809 0.783604
+ 2.993e+11Hz 0.529236 0.782657
+ 2.994e+11Hz 0.530661 0.781707
+ 2.995e+11Hz 0.532084 0.780754
+ 2.996e+11Hz 0.533505 0.779797
+ 2.997e+11Hz 0.534925 0.778838
+ 2.998e+11Hz 0.536342 0.777876
+ 2.999e+11Hz 0.537758 0.77691
+ 3e+11Hz 0.539172 0.775942
+ ]

A22 %vd(20 3) %vd(22, 3) xfer4
.model xfer4 xfer R_I=true table=[
+ 0Hz 0.0101636 0
+ 1e+08Hz 0.0101645 2.67419e-05
+ 2e+08Hz 0.010167 5.34355e-05
+ 3e+08Hz 0.0101713 8.00327e-05
+ 4e+08Hz 0.0101773 0.000106485
+ 5e+08Hz 0.010185 0.000132746
+ 6e+08Hz 0.0101944 0.000158766
+ 7e+08Hz 0.0102055 0.000184498
+ 8e+08Hz 0.0102183 0.000209896
+ 9e+08Hz 0.0102327 0.000234912
+ 1e+09Hz 0.0102488 0.0002595
+ 1.1e+09Hz 0.0102665 0.000283614
+ 1.2e+09Hz 0.0102859 0.000307209
+ 1.3e+09Hz 0.0103068 0.000330239
+ 1.4e+09Hz 0.0103294 0.000352661
+ 1.5e+09Hz 0.0103535 0.000374431
+ 1.6e+09Hz 0.0103792 0.000395505
+ 1.7e+09Hz 0.0104064 0.000415842
+ 1.8e+09Hz 0.0104352 0.000435401
+ 1.9e+09Hz 0.0104654 0.000454139
+ 2e+09Hz 0.010497 0.000472019
+ 2.1e+09Hz 0.0105301 0.000489
+ 2.2e+09Hz 0.0105646 0.000505045
+ 2.3e+09Hz 0.0106005 0.000520116
+ 2.4e+09Hz 0.0106377 0.000534178
+ 2.5e+09Hz 0.0106763 0.000547196
+ 2.6e+09Hz 0.0107161 0.000559136
+ 2.7e+09Hz 0.0107572 0.000569964
+ 2.8e+09Hz 0.0107995 0.000579649
+ 2.9e+09Hz 0.0108429 0.000588161
+ 3e+09Hz 0.0108875 0.000595469
+ 3.1e+09Hz 0.0109333 0.000601546
+ 3.2e+09Hz 0.01098 0.000606364
+ 3.3e+09Hz 0.0110279 0.000609898
+ 3.4e+09Hz 0.0110767 0.000612122
+ 3.5e+09Hz 0.0111265 0.000613014
+ 3.6e+09Hz 0.0111772 0.000612551
+ 3.7e+09Hz 0.0112288 0.000610712
+ 3.8e+09Hz 0.0112812 0.000607479
+ 3.9e+09Hz 0.0113345 0.000602831
+ 4e+09Hz 0.0113884 0.000596753
+ 4.1e+09Hz 0.0114431 0.000589229
+ 4.2e+09Hz 0.0114985 0.000580244
+ 4.3e+09Hz 0.0115546 0.000569785
+ 4.4e+09Hz 0.0116112 0.00055784
+ 4.5e+09Hz 0.0116683 0.000544399
+ 4.6e+09Hz 0.011726 0.000529453
+ 4.7e+09Hz 0.0117841 0.000512993
+ 4.8e+09Hz 0.0118427 0.000495014
+ 4.9e+09Hz 0.0119017 0.000475509
+ 5e+09Hz 0.0119609 0.000454474
+ 5.1e+09Hz 0.0120205 0.000431908
+ 5.2e+09Hz 0.0120804 0.000407808
+ 5.3e+09Hz 0.0121404 0.000382173
+ 5.4e+09Hz 0.0122007 0.000355005
+ 5.5e+09Hz 0.0122611 0.000326306
+ 5.6e+09Hz 0.0123215 0.000296079
+ 5.7e+09Hz 0.012382 0.000264329
+ 5.8e+09Hz 0.0124426 0.00023106
+ 5.9e+09Hz 0.0125031 0.00019628
+ 6e+09Hz 0.0125635 0.000159997
+ 6.1e+09Hz 0.0126238 0.000122219
+ 6.2e+09Hz 0.012684 8.29562e-05
+ 6.3e+09Hz 0.012744 4.22199e-05
+ 6.4e+09Hz 0.0128038 2.19349e-08
+ 6.5e+09Hz 0.0128634 -4.36247e-05
+ 6.6e+09Hz 0.0129226 -8.8706e-05
+ 6.7e+09Hz 0.0129815 -0.000135207
+ 6.8e+09Hz 0.0130401 -0.000183112
+ 6.9e+09Hz 0.0130983 -0.000232405
+ 7e+09Hz 0.013156 -0.000283067
+ 7.1e+09Hz 0.0132133 -0.000335081
+ 7.2e+09Hz 0.0132701 -0.000388427
+ 7.3e+09Hz 0.0133264 -0.000443086
+ 7.4e+09Hz 0.0133821 -0.000499036
+ 7.5e+09Hz 0.0134373 -0.000556257
+ 7.6e+09Hz 0.0134918 -0.000614726
+ 7.7e+09Hz 0.0135457 -0.000674421
+ 7.8e+09Hz 0.013599 -0.000735318
+ 7.9e+09Hz 0.0136516 -0.000797393
+ 8e+09Hz 0.0137034 -0.000860623
+ 8.1e+09Hz 0.0137545 -0.000924982
+ 8.2e+09Hz 0.0138049 -0.000990444
+ 8.3e+09Hz 0.0138544 -0.00105698
+ 8.4e+09Hz 0.0139032 -0.00112458
+ 8.5e+09Hz 0.0139511 -0.00119319
+ 8.6e+09Hz 0.0139982 -0.00126281
+ 8.7e+09Hz 0.0140445 -0.00133339
+ 8.8e+09Hz 0.0140898 -0.00140491
+ 8.9e+09Hz 0.0141343 -0.00147736
+ 9e+09Hz 0.0141778 -0.00155068
+ 9.1e+09Hz 0.0142205 -0.00162487
+ 9.2e+09Hz 0.0142622 -0.00169988
+ 9.3e+09Hz 0.0143029 -0.00177569
+ 9.4e+09Hz 0.0143427 -0.00185228
+ 9.5e+09Hz 0.0143814 -0.0019296
+ 9.6e+09Hz 0.0144193 -0.00200764
+ 9.7e+09Hz 0.0144561 -0.00208636
+ 9.8e+09Hz 0.0144919 -0.00216574
+ 9.9e+09Hz 0.0145267 -0.00224574
+ 1e+10Hz 0.0145604 -0.00232634
+ 1.01e+10Hz 0.0145932 -0.00240751
+ 1.02e+10Hz 0.0146249 -0.00248921
+ 1.03e+10Hz 0.0146556 -0.00257143
+ 1.04e+10Hz 0.0146853 -0.00265412
+ 1.05e+10Hz 0.0147139 -0.00273727
+ 1.06e+10Hz 0.0147415 -0.00282084
+ 1.07e+10Hz 0.014768 -0.00290481
+ 1.08e+10Hz 0.0147936 -0.00298915
+ 1.09e+10Hz 0.014818 -0.00307382
+ 1.1e+10Hz 0.0148415 -0.00315881
+ 1.11e+10Hz 0.0148639 -0.00324409
+ 1.12e+10Hz 0.0148853 -0.00332963
+ 1.13e+10Hz 0.0149056 -0.00341539
+ 1.14e+10Hz 0.014925 -0.00350137
+ 1.15e+10Hz 0.0149433 -0.00358753
+ 1.16e+10Hz 0.0149606 -0.00367385
+ 1.17e+10Hz 0.0149769 -0.0037603
+ 1.18e+10Hz 0.0149922 -0.00384686
+ 1.19e+10Hz 0.0150066 -0.0039335
+ 1.2e+10Hz 0.0150199 -0.0040202
+ 1.21e+10Hz 0.0150323 -0.00410694
+ 1.22e+10Hz 0.0150438 -0.0041937
+ 1.23e+10Hz 0.0150543 -0.00428046
+ 1.24e+10Hz 0.0150638 -0.00436719
+ 1.25e+10Hz 0.0150725 -0.00445387
+ 1.26e+10Hz 0.0150802 -0.00454048
+ 1.27e+10Hz 0.0150871 -0.00462701
+ 1.28e+10Hz 0.015093 -0.00471343
+ 1.29e+10Hz 0.0150981 -0.00479973
+ 1.3e+10Hz 0.0151023 -0.00488589
+ 1.31e+10Hz 0.0151057 -0.00497189
+ 1.32e+10Hz 0.0151083 -0.00505772
+ 1.33e+10Hz 0.01511 -0.00514336
+ 1.34e+10Hz 0.015111 -0.0052288
+ 1.35e+10Hz 0.0151112 -0.00531401
+ 1.36e+10Hz 0.0151106 -0.00539899
+ 1.37e+10Hz 0.0151093 -0.00548373
+ 1.38e+10Hz 0.0151072 -0.00556821
+ 1.39e+10Hz 0.0151044 -0.00565242
+ 1.4e+10Hz 0.0151009 -0.00573635
+ 1.41e+10Hz 0.0150968 -0.00581999
+ 1.42e+10Hz 0.015092 -0.00590332
+ 1.43e+10Hz 0.0150865 -0.00598635
+ 1.44e+10Hz 0.0150804 -0.00606906
+ 1.45e+10Hz 0.0150737 -0.00615144
+ 1.46e+10Hz 0.0150664 -0.00623349
+ 1.47e+10Hz 0.0150585 -0.0063152
+ 1.48e+10Hz 0.0150501 -0.00639657
+ 1.49e+10Hz 0.0150411 -0.00647758
+ 1.5e+10Hz 0.0150316 -0.00655824
+ 1.51e+10Hz 0.0150216 -0.00663855
+ 1.52e+10Hz 0.0150111 -0.00671849
+ 1.53e+10Hz 0.0150001 -0.00679806
+ 1.54e+10Hz 0.0149887 -0.00687728
+ 1.55e+10Hz 0.0149768 -0.00695612
+ 1.56e+10Hz 0.0149645 -0.0070346
+ 1.57e+10Hz 0.0149518 -0.00711271
+ 1.58e+10Hz 0.0149387 -0.00719045
+ 1.59e+10Hz 0.0149252 -0.00726782
+ 1.6e+10Hz 0.0149114 -0.00734483
+ 1.61e+10Hz 0.0148972 -0.00742148
+ 1.62e+10Hz 0.0148827 -0.00749777
+ 1.63e+10Hz 0.0148679 -0.0075737
+ 1.64e+10Hz 0.0148528 -0.00764927
+ 1.65e+10Hz 0.0148374 -0.0077245
+ 1.66e+10Hz 0.0148217 -0.00779938
+ 1.67e+10Hz 0.0148058 -0.00787392
+ 1.68e+10Hz 0.0147896 -0.00794813
+ 1.69e+10Hz 0.0147732 -0.00802201
+ 1.7e+10Hz 0.0147565 -0.00809556
+ 1.71e+10Hz 0.0147397 -0.0081688
+ 1.72e+10Hz 0.0147226 -0.00824173
+ 1.73e+10Hz 0.0147054 -0.00831436
+ 1.74e+10Hz 0.014688 -0.00838669
+ 1.75e+10Hz 0.0146704 -0.00845874
+ 1.76e+10Hz 0.0146527 -0.00853051
+ 1.77e+10Hz 0.0146348 -0.00860201
+ 1.78e+10Hz 0.0146168 -0.00867324
+ 1.79e+10Hz 0.0145986 -0.00874423
+ 1.8e+10Hz 0.0145803 -0.00881497
+ 1.81e+10Hz 0.0145619 -0.00888547
+ 1.82e+10Hz 0.0145434 -0.00895575
+ 1.83e+10Hz 0.0145248 -0.00902582
+ 1.84e+10Hz 0.0145061 -0.00909567
+ 1.85e+10Hz 0.0144873 -0.00916533
+ 1.86e+10Hz 0.0144684 -0.00923481
+ 1.87e+10Hz 0.0144494 -0.00930411
+ 1.88e+10Hz 0.0144303 -0.00937324
+ 1.89e+10Hz 0.0144112 -0.00944221
+ 1.9e+10Hz 0.014392 -0.00951104
+ 1.91e+10Hz 0.0143727 -0.00957973
+ 1.92e+10Hz 0.0143533 -0.00964829
+ 1.93e+10Hz 0.0143339 -0.00971673
+ 1.94e+10Hz 0.0143144 -0.00978506
+ 1.95e+10Hz 0.0142948 -0.0098533
+ 1.96e+10Hz 0.0142752 -0.00992144
+ 1.97e+10Hz 0.0142555 -0.00998951
+ 1.98e+10Hz 0.0142357 -0.0100575
+ 1.99e+10Hz 0.0142158 -0.0101254
+ 2e+10Hz 0.0141959 -0.0101933
+ 2.01e+10Hz 0.0141759 -0.0102612
+ 2.02e+10Hz 0.0141558 -0.0103289
+ 2.03e+10Hz 0.0141356 -0.0103967
+ 2.04e+10Hz 0.0141154 -0.0104645
+ 2.05e+10Hz 0.014095 -0.0105322
+ 2.06e+10Hz 0.0140746 -0.0105999
+ 2.07e+10Hz 0.0140541 -0.0106677
+ 2.08e+10Hz 0.0140335 -0.0107354
+ 2.09e+10Hz 0.0140127 -0.0108032
+ 2.1e+10Hz 0.0139919 -0.010871
+ 2.11e+10Hz 0.0139709 -0.0109388
+ 2.12e+10Hz 0.0139498 -0.0110066
+ 2.13e+10Hz 0.0139286 -0.0110745
+ 2.14e+10Hz 0.0139073 -0.0111425
+ 2.15e+10Hz 0.0138858 -0.0112105
+ 2.16e+10Hz 0.0138641 -0.0112785
+ 2.17e+10Hz 0.0138423 -0.0113466
+ 2.18e+10Hz 0.0138204 -0.0114148
+ 2.19e+10Hz 0.0137982 -0.011483
+ 2.2e+10Hz 0.0137759 -0.0115513
+ 2.21e+10Hz 0.0137534 -0.0116196
+ 2.22e+10Hz 0.0137308 -0.0116881
+ 2.23e+10Hz 0.0137079 -0.0117566
+ 2.24e+10Hz 0.0136848 -0.0118252
+ 2.25e+10Hz 0.0136615 -0.0118938
+ 2.26e+10Hz 0.013638 -0.0119626
+ 2.27e+10Hz 0.0136142 -0.0120314
+ 2.28e+10Hz 0.0135902 -0.0121003
+ 2.29e+10Hz 0.013566 -0.0121693
+ 2.3e+10Hz 0.0135415 -0.0122383
+ 2.31e+10Hz 0.0135168 -0.0123074
+ 2.32e+10Hz 0.0134918 -0.0123766
+ 2.33e+10Hz 0.0134665 -0.0124459
+ 2.34e+10Hz 0.0134409 -0.0125153
+ 2.35e+10Hz 0.013415 -0.0125847
+ 2.36e+10Hz 0.0133889 -0.0126542
+ 2.37e+10Hz 0.0133624 -0.0127237
+ 2.38e+10Hz 0.0133356 -0.0127933
+ 2.39e+10Hz 0.0133085 -0.012863
+ 2.4e+10Hz 0.0132811 -0.0129327
+ 2.41e+10Hz 0.0132533 -0.0130024
+ 2.42e+10Hz 0.0132252 -0.0130722
+ 2.43e+10Hz 0.0131968 -0.0131421
+ 2.44e+10Hz 0.013168 -0.0132119
+ 2.45e+10Hz 0.0131388 -0.0132818
+ 2.46e+10Hz 0.0131093 -0.0133517
+ 2.47e+10Hz 0.0130794 -0.0134217
+ 2.48e+10Hz 0.0130492 -0.0134916
+ 2.49e+10Hz 0.0130185 -0.0135615
+ 2.5e+10Hz 0.0129875 -0.0136315
+ 2.51e+10Hz 0.0129561 -0.0137014
+ 2.52e+10Hz 0.0129243 -0.0137713
+ 2.53e+10Hz 0.0128921 -0.0138412
+ 2.54e+10Hz 0.0128595 -0.013911
+ 2.55e+10Hz 0.0128266 -0.0139809
+ 2.56e+10Hz 0.0127932 -0.0140506
+ 2.57e+10Hz 0.0127594 -0.0141203
+ 2.58e+10Hz 0.0127251 -0.01419
+ 2.59e+10Hz 0.0126905 -0.0142595
+ 2.6e+10Hz 0.0126555 -0.014329
+ 2.61e+10Hz 0.01262 -0.0143984
+ 2.62e+10Hz 0.0125841 -0.0144677
+ 2.63e+10Hz 0.0125478 -0.0145369
+ 2.64e+10Hz 0.0125111 -0.014606
+ 2.65e+10Hz 0.012474 -0.014675
+ 2.66e+10Hz 0.0124365 -0.0147438
+ 2.67e+10Hz 0.0123985 -0.0148125
+ 2.68e+10Hz 0.0123601 -0.014881
+ 2.69e+10Hz 0.0123213 -0.0149494
+ 2.7e+10Hz 0.0122821 -0.0150177
+ 2.71e+10Hz 0.0122424 -0.0150857
+ 2.72e+10Hz 0.0122024 -0.0151536
+ 2.73e+10Hz 0.0121619 -0.0152213
+ 2.74e+10Hz 0.0121211 -0.0152888
+ 2.75e+10Hz 0.0120798 -0.0153561
+ 2.76e+10Hz 0.0120381 -0.0154232
+ 2.77e+10Hz 0.0119961 -0.01549
+ 2.78e+10Hz 0.0119536 -0.0155567
+ 2.79e+10Hz 0.0119108 -0.0156231
+ 2.8e+10Hz 0.0118675 -0.0156892
+ 2.81e+10Hz 0.0118239 -0.0157551
+ 2.82e+10Hz 0.0117799 -0.0158208
+ 2.83e+10Hz 0.0117355 -0.0158862
+ 2.84e+10Hz 0.0116908 -0.0159513
+ 2.85e+10Hz 0.0116456 -0.0160161
+ 2.86e+10Hz 0.0116002 -0.0160807
+ 2.87e+10Hz 0.0115544 -0.0161449
+ 2.88e+10Hz 0.0115082 -0.0162089
+ 2.89e+10Hz 0.0114617 -0.0162726
+ 2.9e+10Hz 0.0114148 -0.0163359
+ 2.91e+10Hz 0.0113677 -0.016399
+ 2.92e+10Hz 0.0113202 -0.0164617
+ 2.93e+10Hz 0.0112724 -0.0165241
+ 2.94e+10Hz 0.0112243 -0.0165862
+ 2.95e+10Hz 0.0111758 -0.0166479
+ 2.96e+10Hz 0.0111271 -0.0167094
+ 2.97e+10Hz 0.0110781 -0.0167704
+ 2.98e+10Hz 0.0110289 -0.0168312
+ 2.99e+10Hz 0.0109793 -0.0168916
+ 3e+10Hz 0.0109295 -0.0169516
+ 3.01e+10Hz 0.0108794 -0.0170113
+ 3.02e+10Hz 0.0108291 -0.0170706
+ 3.03e+10Hz 0.0107786 -0.0171296
+ 3.04e+10Hz 0.0107278 -0.0171882
+ 3.05e+10Hz 0.0106768 -0.0172464
+ 3.06e+10Hz 0.0106256 -0.0173043
+ 3.07e+10Hz 0.0105741 -0.0173619
+ 3.08e+10Hz 0.0105225 -0.017419
+ 3.09e+10Hz 0.0104707 -0.0174758
+ 3.1e+10Hz 0.0104186 -0.0175323
+ 3.11e+10Hz 0.0103664 -0.0175883
+ 3.12e+10Hz 0.0103141 -0.0176441
+ 3.13e+10Hz 0.0102615 -0.0176994
+ 3.14e+10Hz 0.0102089 -0.0177544
+ 3.15e+10Hz 0.010156 -0.017809
+ 3.16e+10Hz 0.0101031 -0.0178633
+ 3.17e+10Hz 0.0100499 -0.0179172
+ 3.18e+10Hz 0.00999672 -0.0179707
+ 3.19e+10Hz 0.00994337 -0.0180239
+ 3.2e+10Hz 0.00988991 -0.0180767
+ 3.21e+10Hz 0.00983634 -0.0181292
+ 3.22e+10Hz 0.00978268 -0.0181813
+ 3.23e+10Hz 0.00972892 -0.0182331
+ 3.24e+10Hz 0.00967508 -0.0182846
+ 3.25e+10Hz 0.00962116 -0.0183357
+ 3.26e+10Hz 0.00956717 -0.0183865
+ 3.27e+10Hz 0.00951311 -0.0184369
+ 3.28e+10Hz 0.00945899 -0.018487
+ 3.29e+10Hz 0.00940482 -0.0185368
+ 3.3e+10Hz 0.00935059 -0.0185863
+ 3.31e+10Hz 0.00929632 -0.0186355
+ 3.32e+10Hz 0.00924201 -0.0186843
+ 3.33e+10Hz 0.00918767 -0.0187328
+ 3.34e+10Hz 0.00913329 -0.0187811
+ 3.35e+10Hz 0.00907889 -0.018829
+ 3.36e+10Hz 0.00902446 -0.0188767
+ 3.37e+10Hz 0.00897002 -0.0189241
+ 3.38e+10Hz 0.00891556 -0.0189712
+ 3.39e+10Hz 0.00886109 -0.019018
+ 3.4e+10Hz 0.00880661 -0.0190645
+ 3.41e+10Hz 0.00875212 -0.0191108
+ 3.42e+10Hz 0.00869763 -0.0191568
+ 3.43e+10Hz 0.00864314 -0.0192026
+ 3.44e+10Hz 0.00858866 -0.0192481
+ 3.45e+10Hz 0.00853417 -0.0192934
+ 3.46e+10Hz 0.00847969 -0.0193385
+ 3.47e+10Hz 0.00842522 -0.0193833
+ 3.48e+10Hz 0.00837075 -0.0194279
+ 3.49e+10Hz 0.00831629 -0.0194723
+ 3.5e+10Hz 0.00826184 -0.0195165
+ 3.51e+10Hz 0.0082074 -0.0195604
+ 3.52e+10Hz 0.00815297 -0.0196042
+ 3.53e+10Hz 0.00809855 -0.0196477
+ 3.54e+10Hz 0.00804414 -0.0196911
+ 3.55e+10Hz 0.00798974 -0.0197343
+ 3.56e+10Hz 0.00793534 -0.0197773
+ 3.57e+10Hz 0.00788096 -0.0198201
+ 3.58e+10Hz 0.00782657 -0.0198628
+ 3.59e+10Hz 0.0077722 -0.0199053
+ 3.6e+10Hz 0.00771782 -0.0199476
+ 3.61e+10Hz 0.00766345 -0.0199898
+ 3.62e+10Hz 0.00760908 -0.0200319
+ 3.63e+10Hz 0.0075547 -0.0200737
+ 3.64e+10Hz 0.00750032 -0.0201155
+ 3.65e+10Hz 0.00744593 -0.0201571
+ 3.66e+10Hz 0.00739153 -0.0201986
+ 3.67e+10Hz 0.00733712 -0.0202399
+ 3.68e+10Hz 0.00728269 -0.0202812
+ 3.69e+10Hz 0.00722824 -0.0203223
+ 3.7e+10Hz 0.00717376 -0.0203633
+ 3.71e+10Hz 0.00711926 -0.0204041
+ 3.72e+10Hz 0.00706474 -0.0204449
+ 3.73e+10Hz 0.00701017 -0.0204856
+ 3.74e+10Hz 0.00695557 -0.0205261
+ 3.75e+10Hz 0.00690093 -0.0205666
+ 3.76e+10Hz 0.00684624 -0.0206069
+ 3.77e+10Hz 0.00679151 -0.0206471
+ 3.78e+10Hz 0.00673672 -0.0206873
+ 3.79e+10Hz 0.00668187 -0.0207274
+ 3.8e+10Hz 0.00662696 -0.0207673
+ 3.81e+10Hz 0.00657198 -0.0208072
+ 3.82e+10Hz 0.00651693 -0.020847
+ 3.83e+10Hz 0.00646181 -0.0208867
+ 3.84e+10Hz 0.00640661 -0.0209263
+ 3.85e+10Hz 0.00635132 -0.0209658
+ 3.86e+10Hz 0.00629594 -0.0210052
+ 3.87e+10Hz 0.00624047 -0.0210445
+ 3.88e+10Hz 0.0061849 -0.0210838
+ 3.89e+10Hz 0.00612923 -0.0211229
+ 3.9e+10Hz 0.00607346 -0.021162
+ 3.91e+10Hz 0.00601757 -0.0212009
+ 3.92e+10Hz 0.00596156 -0.0212398
+ 3.93e+10Hz 0.00590544 -0.0212786
+ 3.94e+10Hz 0.00584919 -0.0213173
+ 3.95e+10Hz 0.00579281 -0.0213559
+ 3.96e+10Hz 0.0057363 -0.0213944
+ 3.97e+10Hz 0.00567966 -0.0214328
+ 3.98e+10Hz 0.00562287 -0.021471
+ 3.99e+10Hz 0.00556594 -0.0215092
+ 4e+10Hz 0.00550886 -0.0215473
+ 4.01e+10Hz 0.00545163 -0.0215853
+ 4.02e+10Hz 0.00539424 -0.0216231
+ 4.03e+10Hz 0.0053367 -0.0216608
+ 4.04e+10Hz 0.00527899 -0.0216984
+ 4.05e+10Hz 0.00522112 -0.0217359
+ 4.06e+10Hz 0.00516308 -0.0217733
+ 4.07e+10Hz 0.00510487 -0.0218105
+ 4.08e+10Hz 0.00504649 -0.0218476
+ 4.09e+10Hz 0.00498792 -0.0218845
+ 4.1e+10Hz 0.00492919 -0.0219214
+ 4.11e+10Hz 0.00487026 -0.021958
+ 4.12e+10Hz 0.00481116 -0.0219945
+ 4.13e+10Hz 0.00475187 -0.0220309
+ 4.14e+10Hz 0.0046924 -0.0220671
+ 4.15e+10Hz 0.00463274 -0.0221031
+ 4.16e+10Hz 0.00457288 -0.0221389
+ 4.17e+10Hz 0.00451284 -0.0221746
+ 4.18e+10Hz 0.00445261 -0.0222101
+ 4.19e+10Hz 0.00439218 -0.0222454
+ 4.2e+10Hz 0.00433156 -0.0222805
+ 4.21e+10Hz 0.00427075 -0.0223155
+ 4.22e+10Hz 0.00420974 -0.0223502
+ 4.23e+10Hz 0.00414854 -0.0223847
+ 4.24e+10Hz 0.00408715 -0.022419
+ 4.25e+10Hz 0.00402556 -0.0224531
+ 4.26e+10Hz 0.00396378 -0.022487
+ 4.27e+10Hz 0.00390181 -0.0225206
+ 4.28e+10Hz 0.00383965 -0.022554
+ 4.29e+10Hz 0.0037773 -0.0225872
+ 4.3e+10Hz 0.00371476 -0.0226201
+ 4.31e+10Hz 0.00365204 -0.0226528
+ 4.32e+10Hz 0.00358913 -0.0226852
+ 4.33e+10Hz 0.00352604 -0.0227174
+ 4.34e+10Hz 0.00346276 -0.0227493
+ 4.35e+10Hz 0.00339931 -0.022781
+ 4.36e+10Hz 0.00333569 -0.0228123
+ 4.37e+10Hz 0.00327189 -0.0228434
+ 4.38e+10Hz 0.00320791 -0.0228742
+ 4.39e+10Hz 0.00314378 -0.0229048
+ 4.4e+10Hz 0.00307947 -0.022935
+ 4.41e+10Hz 0.00301501 -0.0229649
+ 4.42e+10Hz 0.00295039 -0.0229946
+ 4.43e+10Hz 0.00288562 -0.0230239
+ 4.44e+10Hz 0.00282069 -0.023053
+ 4.45e+10Hz 0.00275562 -0.0230817
+ 4.46e+10Hz 0.00269041 -0.0231101
+ 4.47e+10Hz 0.00262506 -0.0231382
+ 4.48e+10Hz 0.00255958 -0.0231659
+ 4.49e+10Hz 0.00249397 -0.0231934
+ 4.5e+10Hz 0.00242823 -0.0232205
+ 4.51e+10Hz 0.00236238 -0.0232472
+ 4.52e+10Hz 0.00229641 -0.0232737
+ 4.53e+10Hz 0.00223033 -0.0232998
+ 4.54e+10Hz 0.00216415 -0.0233255
+ 4.55e+10Hz 0.00209787 -0.0233509
+ 4.56e+10Hz 0.00203149 -0.023376
+ 4.57e+10Hz 0.00196503 -0.0234007
+ 4.58e+10Hz 0.00189848 -0.0234251
+ 4.59e+10Hz 0.00183186 -0.0234491
+ 4.6e+10Hz 0.00176516 -0.0234728
+ 4.61e+10Hz 0.00169839 -0.0234961
+ 4.62e+10Hz 0.00163157 -0.023519
+ 4.63e+10Hz 0.00156468 -0.0235416
+ 4.64e+10Hz 0.00149775 -0.0235638
+ 4.65e+10Hz 0.00143078 -0.0235857
+ 4.66e+10Hz 0.00136376 -0.0236072
+ 4.67e+10Hz 0.00129671 -0.0236284
+ 4.68e+10Hz 0.00122964 -0.0236492
+ 4.69e+10Hz 0.00116254 -0.0236696
+ 4.7e+10Hz 0.00109543 -0.0236897
+ 4.71e+10Hz 0.0010283 -0.0237094
+ 4.72e+10Hz 0.000961174 -0.0237287
+ 4.73e+10Hz 0.000894047 -0.0237477
+ 4.74e+10Hz 0.000826927 -0.0237664
+ 4.75e+10Hz 0.000759819 -0.0237846
+ 4.76e+10Hz 0.000692728 -0.0238026
+ 4.77e+10Hz 0.00062566 -0.0238201
+ 4.78e+10Hz 0.000558621 -0.0238373
+ 4.79e+10Hz 0.000491615 -0.0238542
+ 4.8e+10Hz 0.000424648 -0.0238707
+ 4.81e+10Hz 0.000357726 -0.0238869
+ 4.82e+10Hz 0.000290852 -0.0239027
+ 4.83e+10Hz 0.000224033 -0.0239181
+ 4.84e+10Hz 0.000157272 -0.0239333
+ 4.85e+10Hz 9.05754e-05 -0.0239481
+ 4.86e+10Hz 2.39469e-05 -0.0239625
+ 4.87e+10Hz -4.26085e-05 -0.0239766
+ 4.88e+10Hz -0.000109087 -0.0239904
+ 4.89e+10Hz -0.000175483 -0.0240039
+ 4.9e+10Hz -0.000241793 -0.024017
+ 4.91e+10Hz -0.000308014 -0.0240299
+ 4.92e+10Hz -0.00037414 -0.0240424
+ 4.93e+10Hz -0.000440169 -0.0240546
+ 4.94e+10Hz -0.000506097 -0.0240664
+ 4.95e+10Hz -0.000571919 -0.024078
+ 4.96e+10Hz -0.000637633 -0.0240893
+ 4.97e+10Hz -0.000703235 -0.0241003
+ 4.98e+10Hz -0.000768723 -0.0241109
+ 4.99e+10Hz -0.000834093 -0.0241213
+ 5e+10Hz -0.000899342 -0.0241314
+ 5.01e+10Hz -0.000964469 -0.0241412
+ 5.02e+10Hz -0.00102947 -0.0241508
+ 5.03e+10Hz -0.00109434 -0.02416
+ 5.04e+10Hz -0.00115908 -0.024169
+ 5.05e+10Hz -0.00122369 -0.0241778
+ 5.06e+10Hz -0.00128817 -0.0241862
+ 5.07e+10Hz -0.00135251 -0.0241944
+ 5.08e+10Hz -0.00141671 -0.0242024
+ 5.09e+10Hz -0.00148078 -0.0242101
+ 5.1e+10Hz -0.0015447 -0.0242175
+ 5.11e+10Hz -0.00160848 -0.0242247
+ 5.12e+10Hz -0.00167212 -0.0242317
+ 5.13e+10Hz -0.00173562 -0.0242385
+ 5.14e+10Hz -0.00179897 -0.024245
+ 5.15e+10Hz -0.00186218 -0.0242513
+ 5.16e+10Hz -0.00192525 -0.0242574
+ 5.17e+10Hz -0.00198817 -0.0242632
+ 5.18e+10Hz -0.00205094 -0.0242689
+ 5.19e+10Hz -0.00211357 -0.0242743
+ 5.2e+10Hz -0.00217606 -0.0242795
+ 5.21e+10Hz -0.00223839 -0.0242846
+ 5.22e+10Hz -0.00230059 -0.0242894
+ 5.23e+10Hz -0.00236264 -0.0242941
+ 5.24e+10Hz -0.00242455 -0.0242985
+ 5.25e+10Hz -0.00248632 -0.0243028
+ 5.26e+10Hz -0.00254795 -0.0243069
+ 5.27e+10Hz -0.00260943 -0.0243108
+ 5.28e+10Hz -0.00267078 -0.0243145
+ 5.29e+10Hz -0.00273198 -0.0243181
+ 5.3e+10Hz -0.00279306 -0.0243215
+ 5.31e+10Hz -0.00285399 -0.0243247
+ 5.32e+10Hz -0.00291479 -0.0243278
+ 5.33e+10Hz -0.00297546 -0.0243307
+ 5.34e+10Hz -0.003036 -0.0243334
+ 5.35e+10Hz -0.00309641 -0.024336
+ 5.36e+10Hz -0.00315669 -0.0243384
+ 5.37e+10Hz -0.00321685 -0.0243407
+ 5.38e+10Hz -0.00327688 -0.0243428
+ 5.39e+10Hz -0.00333679 -0.0243448
+ 5.4e+10Hz -0.00339658 -0.0243467
+ 5.41e+10Hz -0.00345625 -0.0243484
+ 5.42e+10Hz -0.00351581 -0.0243499
+ 5.43e+10Hz -0.00357525 -0.0243514
+ 5.44e+10Hz -0.00363458 -0.0243526
+ 5.45e+10Hz -0.0036938 -0.0243538
+ 5.46e+10Hz -0.00375291 -0.0243548
+ 5.47e+10Hz -0.00381192 -0.0243557
+ 5.48e+10Hz -0.00387082 -0.0243564
+ 5.49e+10Hz -0.00392962 -0.024357
+ 5.5e+10Hz -0.00398832 -0.0243575
+ 5.51e+10Hz -0.00404693 -0.0243578
+ 5.52e+10Hz -0.00410543 -0.0243581
+ 5.53e+10Hz -0.00416385 -0.0243581
+ 5.54e+10Hz -0.00422217 -0.0243581
+ 5.55e+10Hz -0.0042804 -0.0243579
+ 5.56e+10Hz -0.00433854 -0.0243576
+ 5.57e+10Hz -0.0043966 -0.0243572
+ 5.58e+10Hz -0.00445457 -0.0243566
+ 5.59e+10Hz -0.00451246 -0.0243559
+ 5.6e+10Hz -0.00457027 -0.024355
+ 5.61e+10Hz -0.004628 -0.0243541
+ 5.62e+10Hz -0.00468565 -0.024353
+ 5.63e+10Hz -0.00474323 -0.0243517
+ 5.64e+10Hz -0.00480073 -0.0243504
+ 5.65e+10Hz -0.00485815 -0.0243489
+ 5.66e+10Hz -0.0049155 -0.0243472
+ 5.67e+10Hz -0.00497278 -0.0243454
+ 5.68e+10Hz -0.00502999 -0.0243435
+ 5.69e+10Hz -0.00508713 -0.0243415
+ 5.7e+10Hz -0.0051442 -0.0243393
+ 5.71e+10Hz -0.0052012 -0.0243369
+ 5.72e+10Hz -0.00525814 -0.0243344
+ 5.73e+10Hz -0.005315 -0.0243318
+ 5.74e+10Hz -0.0053718 -0.024329
+ 5.75e+10Hz -0.00542854 -0.0243261
+ 5.76e+10Hz -0.0054852 -0.024323
+ 5.77e+10Hz -0.0055418 -0.0243198
+ 5.78e+10Hz -0.00559834 -0.0243164
+ 5.79e+10Hz -0.0056548 -0.0243129
+ 5.8e+10Hz -0.00571121 -0.0243092
+ 5.81e+10Hz -0.00576754 -0.0243054
+ 5.82e+10Hz -0.00582381 -0.0243014
+ 5.83e+10Hz -0.00588 -0.0242972
+ 5.84e+10Hz -0.00593613 -0.0242929
+ 5.85e+10Hz -0.00599219 -0.0242884
+ 5.86e+10Hz -0.00604818 -0.0242837
+ 5.87e+10Hz -0.0061041 -0.0242789
+ 5.88e+10Hz -0.00615994 -0.0242739
+ 5.89e+10Hz -0.00621571 -0.0242687
+ 5.9e+10Hz -0.0062714 -0.0242634
+ 5.91e+10Hz -0.00632702 -0.0242578
+ 5.92e+10Hz -0.00638256 -0.0242522
+ 5.93e+10Hz -0.00643801 -0.0242463
+ 5.94e+10Hz -0.00649339 -0.0242402
+ 5.95e+10Hz -0.00654868 -0.024234
+ 5.96e+10Hz -0.00660388 -0.0242276
+ 5.97e+10Hz -0.006659 -0.024221
+ 5.98e+10Hz -0.00671402 -0.0242143
+ 5.99e+10Hz -0.00676896 -0.0242073
+ 6e+10Hz -0.00682379 -0.0242002
+ 6.01e+10Hz -0.00687853 -0.0241929
+ 6.02e+10Hz -0.00693317 -0.0241854
+ 6.03e+10Hz -0.00698771 -0.0241777
+ 6.04e+10Hz -0.00704214 -0.0241698
+ 6.05e+10Hz -0.00709647 -0.0241617
+ 6.06e+10Hz -0.00715068 -0.0241535
+ 6.07e+10Hz -0.00720478 -0.024145
+ 6.08e+10Hz -0.00725876 -0.0241364
+ 6.09e+10Hz -0.00731262 -0.0241276
+ 6.1e+10Hz -0.00736636 -0.0241186
+ 6.11e+10Hz -0.00741997 -0.0241094
+ 6.12e+10Hz -0.00747345 -0.0241
+ 6.13e+10Hz -0.0075268 -0.0240904
+ 6.14e+10Hz -0.00758002 -0.0240806
+ 6.15e+10Hz -0.00763309 -0.0240707
+ 6.16e+10Hz -0.00768603 -0.0240606
+ 6.17e+10Hz -0.00773881 -0.0240502
+ 6.18e+10Hz -0.00779145 -0.0240398
+ 6.19e+10Hz -0.00784394 -0.0240291
+ 6.2e+10Hz -0.00789627 -0.0240182
+ 6.21e+10Hz -0.00794845 -0.0240072
+ 6.22e+10Hz -0.00800046 -0.0239959
+ 6.23e+10Hz -0.00805231 -0.0239846
+ 6.24e+10Hz -0.00810399 -0.023973
+ 6.25e+10Hz -0.00815549 -0.0239612
+ 6.26e+10Hz -0.00820683 -0.0239493
+ 6.27e+10Hz -0.00825798 -0.0239372
+ 6.28e+10Hz -0.00830896 -0.023925
+ 6.29e+10Hz -0.00835975 -0.0239126
+ 6.3e+10Hz -0.00841035 -0.0239
+ 6.31e+10Hz -0.00846076 -0.0238873
+ 6.32e+10Hz -0.00851098 -0.0238744
+ 6.33e+10Hz -0.00856101 -0.0238613
+ 6.34e+10Hz -0.00861083 -0.0238481
+ 6.35e+10Hz -0.00866046 -0.0238348
+ 6.36e+10Hz -0.00870988 -0.0238213
+ 6.37e+10Hz -0.00875909 -0.0238077
+ 6.38e+10Hz -0.0088081 -0.0237939
+ 6.39e+10Hz -0.00885689 -0.02378
+ 6.4e+10Hz -0.00890547 -0.023766
+ 6.41e+10Hz -0.00895384 -0.0237519
+ 6.42e+10Hz -0.00900199 -0.0237376
+ 6.43e+10Hz -0.00904991 -0.0237232
+ 6.44e+10Hz -0.00909762 -0.0237087
+ 6.45e+10Hz -0.0091451 -0.0236941
+ 6.46e+10Hz -0.00919235 -0.0236793
+ 6.47e+10Hz -0.00923938 -0.0236645
+ 6.48e+10Hz -0.00928618 -0.0236496
+ 6.49e+10Hz -0.00933276 -0.0236346
+ 6.5e+10Hz -0.0093791 -0.0236194
+ 6.51e+10Hz -0.0094252 -0.0236043
+ 6.52e+10Hz -0.00947108 -0.023589
+ 6.53e+10Hz -0.00951672 -0.0235736
+ 6.54e+10Hz -0.00956213 -0.0235582
+ 6.55e+10Hz -0.0096073 -0.0235427
+ 6.56e+10Hz -0.00965224 -0.0235272
+ 6.57e+10Hz -0.00969694 -0.0235115
+ 6.58e+10Hz -0.00974141 -0.0234959
+ 6.59e+10Hz -0.00978564 -0.0234802
+ 6.6e+10Hz -0.00982963 -0.0234644
+ 6.61e+10Hz -0.00987339 -0.0234486
+ 6.62e+10Hz -0.00991692 -0.0234328
+ 6.63e+10Hz -0.00996021 -0.0234169
+ 6.64e+10Hz -0.0100033 -0.0234011
+ 6.65e+10Hz -0.0100461 -0.0233852
+ 6.66e+10Hz -0.0100887 -0.0233692
+ 6.67e+10Hz -0.010131 -0.0233533
+ 6.68e+10Hz -0.0101732 -0.0233374
+ 6.69e+10Hz -0.0102151 -0.0233214
+ 6.7e+10Hz -0.0102567 -0.0233055
+ 6.71e+10Hz -0.0102982 -0.0232896
+ 6.72e+10Hz -0.0103394 -0.0232737
+ 6.73e+10Hz -0.0103804 -0.0232578
+ 6.74e+10Hz -0.0104212 -0.0232419
+ 6.75e+10Hz -0.0104618 -0.023226
+ 6.76e+10Hz -0.0105021 -0.0232102
+ 6.77e+10Hz -0.0105423 -0.0231944
+ 6.78e+10Hz -0.0105822 -0.0231786
+ 6.79e+10Hz -0.0106219 -0.0231629
+ 6.8e+10Hz -0.0106615 -0.0231473
+ 6.81e+10Hz -0.0107008 -0.0231316
+ 6.82e+10Hz -0.0107399 -0.0231161
+ 6.83e+10Hz -0.0107788 -0.0231006
+ 6.84e+10Hz -0.0108175 -0.0230851
+ 6.85e+10Hz -0.0108561 -0.0230697
+ 6.86e+10Hz -0.0108944 -0.0230544
+ 6.87e+10Hz -0.0109326 -0.0230391
+ 6.88e+10Hz -0.0109706 -0.023024
+ 6.89e+10Hz -0.0110084 -0.0230089
+ 6.9e+10Hz -0.011046 -0.0229938
+ 6.91e+10Hz -0.0110835 -0.0229789
+ 6.92e+10Hz -0.0111208 -0.022964
+ 6.93e+10Hz -0.0111579 -0.0229493
+ 6.94e+10Hz -0.0111949 -0.0229346
+ 6.95e+10Hz -0.0112317 -0.02292
+ 6.96e+10Hz -0.0112684 -0.0229055
+ 6.97e+10Hz -0.011305 -0.0228911
+ 6.98e+10Hz -0.0113414 -0.0228768
+ 6.99e+10Hz -0.0113776 -0.0228626
+ 7e+10Hz -0.0114137 -0.0228485
+ 7.01e+10Hz -0.0114497 -0.0228345
+ 7.02e+10Hz -0.0114856 -0.0228206
+ 7.03e+10Hz -0.0115213 -0.0228068
+ 7.04e+10Hz -0.011557 -0.0227931
+ 7.05e+10Hz -0.0115925 -0.0227795
+ 7.06e+10Hz -0.0116279 -0.022766
+ 7.07e+10Hz -0.0116632 -0.0227527
+ 7.08e+10Hz -0.0116984 -0.0227394
+ 7.09e+10Hz -0.0117335 -0.0227263
+ 7.1e+10Hz -0.0117685 -0.0227133
+ 7.11e+10Hz -0.0118035 -0.0227004
+ 7.12e+10Hz -0.0118383 -0.0226875
+ 7.13e+10Hz -0.0118731 -0.0226749
+ 7.14e+10Hz -0.0119077 -0.0226623
+ 7.15e+10Hz -0.0119424 -0.0226498
+ 7.16e+10Hz -0.0119769 -0.0226374
+ 7.17e+10Hz -0.0120114 -0.0226252
+ 7.18e+10Hz -0.0120458 -0.0226131
+ 7.19e+10Hz -0.0120802 -0.022601
+ 7.2e+10Hz -0.0121145 -0.0225891
+ 7.21e+10Hz -0.0121488 -0.0225773
+ 7.22e+10Hz -0.012183 -0.0225656
+ 7.23e+10Hz -0.0122172 -0.022554
+ 7.24e+10Hz -0.0122513 -0.0225425
+ 7.25e+10Hz -0.0122854 -0.0225311
+ 7.26e+10Hz -0.0123195 -0.0225198
+ 7.27e+10Hz -0.0123535 -0.0225086
+ 7.28e+10Hz -0.0123875 -0.0224976
+ 7.29e+10Hz -0.0124215 -0.0224866
+ 7.3e+10Hz -0.0124555 -0.0224757
+ 7.31e+10Hz -0.0124894 -0.0224649
+ 7.32e+10Hz -0.0125234 -0.0224542
+ 7.33e+10Hz -0.0125573 -0.0224436
+ 7.34e+10Hz -0.0125912 -0.0224331
+ 7.35e+10Hz -0.0126251 -0.0224226
+ 7.36e+10Hz -0.0126591 -0.0224123
+ 7.37e+10Hz -0.012693 -0.022402
+ 7.38e+10Hz -0.0127269 -0.0223919
+ 7.39e+10Hz -0.0127608 -0.0223818
+ 7.4e+10Hz -0.0127947 -0.0223717
+ 7.41e+10Hz -0.0128286 -0.0223618
+ 7.42e+10Hz -0.0128626 -0.0223519
+ 7.43e+10Hz -0.0128965 -0.0223421
+ 7.44e+10Hz -0.0129304 -0.0223324
+ 7.45e+10Hz -0.0129644 -0.0223228
+ 7.46e+10Hz -0.0129984 -0.0223132
+ 7.47e+10Hz -0.0130324 -0.0223036
+ 7.48e+10Hz -0.0130664 -0.0222942
+ 7.49e+10Hz -0.0131004 -0.0222848
+ 7.5e+10Hz -0.0131345 -0.0222754
+ 7.51e+10Hz -0.0131685 -0.0222662
+ 7.52e+10Hz -0.0132026 -0.0222569
+ 7.53e+10Hz -0.0132367 -0.0222477
+ 7.54e+10Hz -0.0132708 -0.0222386
+ 7.55e+10Hz -0.013305 -0.0222295
+ 7.56e+10Hz -0.0133392 -0.0222205
+ 7.57e+10Hz -0.0133734 -0.0222115
+ 7.58e+10Hz -0.0134076 -0.0222026
+ 7.59e+10Hz -0.0134418 -0.0221937
+ 7.6e+10Hz -0.0134761 -0.0221848
+ 7.61e+10Hz -0.0135104 -0.022176
+ 7.62e+10Hz -0.0135447 -0.0221672
+ 7.63e+10Hz -0.013579 -0.0221584
+ 7.64e+10Hz -0.0136134 -0.0221497
+ 7.65e+10Hz -0.0136477 -0.022141
+ 7.66e+10Hz -0.0136821 -0.0221324
+ 7.67e+10Hz -0.0137166 -0.0221237
+ 7.68e+10Hz -0.013751 -0.0221151
+ 7.69e+10Hz -0.0137855 -0.0221066
+ 7.7e+10Hz -0.01382 -0.022098
+ 7.71e+10Hz -0.0138545 -0.0220895
+ 7.72e+10Hz -0.013889 -0.022081
+ 7.73e+10Hz -0.0139236 -0.0220726
+ 7.74e+10Hz -0.0139581 -0.0220642
+ 7.75e+10Hz -0.0139927 -0.0220557
+ 7.76e+10Hz -0.0140273 -0.0220474
+ 7.77e+10Hz -0.0140619 -0.022039
+ 7.78e+10Hz -0.0140966 -0.0220307
+ 7.79e+10Hz -0.0141312 -0.0220224
+ 7.8e+10Hz -0.0141659 -0.0220141
+ 7.81e+10Hz -0.0142006 -0.0220058
+ 7.82e+10Hz -0.0142353 -0.0219976
+ 7.83e+10Hz -0.01427 -0.0219893
+ 7.84e+10Hz -0.0143047 -0.0219812
+ 7.85e+10Hz -0.0143394 -0.021973
+ 7.86e+10Hz -0.0143742 -0.0219648
+ 7.87e+10Hz -0.0144089 -0.0219567
+ 7.88e+10Hz -0.0144437 -0.0219486
+ 7.89e+10Hz -0.0144785 -0.0219406
+ 7.9e+10Hz -0.0145133 -0.0219326
+ 7.91e+10Hz -0.0145481 -0.0219246
+ 7.92e+10Hz -0.0145829 -0.0219166
+ 7.93e+10Hz -0.0146177 -0.0219087
+ 7.94e+10Hz -0.0146525 -0.0219008
+ 7.95e+10Hz -0.0146874 -0.0218929
+ 7.96e+10Hz -0.0147222 -0.0218851
+ 7.97e+10Hz -0.0147571 -0.0218773
+ 7.98e+10Hz -0.014792 -0.0218695
+ 7.99e+10Hz -0.0148268 -0.0218618
+ 8e+10Hz -0.0148617 -0.0218542
+ 8.01e+10Hz -0.0148966 -0.0218465
+ 8.02e+10Hz -0.0149315 -0.021839
+ 8.03e+10Hz -0.0149665 -0.0218315
+ 8.04e+10Hz -0.0150014 -0.021824
+ 8.05e+10Hz -0.0150363 -0.0218166
+ 8.06e+10Hz -0.0150713 -0.0218092
+ 8.07e+10Hz -0.0151063 -0.0218019
+ 8.08e+10Hz -0.0151413 -0.0217946
+ 8.09e+10Hz -0.0151763 -0.0217874
+ 8.1e+10Hz -0.0152114 -0.0217803
+ 8.11e+10Hz -0.0152464 -0.0217732
+ 8.12e+10Hz -0.0152815 -0.0217663
+ 8.13e+10Hz -0.0153166 -0.0217593
+ 8.14e+10Hz -0.0153518 -0.0217525
+ 8.15e+10Hz -0.0153869 -0.0217457
+ 8.16e+10Hz -0.0154221 -0.021739
+ 8.17e+10Hz -0.0154574 -0.0217324
+ 8.18e+10Hz -0.0154926 -0.0217258
+ 8.19e+10Hz -0.0155279 -0.0217193
+ 8.2e+10Hz -0.0155633 -0.021713
+ 8.21e+10Hz -0.0155987 -0.0217067
+ 8.22e+10Hz -0.0156341 -0.0217005
+ 8.23e+10Hz -0.0156696 -0.0216943
+ 8.24e+10Hz -0.0157052 -0.0216883
+ 8.25e+10Hz -0.0157408 -0.0216824
+ 8.26e+10Hz -0.0157765 -0.0216766
+ 8.27e+10Hz -0.0158122 -0.0216708
+ 8.28e+10Hz -0.015848 -0.0216652
+ 8.29e+10Hz -0.0158839 -0.0216596
+ 8.3e+10Hz -0.0159198 -0.0216542
+ 8.31e+10Hz -0.0159559 -0.0216489
+ 8.32e+10Hz -0.015992 -0.0216436
+ 8.33e+10Hz -0.0160282 -0.0216385
+ 8.34e+10Hz -0.0160645 -0.0216335
+ 8.35e+10Hz -0.0161009 -0.0216286
+ 8.36e+10Hz -0.0161374 -0.0216238
+ 8.37e+10Hz -0.0161741 -0.0216191
+ 8.38e+10Hz -0.0162108 -0.0216146
+ 8.39e+10Hz -0.0162476 -0.0216101
+ 8.4e+10Hz -0.0162846 -0.0216057
+ 8.41e+10Hz -0.0163217 -0.0216015
+ 8.42e+10Hz -0.016359 -0.0215974
+ 8.43e+10Hz -0.0163963 -0.0215934
+ 8.44e+10Hz -0.0164339 -0.0215894
+ 8.45e+10Hz -0.0164716 -0.0215857
+ 8.46e+10Hz -0.0165094 -0.021582
+ 8.47e+10Hz -0.0165474 -0.0215784
+ 8.48e+10Hz -0.0165856 -0.0215749
+ 8.49e+10Hz -0.0166239 -0.0215716
+ 8.5e+10Hz -0.0166625 -0.0215683
+ 8.51e+10Hz -0.0167012 -0.0215652
+ 8.52e+10Hz -0.0167401 -0.0215622
+ 8.53e+10Hz -0.0167792 -0.0215592
+ 8.54e+10Hz -0.0168185 -0.0215564
+ 8.55e+10Hz -0.016858 -0.0215537
+ 8.56e+10Hz -0.0168978 -0.021551
+ 8.57e+10Hz -0.0169378 -0.0215485
+ 8.58e+10Hz -0.016978 -0.021546
+ 8.59e+10Hz -0.0170184 -0.0215437
+ 8.6e+10Hz -0.0170591 -0.0215414
+ 8.61e+10Hz -0.0171 -0.0215392
+ 8.62e+10Hz -0.0171412 -0.0215371
+ 8.63e+10Hz -0.0171827 -0.0215351
+ 8.64e+10Hz -0.0172244 -0.0215331
+ 8.65e+10Hz -0.0172664 -0.0215312
+ 8.66e+10Hz -0.0173087 -0.0215294
+ 8.67e+10Hz -0.0173512 -0.0215276
+ 8.68e+10Hz -0.0173941 -0.0215259
+ 8.69e+10Hz -0.0174373 -0.0215242
+ 8.7e+10Hz -0.0174807 -0.0215226
+ 8.71e+10Hz -0.0175245 -0.021521
+ 8.72e+10Hz -0.0175686 -0.0215194
+ 8.73e+10Hz -0.017613 -0.0215179
+ 8.74e+10Hz -0.0176578 -0.0215164
+ 8.75e+10Hz -0.0177029 -0.0215149
+ 8.76e+10Hz -0.0177483 -0.0215134
+ 8.77e+10Hz -0.0177941 -0.0215119
+ 8.78e+10Hz -0.0178402 -0.0215104
+ 8.79e+10Hz -0.0178867 -0.0215089
+ 8.8e+10Hz -0.0179335 -0.0215074
+ 8.81e+10Hz -0.0179807 -0.0215059
+ 8.82e+10Hz -0.0180283 -0.0215043
+ 8.83e+10Hz -0.0180762 -0.0215027
+ 8.84e+10Hz -0.0181246 -0.0215011
+ 8.85e+10Hz -0.0181733 -0.0214994
+ 8.86e+10Hz -0.0182224 -0.0214976
+ 8.87e+10Hz -0.0182719 -0.0214957
+ 8.88e+10Hz -0.0183218 -0.0214938
+ 8.89e+10Hz -0.0183721 -0.0214918
+ 8.9e+10Hz -0.0184228 -0.0214897
+ 8.91e+10Hz -0.0184739 -0.0214875
+ 8.92e+10Hz -0.0185254 -0.0214851
+ 8.93e+10Hz -0.0185773 -0.0214827
+ 8.94e+10Hz -0.0186297 -0.0214801
+ 8.95e+10Hz -0.0186824 -0.0214773
+ 8.96e+10Hz -0.0187356 -0.0214744
+ 8.97e+10Hz -0.0187892 -0.0214714
+ 8.98e+10Hz -0.0188432 -0.0214682
+ 8.99e+10Hz -0.0188977 -0.0214648
+ 9e+10Hz -0.0189526 -0.0214612
+ 9.01e+10Hz -0.0190079 -0.0214574
+ 9.02e+10Hz -0.0190636 -0.0214533
+ 9.03e+10Hz -0.0191198 -0.0214491
+ 9.04e+10Hz -0.0191764 -0.0214446
+ 9.05e+10Hz -0.0192335 -0.0214399
+ 9.06e+10Hz -0.0192909 -0.0214349
+ 9.07e+10Hz -0.0193488 -0.0214297
+ 9.08e+10Hz -0.0194071 -0.0214242
+ 9.09e+10Hz -0.0194659 -0.0214184
+ 9.1e+10Hz -0.0195251 -0.0214123
+ 9.11e+10Hz -0.0195847 -0.0214059
+ 9.12e+10Hz -0.0196447 -0.0213991
+ 9.13e+10Hz -0.0197052 -0.0213921
+ 9.14e+10Hz -0.0197661 -0.0213847
+ 9.15e+10Hz -0.0198274 -0.0213769
+ 9.16e+10Hz -0.0198891 -0.0213688
+ 9.17e+10Hz -0.0199512 -0.0213603
+ 9.18e+10Hz -0.0200138 -0.0213515
+ 9.19e+10Hz -0.0200767 -0.0213422
+ 9.2e+10Hz -0.0201401 -0.0213325
+ 9.21e+10Hz -0.0202038 -0.0213225
+ 9.22e+10Hz -0.020268 -0.0213119
+ 9.23e+10Hz -0.0203325 -0.021301
+ 9.24e+10Hz -0.0203974 -0.0212896
+ 9.25e+10Hz -0.0204627 -0.0212778
+ 9.26e+10Hz -0.0205284 -0.0212654
+ 9.27e+10Hz -0.0205945 -0.0212526
+ 9.28e+10Hz -0.0206609 -0.0212393
+ 9.29e+10Hz -0.0207277 -0.0212255
+ 9.3e+10Hz -0.0207948 -0.0212112
+ 9.31e+10Hz -0.0208623 -0.0211964
+ 9.32e+10Hz -0.0209301 -0.0211811
+ 9.33e+10Hz -0.0209983 -0.0211652
+ 9.34e+10Hz -0.0210667 -0.0211487
+ 9.35e+10Hz -0.0211355 -0.0211318
+ 9.36e+10Hz -0.0212046 -0.0211142
+ 9.37e+10Hz -0.021274 -0.021096
+ 9.38e+10Hz -0.0213437 -0.0210773
+ 9.39e+10Hz -0.0214137 -0.021058
+ 9.4e+10Hz -0.021484 -0.0210381
+ 9.41e+10Hz -0.0215545 -0.0210175
+ 9.42e+10Hz -0.0216253 -0.0209964
+ 9.43e+10Hz -0.0216963 -0.0209746
+ 9.44e+10Hz -0.0217676 -0.0209522
+ 9.45e+10Hz -0.0218391 -0.0209291
+ 9.46e+10Hz -0.0219108 -0.0209054
+ 9.47e+10Hz -0.0219828 -0.020881
+ 9.48e+10Hz -0.0220549 -0.020856
+ 9.49e+10Hz -0.0221272 -0.0208303
+ 9.5e+10Hz -0.0221997 -0.0208039
+ 9.51e+10Hz -0.0222724 -0.0207768
+ 9.52e+10Hz -0.0223452 -0.0207491
+ 9.53e+10Hz -0.0224182 -0.0207206
+ 9.54e+10Hz -0.0224913 -0.0206914
+ 9.55e+10Hz -0.0225646 -0.0206615
+ 9.56e+10Hz -0.0226379 -0.0206309
+ 9.57e+10Hz -0.0227114 -0.0205996
+ 9.58e+10Hz -0.0227849 -0.0205676
+ 9.59e+10Hz -0.0228585 -0.0205348
+ 9.6e+10Hz -0.0229322 -0.0205013
+ 9.61e+10Hz -0.0230059 -0.0204671
+ 9.62e+10Hz -0.0230797 -0.0204321
+ 9.63e+10Hz -0.0231535 -0.0203963
+ 9.64e+10Hz -0.0232273 -0.0203599
+ 9.65e+10Hz -0.0233012 -0.0203226
+ 9.66e+10Hz -0.023375 -0.0202846
+ 9.67e+10Hz -0.0234488 -0.0202459
+ 9.68e+10Hz -0.0235225 -0.0202064
+ 9.69e+10Hz -0.0235962 -0.0201661
+ 9.7e+10Hz -0.0236699 -0.0201251
+ 9.71e+10Hz -0.0237434 -0.0200833
+ 9.72e+10Hz -0.0238169 -0.0200408
+ 9.73e+10Hz -0.0238903 -0.0199974
+ 9.74e+10Hz -0.0239636 -0.0199533
+ 9.75e+10Hz -0.0240367 -0.0199085
+ 9.76e+10Hz -0.0241097 -0.0198629
+ 9.77e+10Hz -0.0241826 -0.0198165
+ 9.78e+10Hz -0.0242553 -0.0197693
+ 9.79e+10Hz -0.0243278 -0.0197214
+ 9.8e+10Hz -0.0244002 -0.0196727
+ 9.81e+10Hz -0.0244723 -0.0196232
+ 9.82e+10Hz -0.0245442 -0.019573
+ 9.83e+10Hz -0.0246159 -0.0195221
+ 9.84e+10Hz -0.0246873 -0.0194703
+ 9.85e+10Hz -0.0247585 -0.0194178
+ 9.86e+10Hz -0.0248294 -0.0193646
+ 9.87e+10Hz -0.0249001 -0.0193106
+ 9.88e+10Hz -0.0249704 -0.0192559
+ 9.89e+10Hz -0.0250405 -0.0192004
+ 9.9e+10Hz -0.0251102 -0.0191442
+ 9.91e+10Hz -0.0251796 -0.0190872
+ 9.92e+10Hz -0.0252487 -0.0190296
+ 9.93e+10Hz -0.0253174 -0.0189712
+ 9.94e+10Hz -0.0253858 -0.018912
+ 9.95e+10Hz -0.0254537 -0.0188522
+ 9.96e+10Hz -0.0255213 -0.0187916
+ 9.97e+10Hz -0.0255885 -0.0187304
+ 9.98e+10Hz -0.0256553 -0.0186684
+ 9.99e+10Hz -0.0257216 -0.0186057
+ 1e+11Hz -0.0257876 -0.0185424
+ 1.001e+11Hz -0.025853 -0.0184784
+ 1.002e+11Hz -0.0259181 -0.0184136
+ 1.003e+11Hz -0.0259826 -0.0183483
+ 1.004e+11Hz -0.0260467 -0.0182822
+ 1.005e+11Hz -0.0261103 -0.0182155
+ 1.006e+11Hz -0.0261734 -0.0181482
+ 1.007e+11Hz -0.0262359 -0.0180802
+ 1.008e+11Hz -0.026298 -0.0180116
+ 1.009e+11Hz -0.0263595 -0.0179424
+ 1.01e+11Hz -0.0264205 -0.0178725
+ 1.011e+11Hz -0.026481 -0.0178021
+ 1.012e+11Hz -0.0265409 -0.017731
+ 1.013e+11Hz -0.0266002 -0.0176593
+ 1.014e+11Hz -0.026659 -0.0175871
+ 1.015e+11Hz -0.0267171 -0.0175143
+ 1.016e+11Hz -0.0267747 -0.0174409
+ 1.017e+11Hz -0.0268317 -0.017367
+ 1.018e+11Hz -0.0268881 -0.0172925
+ 1.019e+11Hz -0.0269438 -0.0172175
+ 1.02e+11Hz -0.026999 -0.017142
+ 1.021e+11Hz -0.0270535 -0.0170659
+ 1.022e+11Hz -0.0271073 -0.0169894
+ 1.023e+11Hz -0.0271606 -0.0169123
+ 1.024e+11Hz -0.0272131 -0.0168347
+ 1.025e+11Hz -0.0272651 -0.0167567
+ 1.026e+11Hz -0.0273163 -0.0166782
+ 1.027e+11Hz -0.0273669 -0.0165993
+ 1.028e+11Hz -0.0274168 -0.0165199
+ 1.029e+11Hz -0.027466 -0.0164401
+ 1.03e+11Hz -0.0275146 -0.0163598
+ 1.031e+11Hz -0.0275624 -0.0162791
+ 1.032e+11Hz -0.0276095 -0.0161981
+ 1.033e+11Hz -0.027656 -0.0161166
+ 1.034e+11Hz -0.0277017 -0.0160347
+ 1.035e+11Hz -0.0277467 -0.0159525
+ 1.036e+11Hz -0.027791 -0.0158699
+ 1.037e+11Hz -0.0278346 -0.015787
+ 1.038e+11Hz -0.0278775 -0.0157037
+ 1.039e+11Hz -0.0279196 -0.0156201
+ 1.04e+11Hz -0.027961 -0.0155362
+ 1.041e+11Hz -0.0280017 -0.015452
+ 1.042e+11Hz -0.0280416 -0.0153675
+ 1.043e+11Hz -0.0280808 -0.0152827
+ 1.044e+11Hz -0.0281193 -0.0151976
+ 1.045e+11Hz -0.028157 -0.0151123
+ 1.046e+11Hz -0.028194 -0.0150267
+ 1.047e+11Hz -0.0282302 -0.0149409
+ 1.048e+11Hz -0.0282657 -0.0148549
+ 1.049e+11Hz -0.0283004 -0.0147686
+ 1.05e+11Hz -0.0283344 -0.0146821
+ 1.051e+11Hz -0.0283676 -0.0145955
+ 1.052e+11Hz -0.0284 -0.0145086
+ 1.053e+11Hz -0.0284317 -0.0144216
+ 1.054e+11Hz -0.0284627 -0.0143344
+ 1.055e+11Hz -0.0284929 -0.0142471
+ 1.056e+11Hz -0.0285223 -0.0141596
+ 1.057e+11Hz -0.028551 -0.014072
+ 1.058e+11Hz -0.028579 -0.0139843
+ 1.059e+11Hz -0.0286062 -0.0138965
+ 1.06e+11Hz -0.0286326 -0.0138086
+ 1.061e+11Hz -0.0286583 -0.0137206
+ 1.062e+11Hz -0.0286832 -0.0136325
+ 1.063e+11Hz -0.0287074 -0.0135443
+ 1.064e+11Hz -0.0287309 -0.0134561
+ 1.065e+11Hz -0.0287536 -0.0133679
+ 1.066e+11Hz -0.0287755 -0.0132796
+ 1.067e+11Hz -0.0287967 -0.0131913
+ 1.068e+11Hz -0.0288172 -0.013103
+ 1.069e+11Hz -0.0288369 -0.0130147
+ 1.07e+11Hz -0.0288559 -0.0129263
+ 1.071e+11Hz -0.0288742 -0.012838
+ 1.072e+11Hz -0.0288918 -0.0127497
+ 1.073e+11Hz -0.0289086 -0.0126615
+ 1.074e+11Hz -0.0289247 -0.0125733
+ 1.075e+11Hz -0.0289401 -0.0124851
+ 1.076e+11Hz -0.0289547 -0.0123971
+ 1.077e+11Hz -0.0289687 -0.012309
+ 1.078e+11Hz -0.028982 -0.0122211
+ 1.079e+11Hz -0.0289945 -0.0121333
+ 1.08e+11Hz -0.0290064 -0.0120455
+ 1.081e+11Hz -0.0290175 -0.0119579
+ 1.082e+11Hz -0.029028 -0.0118703
+ 1.083e+11Hz -0.0290378 -0.0117829
+ 1.084e+11Hz -0.0290469 -0.0116957
+ 1.085e+11Hz -0.0290553 -0.0116085
+ 1.086e+11Hz -0.029063 -0.0115216
+ 1.087e+11Hz -0.0290701 -0.0114347
+ 1.088e+11Hz -0.0290766 -0.0113481
+ 1.089e+11Hz -0.0290823 -0.0112616
+ 1.09e+11Hz -0.0290874 -0.0111753
+ 1.091e+11Hz -0.0290919 -0.0110892
+ 1.092e+11Hz -0.0290958 -0.0110032
+ 1.093e+11Hz -0.029099 -0.0109175
+ 1.094e+11Hz -0.0291015 -0.010832
+ 1.095e+11Hz -0.0291035 -0.0107467
+ 1.096e+11Hz -0.0291048 -0.0106616
+ 1.097e+11Hz -0.0291055 -0.0105768
+ 1.098e+11Hz -0.0291056 -0.0104922
+ 1.099e+11Hz -0.0291052 -0.0104078
+ 1.1e+11Hz -0.0291041 -0.0103237
+ 1.101e+11Hz -0.0291024 -0.0102398
+ 1.102e+11Hz -0.0291002 -0.0101562
+ 1.103e+11Hz -0.0290974 -0.0100728
+ 1.104e+11Hz -0.029094 -0.00998977
+ 1.105e+11Hz -0.02909 -0.00990698
+ 1.106e+11Hz -0.0290855 -0.00982446
+ 1.107e+11Hz -0.0290805 -0.00974224
+ 1.108e+11Hz -0.0290749 -0.0096603
+ 1.109e+11Hz -0.0290688 -0.00957867
+ 1.11e+11Hz -0.0290621 -0.00949733
+ 1.111e+11Hz -0.029055 -0.0094163
+ 1.112e+11Hz -0.0290473 -0.00933559
+ 1.113e+11Hz -0.0290391 -0.00925519
+ 1.114e+11Hz -0.0290304 -0.0091751
+ 1.115e+11Hz -0.0290212 -0.00909535
+ 1.116e+11Hz -0.0290116 -0.00901592
+ 1.117e+11Hz -0.0290014 -0.00893682
+ 1.118e+11Hz -0.0289908 -0.00885805
+ 1.119e+11Hz -0.0289797 -0.00877963
+ 1.12e+11Hz -0.0289682 -0.00870155
+ 1.121e+11Hz -0.0289562 -0.00862381
+ 1.122e+11Hz -0.0289438 -0.00854642
+ 1.123e+11Hz -0.0289309 -0.00846938
+ 1.124e+11Hz -0.0289176 -0.00839269
+ 1.125e+11Hz -0.0289039 -0.00831636
+ 1.126e+11Hz -0.0288898 -0.00824039
+ 1.127e+11Hz -0.0288752 -0.00816478
+ 1.128e+11Hz -0.0288603 -0.00808953
+ 1.129e+11Hz -0.028845 -0.00801465
+ 1.13e+11Hz -0.0288293 -0.00794013
+ 1.131e+11Hz -0.0288132 -0.00786599
+ 1.132e+11Hz -0.0287967 -0.00779221
+ 1.133e+11Hz -0.0287798 -0.00771881
+ 1.134e+11Hz -0.0287626 -0.00764578
+ 1.135e+11Hz -0.0287451 -0.00757312
+ 1.136e+11Hz -0.0287272 -0.00750084
+ 1.137e+11Hz -0.028709 -0.00742894
+ 1.138e+11Hz -0.0286904 -0.00735742
+ 1.139e+11Hz -0.0286715 -0.00728627
+ 1.14e+11Hz -0.0286523 -0.0072155
+ 1.141e+11Hz -0.0286328 -0.00714512
+ 1.142e+11Hz -0.028613 -0.00707511
+ 1.143e+11Hz -0.0285929 -0.00700548
+ 1.144e+11Hz -0.0285725 -0.00693623
+ 1.145e+11Hz -0.0285518 -0.00686737
+ 1.146e+11Hz -0.0285308 -0.00679888
+ 1.147e+11Hz -0.0285096 -0.00673077
+ 1.148e+11Hz -0.0284881 -0.00666305
+ 1.149e+11Hz -0.0284664 -0.0065957
+ 1.15e+11Hz -0.0284444 -0.00652873
+ 1.151e+11Hz -0.0284221 -0.00646214
+ 1.152e+11Hz -0.0283996 -0.00639592
+ 1.153e+11Hz -0.0283769 -0.00633009
+ 1.154e+11Hz -0.028354 -0.00626462
+ 1.155e+11Hz -0.0283308 -0.00619954
+ 1.156e+11Hz -0.0283074 -0.00613482
+ 1.157e+11Hz -0.0282838 -0.00607048
+ 1.158e+11Hz -0.02826 -0.00600651
+ 1.159e+11Hz -0.028236 -0.0059429
+ 1.16e+11Hz -0.0282118 -0.00587967
+ 1.161e+11Hz -0.0281875 -0.0058168
+ 1.162e+11Hz -0.0281629 -0.00575429
+ 1.163e+11Hz -0.0281382 -0.00569215
+ 1.164e+11Hz -0.0281133 -0.00563037
+ 1.165e+11Hz -0.0280882 -0.00556894
+ 1.166e+11Hz -0.028063 -0.00550788
+ 1.167e+11Hz -0.0280376 -0.00544716
+ 1.168e+11Hz -0.0280121 -0.0053868
+ 1.169e+11Hz -0.0279865 -0.00532679
+ 1.17e+11Hz -0.0279607 -0.00526713
+ 1.171e+11Hz -0.0279347 -0.00520781
+ 1.172e+11Hz -0.0279086 -0.00514884
+ 1.173e+11Hz -0.0278825 -0.00509021
+ 1.174e+11Hz -0.0278561 -0.00503191
+ 1.175e+11Hz -0.0278297 -0.00497395
+ 1.176e+11Hz -0.0278032 -0.00491632
+ 1.177e+11Hz -0.0277765 -0.00485902
+ 1.178e+11Hz -0.0277498 -0.00480205
+ 1.179e+11Hz -0.0277229 -0.00474541
+ 1.18e+11Hz -0.027696 -0.00468908
+ 1.181e+11Hz -0.0276689 -0.00463308
+ 1.182e+11Hz -0.0276418 -0.00457739
+ 1.183e+11Hz -0.0276146 -0.00452201
+ 1.184e+11Hz -0.0275873 -0.00446694
+ 1.185e+11Hz -0.0275599 -0.00441218
+ 1.186e+11Hz -0.0275325 -0.00435772
+ 1.187e+11Hz -0.0275049 -0.00430357
+ 1.188e+11Hz -0.0274774 -0.00424971
+ 1.189e+11Hz -0.0274497 -0.00419614
+ 1.19e+11Hz -0.027422 -0.00414287
+ 1.191e+11Hz -0.0273942 -0.00408989
+ 1.192e+11Hz -0.0273664 -0.00403719
+ 1.193e+11Hz -0.0273385 -0.00398477
+ 1.194e+11Hz -0.0273106 -0.00393263
+ 1.195e+11Hz -0.0272826 -0.00388077
+ 1.196e+11Hz -0.0272546 -0.00382918
+ 1.197e+11Hz -0.0272265 -0.00377786
+ 1.198e+11Hz -0.0271984 -0.0037268
+ 1.199e+11Hz -0.0271703 -0.00367601
+ 1.2e+11Hz -0.0271421 -0.00362547
+ 1.201e+11Hz -0.0271139 -0.0035752
+ 1.202e+11Hz -0.0270857 -0.00352517
+ 1.203e+11Hz -0.0270574 -0.0034754
+ 1.204e+11Hz -0.0270291 -0.00342587
+ 1.205e+11Hz -0.0270008 -0.00337659
+ 1.206e+11Hz -0.0269724 -0.00332755
+ 1.207e+11Hz -0.0269441 -0.00327874
+ 1.208e+11Hz -0.0269157 -0.00323017
+ 1.209e+11Hz -0.0268873 -0.00318183
+ 1.21e+11Hz -0.0268588 -0.00313372
+ 1.211e+11Hz -0.0268304 -0.00308584
+ 1.212e+11Hz -0.0268019 -0.00303817
+ 1.213e+11Hz -0.0267734 -0.00299073
+ 1.214e+11Hz -0.0267449 -0.0029435
+ 1.215e+11Hz -0.0267164 -0.00289649
+ 1.216e+11Hz -0.0266879 -0.00284969
+ 1.217e+11Hz -0.0266594 -0.00280309
+ 1.218e+11Hz -0.0266308 -0.0027567
+ 1.219e+11Hz -0.0266023 -0.00271051
+ 1.22e+11Hz -0.0265737 -0.00266452
+ 1.221e+11Hz -0.0265452 -0.00261873
+ 1.222e+11Hz -0.0265166 -0.00257313
+ 1.223e+11Hz -0.026488 -0.00252772
+ 1.224e+11Hz -0.0264594 -0.00248251
+ 1.225e+11Hz -0.0264309 -0.00243747
+ 1.226e+11Hz -0.0264023 -0.00239263
+ 1.227e+11Hz -0.0263737 -0.00234796
+ 1.228e+11Hz -0.0263451 -0.00230347
+ 1.229e+11Hz -0.0263165 -0.00225916
+ 1.23e+11Hz -0.0262878 -0.00221502
+ 1.231e+11Hz -0.0262592 -0.00217105
+ 1.232e+11Hz -0.0262306 -0.00212725
+ 1.233e+11Hz -0.026202 -0.00208362
+ 1.234e+11Hz -0.0261734 -0.00204016
+ 1.235e+11Hz -0.0261448 -0.00199686
+ 1.236e+11Hz -0.0261162 -0.00195371
+ 1.237e+11Hz -0.0260875 -0.00191073
+ 1.238e+11Hz -0.0260589 -0.0018679
+ 1.239e+11Hz -0.0260303 -0.00182523
+ 1.24e+11Hz -0.0260017 -0.00178271
+ 1.241e+11Hz -0.025973 -0.00174034
+ 1.242e+11Hz -0.0259444 -0.00169812
+ 1.243e+11Hz -0.0259158 -0.00165605
+ 1.244e+11Hz -0.0258872 -0.00161412
+ 1.245e+11Hz -0.0258585 -0.00157233
+ 1.246e+11Hz -0.0258299 -0.00153069
+ 1.247e+11Hz -0.0258013 -0.00148918
+ 1.248e+11Hz -0.0257726 -0.00144782
+ 1.249e+11Hz -0.025744 -0.00140659
+ 1.25e+11Hz -0.0257154 -0.00136549
+ 1.251e+11Hz -0.0256868 -0.00132453
+ 1.252e+11Hz -0.0256581 -0.0012837
+ 1.253e+11Hz -0.0256295 -0.001243
+ 1.254e+11Hz -0.0256009 -0.00120243
+ 1.255e+11Hz -0.0255722 -0.00116198
+ 1.256e+11Hz -0.0255436 -0.00112166
+ 1.257e+11Hz -0.025515 -0.00108147
+ 1.258e+11Hz -0.0254863 -0.00104139
+ 1.259e+11Hz -0.0254577 -0.00100144
+ 1.26e+11Hz -0.0254291 -0.000961613
+ 1.261e+11Hz -0.0254005 -0.0009219
+ 1.262e+11Hz -0.0253718 -0.000882305
+ 1.263e+11Hz -0.0253432 -0.000842826
+ 1.264e+11Hz -0.0253146 -0.000803461
+ 1.265e+11Hz -0.025286 -0.000764209
+ 1.266e+11Hz -0.0252573 -0.000725069
+ 1.267e+11Hz -0.0252287 -0.00068604
+ 1.268e+11Hz -0.0252001 -0.000647119
+ 1.269e+11Hz -0.0251715 -0.000608307
+ 1.27e+11Hz -0.0251429 -0.0005696
+ 1.271e+11Hz -0.0251143 -0.000530999
+ 1.272e+11Hz -0.0250857 -0.000492502
+ 1.273e+11Hz -0.0250571 -0.000454107
+ 1.274e+11Hz -0.0250285 -0.000415812
+ 1.275e+11Hz -0.0249999 -0.000377618
+ 1.276e+11Hz -0.0249713 -0.000339522
+ 1.277e+11Hz -0.0249428 -0.000301522
+ 1.278e+11Hz -0.0249142 -0.000263618
+ 1.279e+11Hz -0.0248856 -0.000225807
+ 1.28e+11Hz -0.0248571 -0.000188089
+ 1.281e+11Hz -0.0248285 -0.000150462
+ 1.282e+11Hz -0.0248 -0.000112925
+ 1.283e+11Hz -0.0247715 -7.54747e-05
+ 1.284e+11Hz -0.0247429 -3.81111e-05
+ 1.285e+11Hz -0.0247144 -8.32039e-07
+ 1.286e+11Hz -0.0246859 3.6364e-05
+ 1.287e+11Hz -0.0246575 7.34787e-05
+ 1.288e+11Hz -0.024629 0.000110514
+ 1.289e+11Hz -0.0246005 0.000147471
+ 1.29e+11Hz -0.0245721 0.000184353
+ 1.291e+11Hz -0.0245436 0.00022116
+ 1.292e+11Hz -0.0245152 0.000257894
+ 1.293e+11Hz -0.0244868 0.000294559
+ 1.294e+11Hz -0.0244584 0.000331155
+ 1.295e+11Hz -0.02443 0.000367684
+ 1.296e+11Hz -0.0244017 0.000404149
+ 1.297e+11Hz -0.0243733 0.000440552
+ 1.298e+11Hz -0.024345 0.000476895
+ 1.299e+11Hz -0.0243167 0.000513179
+ 1.3e+11Hz -0.0242884 0.000549408
+ 1.301e+11Hz -0.0242601 0.000585584
+ 1.302e+11Hz -0.0242319 0.000621709
+ 1.303e+11Hz -0.0242036 0.000657784
+ 1.304e+11Hz -0.0241754 0.000693814
+ 1.305e+11Hz -0.0241472 0.0007298
+ 1.306e+11Hz -0.0241191 0.000765745
+ 1.307e+11Hz -0.0240909 0.000801651
+ 1.308e+11Hz -0.0240628 0.000837522
+ 1.309e+11Hz -0.0240347 0.000873359
+ 1.31e+11Hz -0.0240066 0.000909166
+ 1.311e+11Hz -0.0239785 0.000944945
+ 1.312e+11Hz -0.0239504 0.0009807
+ 1.313e+11Hz -0.0239224 0.00101643
+ 1.314e+11Hz -0.0238944 0.00105215
+ 1.315e+11Hz -0.0238664 0.00108785
+ 1.316e+11Hz -0.0238385 0.00112353
+ 1.317e+11Hz -0.0238105 0.00115921
+ 1.318e+11Hz -0.0237826 0.00119488
+ 1.319e+11Hz -0.0237547 0.00123054
+ 1.32e+11Hz -0.0237268 0.00126621
+ 1.321e+11Hz -0.023699 0.00130188
+ 1.322e+11Hz -0.0236711 0.00133755
+ 1.323e+11Hz -0.0236433 0.00137324
+ 1.324e+11Hz -0.0236155 0.00140894
+ 1.325e+11Hz -0.0235877 0.00144466
+ 1.326e+11Hz -0.0235599 0.00148039
+ 1.327e+11Hz -0.0235321 0.00151616
+ 1.328e+11Hz -0.0235044 0.00155194
+ 1.329e+11Hz -0.0234766 0.00158776
+ 1.33e+11Hz -0.0234489 0.00162362
+ 1.331e+11Hz -0.0234212 0.00165951
+ 1.332e+11Hz -0.0233935 0.00169545
+ 1.333e+11Hz -0.0233658 0.00173143
+ 1.334e+11Hz -0.0233381 0.00176746
+ 1.335e+11Hz -0.0233103 0.00180354
+ 1.336e+11Hz -0.0232826 0.00183968
+ 1.337e+11Hz -0.0232549 0.00187588
+ 1.338e+11Hz -0.0232272 0.00191214
+ 1.339e+11Hz -0.0231995 0.00194847
+ 1.34e+11Hz -0.0231718 0.00198488
+ 1.341e+11Hz -0.0231441 0.00202135
+ 1.342e+11Hz -0.0231163 0.00205791
+ 1.343e+11Hz -0.0230885 0.00209455
+ 1.344e+11Hz -0.0230608 0.00213128
+ 1.345e+11Hz -0.0230329 0.0021681
+ 1.346e+11Hz -0.0230051 0.002205
+ 1.347e+11Hz -0.0229772 0.00224201
+ 1.348e+11Hz -0.0229493 0.00227912
+ 1.349e+11Hz -0.0229214 0.00231633
+ 1.35e+11Hz -0.0228934 0.00235365
+ 1.351e+11Hz -0.0228654 0.00239108
+ 1.352e+11Hz -0.0228374 0.00242863
+ 1.353e+11Hz -0.0228092 0.00246629
+ 1.354e+11Hz -0.0227811 0.00250408
+ 1.355e+11Hz -0.0227528 0.00254198
+ 1.356e+11Hz -0.0227245 0.00258002
+ 1.357e+11Hz -0.0226962 0.00261819
+ 1.358e+11Hz -0.0226677 0.00265649
+ 1.359e+11Hz -0.0226392 0.00269492
+ 1.36e+11Hz -0.0226106 0.0027335
+ 1.361e+11Hz -0.0225819 0.00277222
+ 1.362e+11Hz -0.0225532 0.00281108
+ 1.363e+11Hz -0.0225243 0.00285009
+ 1.364e+11Hz -0.0224953 0.00288925
+ 1.365e+11Hz -0.0224662 0.00292856
+ 1.366e+11Hz -0.022437 0.00296803
+ 1.367e+11Hz -0.0224077 0.00300765
+ 1.368e+11Hz -0.0223782 0.00304743
+ 1.369e+11Hz -0.0223486 0.00308737
+ 1.37e+11Hz -0.0223189 0.00312747
+ 1.371e+11Hz -0.022289 0.00316774
+ 1.372e+11Hz -0.022259 0.00320817
+ 1.373e+11Hz -0.0222288 0.00324877
+ 1.374e+11Hz -0.0221984 0.00328954
+ 1.375e+11Hz -0.0221679 0.00333047
+ 1.376e+11Hz -0.0221372 0.00337158
+ 1.377e+11Hz -0.0221063 0.00341286
+ 1.378e+11Hz -0.0220752 0.0034543
+ 1.379e+11Hz -0.022044 0.00349592
+ 1.38e+11Hz -0.0220125 0.00353771
+ 1.381e+11Hz -0.0219808 0.00357968
+ 1.382e+11Hz -0.0219489 0.00362181
+ 1.383e+11Hz -0.0219167 0.00366412
+ 1.384e+11Hz -0.0218843 0.0037066
+ 1.385e+11Hz -0.0218517 0.00374925
+ 1.386e+11Hz -0.0218189 0.00379207
+ 1.387e+11Hz -0.0217857 0.00383506
+ 1.388e+11Hz -0.0217524 0.00387822
+ 1.389e+11Hz -0.0217187 0.00392154
+ 1.39e+11Hz -0.0216848 0.00396503
+ 1.391e+11Hz -0.0216505 0.00400868
+ 1.392e+11Hz -0.021616 0.0040525
+ 1.393e+11Hz -0.0215812 0.00409647
+ 1.394e+11Hz -0.0215461 0.00414061
+ 1.395e+11Hz -0.0215106 0.00418489
+ 1.396e+11Hz -0.0214749 0.00422933
+ 1.397e+11Hz -0.0214388 0.00427392
+ 1.398e+11Hz -0.0214023 0.00431865
+ 1.399e+11Hz -0.0213655 0.00436353
+ 1.4e+11Hz -0.0213284 0.00440855
+ 1.401e+11Hz -0.0212909 0.0044537
+ 1.402e+11Hz -0.021253 0.00449898
+ 1.403e+11Hz -0.0212147 0.00454439
+ 1.404e+11Hz -0.0211761 0.00458993
+ 1.405e+11Hz -0.0211371 0.00463558
+ 1.406e+11Hz -0.0210976 0.00468135
+ 1.407e+11Hz -0.0210578 0.00472722
+ 1.408e+11Hz -0.0210176 0.0047732
+ 1.409e+11Hz -0.0209769 0.00481928
+ 1.41e+11Hz -0.0209358 0.00486545
+ 1.411e+11Hz -0.0208942 0.0049117
+ 1.412e+11Hz -0.0208523 0.00495804
+ 1.413e+11Hz -0.0208098 0.00500445
+ 1.414e+11Hz -0.020767 0.00505093
+ 1.415e+11Hz -0.0207236 0.00509747
+ 1.416e+11Hz -0.0206798 0.00514406
+ 1.417e+11Hz -0.0206355 0.00519071
+ 1.418e+11Hz -0.0205907 0.00523739
+ 1.419e+11Hz -0.0205455 0.00528411
+ 1.42e+11Hz -0.0204997 0.00533085
+ 1.421e+11Hz -0.0204535 0.00537761
+ 1.422e+11Hz -0.0204068 0.00542438
+ 1.423e+11Hz -0.0203595 0.00547115
+ 1.424e+11Hz -0.0203117 0.00551791
+ 1.425e+11Hz -0.0202634 0.00556466
+ 1.426e+11Hz -0.0202146 0.00561139
+ 1.427e+11Hz -0.0201653 0.00565808
+ 1.428e+11Hz -0.0201154 0.00570473
+ 1.429e+11Hz -0.0200649 0.00575133
+ 1.43e+11Hz -0.020014 0.00579787
+ 1.431e+11Hz -0.0199625 0.00584435
+ 1.432e+11Hz -0.0199104 0.00589074
+ 1.433e+11Hz -0.0198578 0.00593704
+ 1.434e+11Hz -0.0198046 0.00598325
+ 1.435e+11Hz -0.0197509 0.00602935
+ 1.436e+11Hz -0.0196966 0.00607533
+ 1.437e+11Hz -0.0196417 0.00612118
+ 1.438e+11Hz -0.0195863 0.00616689
+ 1.439e+11Hz -0.0195302 0.00621246
+ 1.44e+11Hz -0.0194737 0.00625786
+ 1.441e+11Hz -0.0194165 0.0063031
+ 1.442e+11Hz -0.0193588 0.00634815
+ 1.443e+11Hz -0.0193005 0.00639301
+ 1.444e+11Hz -0.0192416 0.00643768
+ 1.445e+11Hz -0.0191821 0.00648212
+ 1.446e+11Hz -0.019122 0.00652635
+ 1.447e+11Hz -0.0190614 0.00657033
+ 1.448e+11Hz -0.0190002 0.00661408
+ 1.449e+11Hz -0.0189384 0.00665756
+ 1.45e+11Hz -0.018876 0.00670078
+ 1.451e+11Hz -0.018813 0.00674371
+ 1.452e+11Hz -0.0187495 0.00678636
+ 1.453e+11Hz -0.0186853 0.00682871
+ 1.454e+11Hz -0.0186206 0.00687074
+ 1.455e+11Hz -0.0185554 0.00691245
+ 1.456e+11Hz -0.0184895 0.00695382
+ 1.457e+11Hz -0.0184231 0.00699485
+ 1.458e+11Hz -0.0183561 0.00703551
+ 1.459e+11Hz -0.0182885 0.00707581
+ 1.46e+11Hz -0.0182204 0.00711573
+ 1.461e+11Hz -0.0181517 0.00715526
+ 1.462e+11Hz -0.0180825 0.00719439
+ 1.463e+11Hz -0.0180127 0.00723311
+ 1.464e+11Hz -0.0179424 0.0072714
+ 1.465e+11Hz -0.0178715 0.00730925
+ 1.466e+11Hz -0.0178 0.00734667
+ 1.467e+11Hz -0.0177281 0.00738362
+ 1.468e+11Hz -0.0176556 0.00742011
+ 1.469e+11Hz -0.0175826 0.00745612
+ 1.47e+11Hz -0.017509 0.00749165
+ 1.471e+11Hz -0.017435 0.00752668
+ 1.472e+11Hz -0.0173604 0.0075612
+ 1.473e+11Hz -0.0172854 0.0075952
+ 1.474e+11Hz -0.0172098 0.00762867
+ 1.475e+11Hz -0.0171337 0.00766161
+ 1.476e+11Hz -0.0170572 0.007694
+ 1.477e+11Hz -0.0169802 0.00772583
+ 1.478e+11Hz -0.0169027 0.0077571
+ 1.479e+11Hz -0.0168248 0.00778779
+ 1.48e+11Hz -0.0167464 0.0078179
+ 1.481e+11Hz -0.0166676 0.00784742
+ 1.482e+11Hz -0.0165883 0.00787633
+ 1.483e+11Hz -0.0165087 0.00790463
+ 1.484e+11Hz -0.0164285 0.00793232
+ 1.485e+11Hz -0.016348 0.00795938
+ 1.486e+11Hz -0.0162671 0.0079858
+ 1.487e+11Hz -0.0161858 0.00801158
+ 1.488e+11Hz -0.0161041 0.00803671
+ 1.489e+11Hz -0.016022 0.00806119
+ 1.49e+11Hz -0.0159396 0.008085
+ 1.491e+11Hz -0.0158568 0.00810814
+ 1.492e+11Hz -0.0157737 0.0081306
+ 1.493e+11Hz -0.0156902 0.00815238
+ 1.494e+11Hz -0.0156064 0.00817346
+ 1.495e+11Hz -0.0155223 0.00819385
+ 1.496e+11Hz -0.0154379 0.00821354
+ 1.497e+11Hz -0.0153532 0.00823252
+ 1.498e+11Hz -0.0152682 0.00825078
+ 1.499e+11Hz -0.015183 0.00826833
+ 1.5e+11Hz -0.0150975 0.00828515
+ 1.501e+11Hz -0.0150117 0.00830125
+ 1.502e+11Hz -0.0149257 0.00831661
+ 1.503e+11Hz -0.0148395 0.00833124
+ 1.504e+11Hz -0.0147531 0.00834513
+ 1.505e+11Hz -0.0146664 0.00835827
+ 1.506e+11Hz -0.0145796 0.00837067
+ 1.507e+11Hz -0.0144926 0.00838231
+ 1.508e+11Hz -0.0144054 0.0083932
+ 1.509e+11Hz -0.014318 0.00840334
+ 1.51e+11Hz -0.0142305 0.00841272
+ 1.511e+11Hz -0.0141429 0.00842134
+ 1.512e+11Hz -0.0140552 0.00842919
+ 1.513e+11Hz -0.0139673 0.00843628
+ 1.514e+11Hz -0.0138793 0.00844261
+ 1.515e+11Hz -0.0137913 0.00844817
+ 1.516e+11Hz -0.0137031 0.00845296
+ 1.517e+11Hz -0.0136149 0.00845699
+ 1.518e+11Hz -0.0135267 0.00846025
+ 1.519e+11Hz -0.0134384 0.00846274
+ 1.52e+11Hz -0.0133501 0.00846446
+ 1.521e+11Hz -0.0132617 0.00846542
+ 1.522e+11Hz -0.0131734 0.0084656
+ 1.523e+11Hz -0.013085 0.00846503
+ 1.524e+11Hz -0.0129967 0.00846368
+ 1.525e+11Hz -0.0129084 0.00846158
+ 1.526e+11Hz -0.0128201 0.00845871
+ 1.527e+11Hz -0.0127319 0.00845508
+ 1.528e+11Hz -0.0126438 0.00845069
+ 1.529e+11Hz -0.0125557 0.00844555
+ 1.53e+11Hz -0.0124677 0.00843966
+ 1.531e+11Hz -0.0123797 0.00843301
+ 1.532e+11Hz -0.0122919 0.00842562
+ 1.533e+11Hz -0.0122042 0.00841748
+ 1.534e+11Hz -0.0121167 0.0084086
+ 1.535e+11Hz -0.0120292 0.00839898
+ 1.536e+11Hz -0.0119419 0.00838863
+ 1.537e+11Hz -0.0118548 0.00837755
+ 1.538e+11Hz -0.0117678 0.00836575
+ 1.539e+11Hz -0.011681 0.00835322
+ 1.54e+11Hz -0.0115944 0.00833998
+ 1.541e+11Hz -0.011508 0.00832602
+ 1.542e+11Hz -0.0114217 0.00831136
+ 1.543e+11Hz -0.0113357 0.00829599
+ 1.544e+11Hz -0.01125 0.00827993
+ 1.545e+11Hz -0.0111644 0.00826318
+ 1.546e+11Hz -0.0110791 0.00824574
+ 1.547e+11Hz -0.010994 0.00822762
+ 1.548e+11Hz -0.0109092 0.00820882
+ 1.549e+11Hz -0.0108247 0.00818936
+ 1.55e+11Hz -0.0107404 0.00816924
+ 1.551e+11Hz -0.0106564 0.00814845
+ 1.552e+11Hz -0.0105728 0.00812702
+ 1.553e+11Hz -0.0104894 0.00810495
+ 1.554e+11Hz -0.0104063 0.00808223
+ 1.555e+11Hz -0.0103235 0.00805889
+ 1.556e+11Hz -0.010241 0.00803493
+ 1.557e+11Hz -0.0101589 0.00801035
+ 1.558e+11Hz -0.0100771 0.00798515
+ 1.559e+11Hz -0.00999564 0.00795936
+ 1.56e+11Hz -0.00991453 0.00793297
+ 1.561e+11Hz -0.00983377 0.007906
+ 1.562e+11Hz -0.00975337 0.00787844
+ 1.563e+11Hz -0.00967333 0.00785031
+ 1.564e+11Hz -0.00959367 0.00782161
+ 1.565e+11Hz -0.00951437 0.00779236
+ 1.566e+11Hz -0.00943546 0.00776255
+ 1.567e+11Hz -0.00935694 0.00773221
+ 1.568e+11Hz -0.00927881 0.00770132
+ 1.569e+11Hz -0.00920107 0.00766991
+ 1.57e+11Hz -0.00912374 0.00763798
+ 1.571e+11Hz -0.0090468 0.00760554
+ 1.572e+11Hz -0.00897028 0.00757259
+ 1.573e+11Hz -0.00889417 0.00753915
+ 1.574e+11Hz -0.00881848 0.00750522
+ 1.575e+11Hz -0.00874321 0.0074708
+ 1.576e+11Hz -0.00866836 0.00743592
+ 1.577e+11Hz -0.00859394 0.00740057
+ 1.578e+11Hz -0.00851995 0.00736476
+ 1.579e+11Hz -0.00844639 0.0073285
+ 1.58e+11Hz -0.00837327 0.0072918
+ 1.581e+11Hz -0.00830058 0.00725466
+ 1.582e+11Hz -0.00822834 0.0072171
+ 1.583e+11Hz -0.00815654 0.00717912
+ 1.584e+11Hz -0.00808519 0.00714073
+ 1.585e+11Hz -0.00801429 0.00710194
+ 1.586e+11Hz -0.00794383 0.00706275
+ 1.587e+11Hz -0.00787383 0.00702317
+ 1.588e+11Hz -0.00780427 0.00698321
+ 1.589e+11Hz -0.00773518 0.00694288
+ 1.59e+11Hz -0.00766653 0.00690218
+ 1.591e+11Hz -0.00759834 0.00686112
+ 1.592e+11Hz -0.00753061 0.00681972
+ 1.593e+11Hz -0.00746334 0.00677797
+ 1.594e+11Hz -0.00739653 0.00673588
+ 1.595e+11Hz -0.00733017 0.00669347
+ 1.596e+11Hz -0.00726427 0.00665073
+ 1.597e+11Hz -0.00719884 0.00660767
+ 1.598e+11Hz -0.00713386 0.00656431
+ 1.599e+11Hz -0.00706934 0.00652065
+ 1.6e+11Hz -0.00700528 0.00647669
+ 1.601e+11Hz -0.00694169 0.00643245
+ 1.602e+11Hz -0.00687855 0.00638792
+ 1.603e+11Hz -0.00681586 0.00634312
+ 1.604e+11Hz -0.00675364 0.00629805
+ 1.605e+11Hz -0.00669187 0.00625272
+ 1.606e+11Hz -0.00663056 0.00620713
+ 1.607e+11Hz -0.00656971 0.0061613
+ 1.608e+11Hz -0.00650931 0.00611522
+ 1.609e+11Hz -0.00644937 0.0060689
+ 1.61e+11Hz -0.00638988 0.00602235
+ 1.611e+11Hz -0.00633084 0.00597558
+ 1.612e+11Hz -0.00627225 0.00592859
+ 1.613e+11Hz -0.0062141 0.00588138
+ 1.614e+11Hz -0.00615641 0.00583397
+ 1.615e+11Hz -0.00609916 0.00578635
+ 1.616e+11Hz -0.00604236 0.00573854
+ 1.617e+11Hz -0.005986 0.00569053
+ 1.618e+11Hz -0.00593009 0.00564234
+ 1.619e+11Hz -0.00587461 0.00559396
+ 1.62e+11Hz -0.00581957 0.00554541
+ 1.621e+11Hz -0.00576497 0.00549668
+ 1.622e+11Hz -0.0057108 0.00544779
+ 1.623e+11Hz -0.00565707 0.00539874
+ 1.624e+11Hz -0.00560376 0.00534953
+ 1.625e+11Hz -0.00555089 0.00530017
+ 1.626e+11Hz -0.00549844 0.00525066
+ 1.627e+11Hz -0.00544642 0.005201
+ 1.628e+11Hz -0.00539482 0.00515121
+ 1.629e+11Hz -0.00534364 0.00510128
+ 1.63e+11Hz -0.00529288 0.00505122
+ 1.631e+11Hz -0.00524253 0.00500103
+ 1.632e+11Hz -0.00519261 0.00495072
+ 1.633e+11Hz -0.00514309 0.00490029
+ 1.634e+11Hz -0.00509398 0.00484974
+ 1.635e+11Hz -0.00504529 0.00479909
+ 1.636e+11Hz -0.004997 0.00474832
+ 1.637e+11Hz -0.00494911 0.00469746
+ 1.638e+11Hz -0.00490162 0.00464649
+ 1.639e+11Hz -0.00485454 0.00459542
+ 1.64e+11Hz -0.00480785 0.00454426
+ 1.641e+11Hz -0.00476156 0.00449301
+ 1.642e+11Hz -0.00471566 0.00444167
+ 1.643e+11Hz -0.00467015 0.00439025
+ 1.644e+11Hz -0.00462503 0.00433875
+ 1.645e+11Hz -0.0045803 0.00428717
+ 1.646e+11Hz -0.00453595 0.00423551
+ 1.647e+11Hz -0.00449198 0.00418379
+ 1.648e+11Hz -0.0044484 0.00413199
+ 1.649e+11Hz -0.00440519 0.00408013
+ 1.65e+11Hz -0.00436236 0.00402821
+ 1.651e+11Hz -0.0043199 0.00397622
+ 1.652e+11Hz -0.00427781 0.00392418
+ 1.653e+11Hz -0.00423609 0.00387208
+ 1.654e+11Hz -0.00419474 0.00381993
+ 1.655e+11Hz -0.00415376 0.00376773
+ 1.656e+11Hz -0.00411313 0.00371548
+ 1.657e+11Hz -0.00407287 0.00366319
+ 1.658e+11Hz -0.00403297 0.00361086
+ 1.659e+11Hz -0.00399343 0.00355848
+ 1.66e+11Hz -0.00395424 0.00350607
+ 1.661e+11Hz -0.0039154 0.00345362
+ 1.662e+11Hz -0.00387692 0.00340114
+ 1.663e+11Hz -0.00383878 0.00334863
+ 1.664e+11Hz -0.00380099 0.00329608
+ 1.665e+11Hz -0.00376355 0.00324352
+ 1.666e+11Hz -0.00372645 0.00319092
+ 1.667e+11Hz -0.00368969 0.00313831
+ 1.668e+11Hz -0.00365327 0.00308567
+ 1.669e+11Hz -0.00361719 0.00303302
+ 1.67e+11Hz -0.00358144 0.00298035
+ 1.671e+11Hz -0.00354603 0.00292767
+ 1.672e+11Hz -0.00351095 0.00287497
+ 1.673e+11Hz -0.0034762 0.00282227
+ 1.674e+11Hz -0.00344178 0.00276955
+ 1.675e+11Hz -0.00340768 0.00271683
+ 1.676e+11Hz -0.00337391 0.00266411
+ 1.677e+11Hz -0.00334046 0.00261138
+ 1.678e+11Hz -0.00330733 0.00255866
+ 1.679e+11Hz -0.00327452 0.00250593
+ 1.68e+11Hz -0.00324203 0.00245321
+ 1.681e+11Hz -0.00320985 0.00240049
+ 1.682e+11Hz -0.00317799 0.00234778
+ 1.683e+11Hz -0.00314644 0.00229508
+ 1.684e+11Hz -0.0031152 0.00224239
+ 1.685e+11Hz -0.00308427 0.00218971
+ 1.686e+11Hz -0.00305364 0.00213705
+ 1.687e+11Hz -0.00302332 0.0020844
+ 1.688e+11Hz -0.0029933 0.00203177
+ 1.689e+11Hz -0.00296358 0.00197916
+ 1.69e+11Hz -0.00293416 0.00192657
+ 1.691e+11Hz -0.00290504 0.001874
+ 1.692e+11Hz -0.00287621 0.00182146
+ 1.693e+11Hz -0.00284768 0.00176894
+ 1.694e+11Hz -0.00281944 0.00171645
+ 1.695e+11Hz -0.00279149 0.00166399
+ 1.696e+11Hz -0.00276383 0.00161156
+ 1.697e+11Hz -0.00273645 0.00155917
+ 1.698e+11Hz -0.00270936 0.00150681
+ 1.699e+11Hz -0.00268255 0.00145448
+ 1.7e+11Hz -0.00265602 0.00140219
+ 1.701e+11Hz -0.00262977 0.00134994
+ 1.702e+11Hz -0.0026038 0.00129774
+ 1.703e+11Hz -0.00257811 0.00124557
+ 1.704e+11Hz -0.00255268 0.00119345
+ 1.705e+11Hz -0.00252753 0.00114137
+ 1.706e+11Hz -0.00250265 0.00108934
+ 1.707e+11Hz -0.00247804 0.00103735
+ 1.708e+11Hz -0.00245369 0.00098542
+ 1.709e+11Hz -0.0024296 0.000933538
+ 1.71e+11Hz -0.00240578 0.000881707
+ 1.711e+11Hz -0.00238222 0.00082993
+ 1.712e+11Hz -0.00235891 0.000778209
+ 1.713e+11Hz -0.00233586 0.000726543
+ 1.714e+11Hz -0.00231306 0.000674936
+ 1.715e+11Hz -0.00229052 0.000623387
+ 1.716e+11Hz -0.00226823 0.000571899
+ 1.717e+11Hz -0.00224618 0.000520472
+ 1.718e+11Hz -0.00222438 0.000469108
+ 1.719e+11Hz -0.00220282 0.000417807
+ 1.72e+11Hz -0.00218151 0.000366572
+ 1.721e+11Hz -0.00216043 0.000315403
+ 1.722e+11Hz -0.00213959 0.000264302
+ 1.723e+11Hz -0.00211899 0.000213268
+ 1.724e+11Hz -0.00209862 0.000162304
+ 1.725e+11Hz -0.00207848 0.000111411
+ 1.726e+11Hz -0.00205857 6.0589e-05
+ 1.727e+11Hz -0.00203889 9.83952e-06
+ 1.728e+11Hz -0.00201943 -4.08367e-05
+ 1.729e+11Hz -0.0020002 -9.14386e-05
+ 1.73e+11Hz -0.00198118 -0.000141965
+ 1.731e+11Hz -0.00196239 -0.000192416
+ 1.732e+11Hz -0.00194381 -0.00024279
+ 1.733e+11Hz -0.00192544 -0.000293087
+ 1.734e+11Hz -0.00190729 -0.000343305
+ 1.735e+11Hz -0.00188934 -0.000393445
+ 1.736e+11Hz -0.00187161 -0.000443505
+ 1.737e+11Hz -0.00185408 -0.000493484
+ 1.738e+11Hz -0.00183675 -0.000543383
+ 1.739e+11Hz -0.00181963 -0.0005932
+ 1.74e+11Hz -0.0018027 -0.000642935
+ 1.741e+11Hz -0.00178597 -0.000692588
+ 1.742e+11Hz -0.00176944 -0.000742158
+ 1.743e+11Hz -0.0017531 -0.000791644
+ 1.744e+11Hz -0.00173695 -0.000841047
+ 1.745e+11Hz -0.00172099 -0.000890365
+ 1.746e+11Hz -0.00170521 -0.000939599
+ 1.747e+11Hz -0.00168962 -0.000988748
+ 1.748e+11Hz -0.00167421 -0.00103781
+ 1.749e+11Hz -0.00165899 -0.00108679
+ 1.75e+11Hz -0.00164394 -0.00113568
+ 1.751e+11Hz -0.00162907 -0.00118449
+ 1.752e+11Hz -0.00161437 -0.00123321
+ 1.753e+11Hz -0.00159985 -0.00128185
+ 1.754e+11Hz -0.00158549 -0.0013304
+ 1.755e+11Hz -0.00157131 -0.00137886
+ 1.756e+11Hz -0.00155729 -0.00142724
+ 1.757e+11Hz -0.00154344 -0.00147553
+ 1.758e+11Hz -0.00152975 -0.00152374
+ 1.759e+11Hz -0.00151622 -0.00157186
+ 1.76e+11Hz -0.00150285 -0.00161989
+ 1.761e+11Hz -0.00148964 -0.00166784
+ 1.762e+11Hz -0.00147658 -0.0017157
+ 1.763e+11Hz -0.00146368 -0.00176348
+ 1.764e+11Hz -0.00145093 -0.00181117
+ 1.765e+11Hz -0.00143833 -0.00185877
+ 1.766e+11Hz -0.00142588 -0.00190629
+ 1.767e+11Hz -0.00141358 -0.00195373
+ 1.768e+11Hz -0.00140142 -0.00200108
+ 1.769e+11Hz -0.00138941 -0.00204834
+ 1.77e+11Hz -0.00137754 -0.00209552
+ 1.771e+11Hz -0.00136581 -0.00214262
+ 1.772e+11Hz -0.00135422 -0.00218964
+ 1.773e+11Hz -0.00134277 -0.00223657
+ 1.774e+11Hz -0.00133146 -0.00228341
+ 1.775e+11Hz -0.00132028 -0.00233018
+ 1.776e+11Hz -0.00130923 -0.00237686
+ 1.777e+11Hz -0.00129832 -0.00242346
+ 1.778e+11Hz -0.00128754 -0.00246998
+ 1.779e+11Hz -0.00127689 -0.00251641
+ 1.78e+11Hz -0.00126637 -0.00256277
+ 1.781e+11Hz -0.00125597 -0.00260904
+ 1.782e+11Hz -0.0012457 -0.00265523
+ 1.783e+11Hz -0.00123556 -0.00270134
+ 1.784e+11Hz -0.00122554 -0.00274738
+ 1.785e+11Hz -0.00121564 -0.00279333
+ 1.786e+11Hz -0.00120587 -0.0028392
+ 1.787e+11Hz -0.00119621 -0.00288499
+ 1.788e+11Hz -0.00118668 -0.0029307
+ 1.789e+11Hz -0.00117726 -0.00297634
+ 1.79e+11Hz -0.00116796 -0.00302189
+ 1.791e+11Hz -0.00115878 -0.00306737
+ 1.792e+11Hz -0.00114971 -0.00311276
+ 1.793e+11Hz -0.00114076 -0.00315808
+ 1.794e+11Hz -0.00113192 -0.00320332
+ 1.795e+11Hz -0.00112319 -0.00324849
+ 1.796e+11Hz -0.00111457 -0.00329357
+ 1.797e+11Hz -0.00110607 -0.00333858
+ 1.798e+11Hz -0.00109767 -0.00338351
+ 1.799e+11Hz -0.00108939 -0.00342836
+ 1.8e+11Hz -0.00108121 -0.00347313
+ 1.801e+11Hz -0.00107313 -0.00351782
+ 1.802e+11Hz -0.00106517 -0.00356244
+ 1.803e+11Hz -0.00105731 -0.00360698
+ 1.804e+11Hz -0.00104955 -0.00365144
+ 1.805e+11Hz -0.0010419 -0.00369582
+ 1.806e+11Hz -0.00103435 -0.00374012
+ 1.807e+11Hz -0.0010269 -0.00378435
+ 1.808e+11Hz -0.00101955 -0.00382849
+ 1.809e+11Hz -0.00101231 -0.00387256
+ 1.81e+11Hz -0.00100516 -0.00391655
+ 1.811e+11Hz -0.000998105 -0.00396045
+ 1.812e+11Hz -0.000991151 -0.00400428
+ 1.813e+11Hz -0.000984293 -0.00404803
+ 1.814e+11Hz -0.00097753 -0.00409169
+ 1.815e+11Hz -0.000970861 -0.00413528
+ 1.816e+11Hz -0.000964285 -0.00417878
+ 1.817e+11Hz -0.0009578 -0.0042222
+ 1.818e+11Hz -0.000951406 -0.00426554
+ 1.819e+11Hz -0.000945102 -0.00430879
+ 1.82e+11Hz -0.000938886 -0.00435196
+ 1.821e+11Hz -0.000932757 -0.00439504
+ 1.822e+11Hz -0.000926714 -0.00443804
+ 1.823e+11Hz -0.000920755 -0.00448096
+ 1.824e+11Hz -0.00091488 -0.00452379
+ 1.825e+11Hz -0.000909087 -0.00456653
+ 1.826e+11Hz -0.000903374 -0.00460919
+ 1.827e+11Hz -0.00089774 -0.00465175
+ 1.828e+11Hz -0.000892183 -0.00469423
+ 1.829e+11Hz -0.000886702 -0.00473662
+ 1.83e+11Hz -0.000881296 -0.00477892
+ 1.831e+11Hz -0.000875962 -0.00482112
+ 1.832e+11Hz -0.000870698 -0.00486324
+ 1.833e+11Hz -0.000865504 -0.00490526
+ 1.834e+11Hz -0.000860377 -0.00494719
+ 1.835e+11Hz -0.000855315 -0.00498903
+ 1.836e+11Hz -0.000850316 -0.00503077
+ 1.837e+11Hz -0.000845378 -0.00507242
+ 1.838e+11Hz -0.000840499 -0.00511397
+ 1.839e+11Hz -0.000835677 -0.00515542
+ 1.84e+11Hz -0.00083091 -0.00519678
+ 1.841e+11Hz -0.000826195 -0.00523804
+ 1.842e+11Hz -0.00082153 -0.0052792
+ 1.843e+11Hz -0.000816912 -0.00532027
+ 1.844e+11Hz -0.000812339 -0.00536123
+ 1.845e+11Hz -0.000807809 -0.0054021
+ 1.846e+11Hz -0.000803318 -0.00544286
+ 1.847e+11Hz -0.000798863 -0.00548352
+ 1.848e+11Hz -0.000794443 -0.00552409
+ 1.849e+11Hz -0.000790054 -0.00556455
+ 1.85e+11Hz -0.000785694 -0.00560491
+ 1.851e+11Hz -0.000781358 -0.00564516
+ 1.852e+11Hz -0.000777045 -0.00568532
+ 1.853e+11Hz -0.00077275 -0.00572537
+ 1.854e+11Hz -0.000768471 -0.00576532
+ 1.855e+11Hz -0.000764205 -0.00580517
+ 1.856e+11Hz -0.000759947 -0.00584492
+ 1.857e+11Hz -0.000755695 -0.00588456
+ 1.858e+11Hz -0.000751445 -0.00592411
+ 1.859e+11Hz -0.000747193 -0.00596355
+ 1.86e+11Hz -0.000742937 -0.00600289
+ 1.861e+11Hz -0.000738671 -0.00604213
+ 1.862e+11Hz -0.000734393 -0.00608127
+ 1.863e+11Hz -0.000730098 -0.00612031
+ 1.864e+11Hz -0.000725782 -0.00615926
+ 1.865e+11Hz -0.000721443 -0.0061981
+ 1.866e+11Hz -0.000717075 -0.00623685
+ 1.867e+11Hz -0.000712675 -0.0062755
+ 1.868e+11Hz -0.000708239 -0.00631406
+ 1.869e+11Hz -0.000703762 -0.00635253
+ 1.87e+11Hz -0.00069924 -0.00639091
+ 1.871e+11Hz -0.00069467 -0.00642919
+ 1.872e+11Hz -0.000690046 -0.00646739
+ 1.873e+11Hz -0.000685366 -0.0065055
+ 1.874e+11Hz -0.000680623 -0.00654353
+ 1.875e+11Hz -0.000675815 -0.00658148
+ 1.876e+11Hz -0.000670937 -0.00661934
+ 1.877e+11Hz -0.000665984 -0.00665713
+ 1.878e+11Hz -0.000660953 -0.00669485
+ 1.879e+11Hz -0.000655838 -0.00673249
+ 1.88e+11Hz -0.000650635 -0.00677006
+ 1.881e+11Hz -0.000645341 -0.00680757
+ 1.882e+11Hz -0.00063995 -0.00684501
+ 1.883e+11Hz -0.000634459 -0.0068824
+ 1.884e+11Hz -0.000628863 -0.00691972
+ 1.885e+11Hz -0.000623158 -0.006957
+ 1.886e+11Hz -0.000617339 -0.00699422
+ 1.887e+11Hz -0.000611403 -0.0070314
+ 1.888e+11Hz -0.000605345 -0.00706854
+ 1.889e+11Hz -0.000599161 -0.00710565
+ 1.89e+11Hz -0.000592846 -0.00714272
+ 1.891e+11Hz -0.000586398 -0.00717976
+ 1.892e+11Hz -0.000579811 -0.00721678
+ 1.893e+11Hz -0.000573083 -0.00725379
+ 1.894e+11Hz -0.000566208 -0.00729078
+ 1.895e+11Hz -0.000559184 -0.00732776
+ 1.896e+11Hz -0.000552006 -0.00736474
+ 1.897e+11Hz -0.000544672 -0.00740172
+ 1.898e+11Hz -0.000537177 -0.00743871
+ 1.899e+11Hz -0.000529518 -0.00747572
+ 1.9e+11Hz -0.000521692 -0.00751275
+ 1.901e+11Hz -0.000513695 -0.00754981
+ 1.902e+11Hz -0.000505526 -0.0075869
+ 1.903e+11Hz -0.000497179 -0.00762403
+ 1.904e+11Hz -0.000488654 -0.00766121
+ 1.905e+11Hz -0.000479946 -0.00769844
+ 1.906e+11Hz -0.000471055 -0.00773573
+ 1.907e+11Hz -0.000461976 -0.00777309
+ 1.908e+11Hz -0.000452709 -0.00781053
+ 1.909e+11Hz -0.00044325 -0.00784804
+ 1.91e+11Hz -0.000433599 -0.00788565
+ 1.911e+11Hz -0.000423752 -0.00792336
+ 1.912e+11Hz -0.00041371 -0.00796118
+ 1.913e+11Hz -0.00040347 -0.0079991
+ 1.914e+11Hz -0.000393031 -0.00803715
+ 1.915e+11Hz -0.000382392 -0.00807533
+ 1.916e+11Hz -0.000371553 -0.00811365
+ 1.917e+11Hz -0.000360512 -0.00815212
+ 1.918e+11Hz -0.00034927 -0.00819074
+ 1.919e+11Hz -0.000337826 -0.00822953
+ 1.92e+11Hz -0.000326181 -0.00826849
+ 1.921e+11Hz -0.000314334 -0.00830763
+ 1.922e+11Hz -0.000302287 -0.00834696
+ 1.923e+11Hz -0.000290039 -0.0083865
+ 1.924e+11Hz -0.000277593 -0.00842624
+ 1.925e+11Hz -0.000264948 -0.0084662
+ 1.926e+11Hz -0.000252108 -0.00850639
+ 1.927e+11Hz -0.000239073 -0.00854681
+ 1.928e+11Hz -0.000225845 -0.00858749
+ 1.929e+11Hz -0.000212427 -0.00862841
+ 1.93e+11Hz -0.000198821 -0.00866961
+ 1.931e+11Hz -0.00018503 -0.00871107
+ 1.932e+11Hz -0.000171057 -0.00875283
+ 1.933e+11Hz -0.000156906 -0.00879487
+ 1.934e+11Hz -0.000142579 -0.00883722
+ 1.935e+11Hz -0.000128082 -0.00887988
+ 1.936e+11Hz -0.000113417 -0.00892286
+ 1.937e+11Hz -9.85897e-05 -0.00896617
+ 1.938e+11Hz -8.36045e-05 -0.00900983
+ 1.939e+11Hz -6.84665e-05 -0.00905383
+ 1.94e+11Hz -5.31808e-05 -0.00909819
+ 1.941e+11Hz -3.77531e-05 -0.00914293
+ 1.942e+11Hz -2.21892e-05 -0.00918804
+ 1.943e+11Hz -6.49523e-06 -0.00923353
+ 1.944e+11Hz 9.3224e-06 -0.00927943
+ 1.945e+11Hz 2.5257e-05 -0.00932573
+ 1.946e+11Hz 4.13015e-05 -0.00937244
+ 1.947e+11Hz 5.74487e-05 -0.00941957
+ 1.948e+11Hz 7.36911e-05 -0.00946714
+ 1.949e+11Hz 9.00207e-05 -0.00951515
+ 1.95e+11Hz 0.00010643 -0.0095636
+ 1.951e+11Hz 0.000122909 -0.00961251
+ 1.952e+11Hz 0.000139451 -0.00966189
+ 1.953e+11Hz 0.000156046 -0.00971174
+ 1.954e+11Hz 0.000172684 -0.00976207
+ 1.955e+11Hz 0.000189358 -0.00981289
+ 1.956e+11Hz 0.000206056 -0.00986421
+ 1.957e+11Hz 0.000222768 -0.00991602
+ 1.958e+11Hz 0.000239485 -0.00996835
+ 1.959e+11Hz 0.000256196 -0.0100212
+ 1.96e+11Hz 0.00027289 -0.0100746
+ 1.961e+11Hz 0.000289556 -0.0101285
+ 1.962e+11Hz 0.000306183 -0.0101829
+ 1.963e+11Hz 0.000322759 -0.0102379
+ 1.964e+11Hz 0.000339273 -0.0102934
+ 1.965e+11Hz 0.000355713 -0.0103495
+ 1.966e+11Hz 0.000372066 -0.0104061
+ 1.967e+11Hz 0.00038832 -0.0104633
+ 1.968e+11Hz 0.000404462 -0.0105211
+ 1.969e+11Hz 0.000420481 -0.0105794
+ 1.97e+11Hz 0.000436362 -0.0106383
+ 1.971e+11Hz 0.000452092 -0.0106978
+ 1.972e+11Hz 0.000467659 -0.0107579
+ 1.973e+11Hz 0.000483049 -0.0108186
+ 1.974e+11Hz 0.000498248 -0.0108798
+ 1.975e+11Hz 0.000513242 -0.0109417
+ 1.976e+11Hz 0.000528018 -0.0110041
+ 1.977e+11Hz 0.000542561 -0.0110672
+ 1.978e+11Hz 0.000556857 -0.0111308
+ 1.979e+11Hz 0.000570891 -0.011195
+ 1.98e+11Hz 0.00058465 -0.0112599
+ 1.981e+11Hz 0.000598119 -0.0113253
+ 1.982e+11Hz 0.000611282 -0.0113913
+ 1.983e+11Hz 0.000624126 -0.0114579
+ 1.984e+11Hz 0.000636636 -0.0115252
+ 1.985e+11Hz 0.000648796 -0.011593
+ 1.986e+11Hz 0.000660592 -0.0116614
+ 1.987e+11Hz 0.000672009 -0.0117304
+ 1.988e+11Hz 0.000683032 -0.0118001
+ 1.989e+11Hz 0.000693646 -0.0118702
+ 1.99e+11Hz 0.000703835 -0.011941
+ 1.991e+11Hz 0.000713586 -0.0120124
+ 1.992e+11Hz 0.000722882 -0.0120843
+ 1.993e+11Hz 0.00073171 -0.0121569
+ 1.994e+11Hz 0.000740054 -0.01223
+ 1.995e+11Hz 0.000747898 -0.0123036
+ 1.996e+11Hz 0.00075523 -0.0123778
+ 1.997e+11Hz 0.000762032 -0.0124526
+ 1.998e+11Hz 0.000768292 -0.0125279
+ 1.999e+11Hz 0.000773994 -0.0126038
+ 2e+11Hz 0.000779124 -0.0126802
+ 2.001e+11Hz 0.000783668 -0.0127571
+ 2.002e+11Hz 0.00078761 -0.0128346
+ 2.003e+11Hz 0.000790938 -0.0129125
+ 2.004e+11Hz 0.000793637 -0.012991
+ 2.005e+11Hz 0.000795693 -0.01307
+ 2.006e+11Hz 0.000797093 -0.0131494
+ 2.007e+11Hz 0.000797823 -0.0132293
+ 2.008e+11Hz 0.00079787 -0.0133097
+ 2.009e+11Hz 0.000797221 -0.0133906
+ 2.01e+11Hz 0.000795862 -0.0134719
+ 2.011e+11Hz 0.000793782 -0.0135536
+ 2.012e+11Hz 0.000790968 -0.0136358
+ 2.013e+11Hz 0.000787407 -0.0137183
+ 2.014e+11Hz 0.000783088 -0.0138013
+ 2.015e+11Hz 0.000777999 -0.0138846
+ 2.016e+11Hz 0.000772129 -0.0139684
+ 2.017e+11Hz 0.000765466 -0.0140525
+ 2.018e+11Hz 0.000757999 -0.0141369
+ 2.019e+11Hz 0.000749719 -0.0142217
+ 2.02e+11Hz 0.000740614 -0.0143068
+ 2.021e+11Hz 0.000730675 -0.0143922
+ 2.022e+11Hz 0.000719892 -0.0144779
+ 2.023e+11Hz 0.000708256 -0.0145638
+ 2.024e+11Hz 0.000695758 -0.0146501
+ 2.025e+11Hz 0.000682389 -0.0147366
+ 2.026e+11Hz 0.000668141 -0.0148233
+ 2.027e+11Hz 0.000653007 -0.0149102
+ 2.028e+11Hz 0.000636978 -0.0149974
+ 2.029e+11Hz 0.000620048 -0.0150847
+ 2.03e+11Hz 0.000602209 -0.0151722
+ 2.031e+11Hz 0.000583456 -0.0152598
+ 2.032e+11Hz 0.000563782 -0.0153476
+ 2.033e+11Hz 0.000543182 -0.0154355
+ 2.034e+11Hz 0.00052165 -0.0155235
+ 2.035e+11Hz 0.000499182 -0.0156116
+ 2.036e+11Hz 0.000475774 -0.0156997
+ 2.037e+11Hz 0.000451421 -0.0157879
+ 2.038e+11Hz 0.00042612 -0.0158762
+ 2.039e+11Hz 0.000399868 -0.0159644
+ 2.04e+11Hz 0.000372661 -0.0160527
+ 2.041e+11Hz 0.000344499 -0.0161409
+ 2.042e+11Hz 0.000315379 -0.0162291
+ 2.043e+11Hz 0.000285299 -0.0163172
+ 2.044e+11Hz 0.00025426 -0.0164053
+ 2.045e+11Hz 0.000222259 -0.0164933
+ 2.046e+11Hz 0.000189297 -0.0165811
+ 2.047e+11Hz 0.000155375 -0.0166688
+ 2.048e+11Hz 0.000120493 -0.0167564
+ 2.049e+11Hz 8.46531e-05 -0.0168438
+ 2.05e+11Hz 4.78559e-05 -0.0169311
+ 2.051e+11Hz 1.0104e-05 -0.0170181
+ 2.052e+11Hz -2.86e-05 -0.0171049
+ 2.053e+11Hz -6.82532e-05 -0.0171915
+ 2.054e+11Hz -0.000108852 -0.0172778
+ 2.055e+11Hz -0.000150393 -0.0173638
+ 2.056e+11Hz -0.000192871 -0.0174496
+ 2.057e+11Hz -0.000236283 -0.017535
+ 2.058e+11Hz -0.000280622 -0.0176202
+ 2.059e+11Hz -0.000325883 -0.0177049
+ 2.06e+11Hz -0.00037206 -0.0177894
+ 2.061e+11Hz -0.000419148 -0.0178734
+ 2.062e+11Hz -0.000467138 -0.0179571
+ 2.063e+11Hz -0.000516025 -0.0180403
+ 2.064e+11Hz -0.000565799 -0.0181231
+ 2.065e+11Hz -0.000616454 -0.0182055
+ 2.066e+11Hz -0.000667981 -0.0182874
+ 2.067e+11Hz -0.000720371 -0.0183689
+ 2.068e+11Hz -0.000773616 -0.0184498
+ 2.069e+11Hz -0.000827705 -0.0185303
+ 2.07e+11Hz -0.000882628 -0.0186102
+ 2.071e+11Hz -0.000938377 -0.0186896
+ 2.072e+11Hz -0.000994939 -0.0187684
+ 2.073e+11Hz -0.00105231 -0.0188467
+ 2.074e+11Hz -0.00111046 -0.0189244
+ 2.075e+11Hz -0.0011694 -0.0190015
+ 2.076e+11Hz -0.00122911 -0.019078
+ 2.077e+11Hz -0.00128957 -0.0191539
+ 2.078e+11Hz -0.00135078 -0.0192291
+ 2.079e+11Hz -0.00141272 -0.0193038
+ 2.08e+11Hz -0.00147538 -0.0193777
+ 2.081e+11Hz -0.00153874 -0.019451
+ 2.082e+11Hz -0.0016028 -0.0195236
+ 2.083e+11Hz -0.00166753 -0.0195955
+ 2.084e+11Hz -0.00173293 -0.0196668
+ 2.085e+11Hz -0.00179898 -0.0197373
+ 2.086e+11Hz -0.00186566 -0.0198071
+ 2.087e+11Hz -0.00193297 -0.0198761
+ 2.088e+11Hz -0.00200088 -0.0199444
+ 2.089e+11Hz -0.00206938 -0.020012
+ 2.09e+11Hz -0.00213846 -0.0200788
+ 2.091e+11Hz -0.0022081 -0.0201449
+ 2.092e+11Hz -0.00227828 -0.0202101
+ 2.093e+11Hz -0.002349 -0.0202746
+ 2.094e+11Hz -0.00242023 -0.0203384
+ 2.095e+11Hz -0.00249196 -0.0204013
+ 2.096e+11Hz -0.00256417 -0.0204634
+ 2.097e+11Hz -0.00263684 -0.0205247
+ 2.098e+11Hz -0.00270997 -0.0205852
+ 2.099e+11Hz -0.00278353 -0.0206449
+ 2.1e+11Hz -0.00285752 -0.0207038
+ 2.101e+11Hz -0.0029319 -0.0207618
+ 2.102e+11Hz -0.00300667 -0.020819
+ 2.103e+11Hz -0.00308181 -0.0208754
+ 2.104e+11Hz -0.0031573 -0.020931
+ 2.105e+11Hz -0.00323313 -0.0209857
+ 2.106e+11Hz -0.00330928 -0.0210396
+ 2.107e+11Hz -0.00338574 -0.0210926
+ 2.108e+11Hz -0.00346248 -0.0211448
+ 2.109e+11Hz -0.00353949 -0.0211962
+ 2.11e+11Hz -0.00361677 -0.0212467
+ 2.111e+11Hz -0.00369428 -0.0212964
+ 2.112e+11Hz -0.00377202 -0.0213452
+ 2.113e+11Hz -0.00384996 -0.0213932
+ 2.114e+11Hz -0.0039281 -0.0214404
+ 2.115e+11Hz -0.00400642 -0.0214867
+ 2.116e+11Hz -0.00408489 -0.0215322
+ 2.117e+11Hz -0.00416352 -0.0215768
+ 2.118e+11Hz -0.00424227 -0.0216207
+ 2.119e+11Hz -0.00432114 -0.0216637
+ 2.12e+11Hz -0.00440011 -0.0217058
+ 2.121e+11Hz -0.00447917 -0.0217472
+ 2.122e+11Hz -0.0045583 -0.0217877
+ 2.123e+11Hz -0.00463749 -0.0218274
+ 2.124e+11Hz -0.00471672 -0.0218663
+ 2.125e+11Hz -0.00479598 -0.0219044
+ 2.126e+11Hz -0.00487525 -0.0219417
+ 2.127e+11Hz -0.00495453 -0.0219782
+ 2.128e+11Hz -0.00503379 -0.0220139
+ 2.129e+11Hz -0.00511303 -0.0220488
+ 2.13e+11Hz -0.00519223 -0.022083
+ 2.131e+11Hz -0.00527138 -0.0221164
+ 2.132e+11Hz -0.00535046 -0.022149
+ 2.133e+11Hz -0.00542947 -0.0221809
+ 2.134e+11Hz -0.0055084 -0.022212
+ 2.135e+11Hz -0.00558722 -0.0222424
+ 2.136e+11Hz -0.00566593 -0.0222721
+ 2.137e+11Hz -0.00574453 -0.022301
+ 2.138e+11Hz -0.00582299 -0.0223292
+ 2.139e+11Hz -0.0059013 -0.0223567
+ 2.14e+11Hz -0.00597946 -0.0223835
+ 2.141e+11Hz -0.00605746 -0.0224096
+ 2.142e+11Hz -0.00613529 -0.022435
+ 2.143e+11Hz -0.00621293 -0.0224598
+ 2.144e+11Hz -0.00629038 -0.0224839
+ 2.145e+11Hz -0.00636763 -0.0225073
+ 2.146e+11Hz -0.00644467 -0.0225301
+ 2.147e+11Hz -0.00652149 -0.0225523
+ 2.148e+11Hz -0.00659808 -0.0225738
+ 2.149e+11Hz -0.00667445 -0.0225947
+ 2.15e+11Hz -0.00675057 -0.022615
+ 2.151e+11Hz -0.00682644 -0.0226347
+ 2.152e+11Hz -0.00690205 -0.0226539
+ 2.153e+11Hz -0.00697741 -0.0226724
+ 2.154e+11Hz -0.00705249 -0.0226904
+ 2.155e+11Hz -0.0071273 -0.0227078
+ 2.156e+11Hz -0.00720184 -0.0227247
+ 2.157e+11Hz -0.00727608 -0.0227411
+ 2.158e+11Hz -0.00735004 -0.0227569
+ 2.159e+11Hz -0.0074237 -0.0227722
+ 2.16e+11Hz -0.00749706 -0.022787
+ 2.161e+11Hz -0.00757012 -0.0228013
+ 2.162e+11Hz -0.00764286 -0.0228151
+ 2.163e+11Hz -0.0077153 -0.0228285
+ 2.164e+11Hz -0.00778742 -0.0228414
+ 2.165e+11Hz -0.00785922 -0.0228538
+ 2.166e+11Hz -0.0079307 -0.0228658
+ 2.167e+11Hz -0.00800186 -0.0228774
+ 2.168e+11Hz -0.00807269 -0.0228885
+ 2.169e+11Hz -0.00814319 -0.0228993
+ 2.17e+11Hz -0.00821337 -0.0229096
+ 2.171e+11Hz -0.0082832 -0.0229196
+ 2.172e+11Hz -0.00835271 -0.0229291
+ 2.173e+11Hz -0.00842188 -0.0229383
+ 2.174e+11Hz -0.00849071 -0.0229471
+ 2.175e+11Hz -0.00855921 -0.0229556
+ 2.176e+11Hz -0.00862737 -0.0229637
+ 2.177e+11Hz -0.00869519 -0.0229715
+ 2.178e+11Hz -0.00876268 -0.022979
+ 2.179e+11Hz -0.00882982 -0.0229862
+ 2.18e+11Hz -0.00889663 -0.022993
+ 2.181e+11Hz -0.00896311 -0.0229996
+ 2.182e+11Hz -0.00902924 -0.0230058
+ 2.183e+11Hz -0.00909504 -0.0230118
+ 2.184e+11Hz -0.00916051 -0.0230176
+ 2.185e+11Hz -0.00922564 -0.023023
+ 2.186e+11Hz -0.00929044 -0.0230282
+ 2.187e+11Hz -0.00935491 -0.0230332
+ 2.188e+11Hz -0.00941905 -0.0230379
+ 2.189e+11Hz -0.00948286 -0.0230424
+ 2.19e+11Hz -0.00954635 -0.0230467
+ 2.191e+11Hz -0.00960952 -0.0230508
+ 2.192e+11Hz -0.00967236 -0.0230546
+ 2.193e+11Hz -0.00973488 -0.0230583
+ 2.194e+11Hz -0.00979709 -0.0230618
+ 2.195e+11Hz -0.00985898 -0.023065
+ 2.196e+11Hz -0.00992057 -0.0230682
+ 2.197e+11Hz -0.00998184 -0.0230711
+ 2.198e+11Hz -0.0100428 -0.0230739
+ 2.199e+11Hz -0.0101035 -0.0230765
+ 2.2e+11Hz -0.0101638 -0.023079
+ 2.201e+11Hz -0.0102239 -0.0230813
+ 2.202e+11Hz -0.0102837 -0.0230835
+ 2.203e+11Hz -0.0103432 -0.0230856
+ 2.204e+11Hz -0.0104023 -0.0230876
+ 2.205e+11Hz -0.0104613 -0.0230894
+ 2.206e+11Hz -0.0105199 -0.0230911
+ 2.207e+11Hz -0.0105782 -0.0230927
+ 2.208e+11Hz -0.0106363 -0.0230942
+ 2.209e+11Hz -0.0106941 -0.0230957
+ 2.21e+11Hz -0.0107516 -0.023097
+ 2.211e+11Hz -0.0108089 -0.0230982
+ 2.212e+11Hz -0.0108659 -0.0230994
+ 2.213e+11Hz -0.0109227 -0.0231005
+ 2.214e+11Hz -0.0109792 -0.0231015
+ 2.215e+11Hz -0.0110355 -0.0231025
+ 2.216e+11Hz -0.0110915 -0.0231033
+ 2.217e+11Hz -0.0111472 -0.0231042
+ 2.218e+11Hz -0.0112028 -0.023105
+ 2.219e+11Hz -0.0112581 -0.0231057
+ 2.22e+11Hz -0.0113131 -0.0231064
+ 2.221e+11Hz -0.011368 -0.0231071
+ 2.222e+11Hz -0.0114226 -0.0231077
+ 2.223e+11Hz -0.011477 -0.0231083
+ 2.224e+11Hz -0.0115311 -0.0231088
+ 2.225e+11Hz -0.0115851 -0.0231094
+ 2.226e+11Hz -0.0116389 -0.0231099
+ 2.227e+11Hz -0.0116924 -0.0231104
+ 2.228e+11Hz -0.0117458 -0.0231109
+ 2.229e+11Hz -0.0117989 -0.0231114
+ 2.23e+11Hz -0.0118519 -0.0231119
+ 2.231e+11Hz -0.0119047 -0.0231124
+ 2.232e+11Hz -0.0119573 -0.0231129
+ 2.233e+11Hz -0.0120097 -0.0231134
+ 2.234e+11Hz -0.0120619 -0.0231139
+ 2.235e+11Hz -0.012114 -0.0231144
+ 2.236e+11Hz -0.0121659 -0.0231149
+ 2.237e+11Hz -0.0122176 -0.0231155
+ 2.238e+11Hz -0.0122692 -0.023116
+ 2.239e+11Hz -0.0123206 -0.0231166
+ 2.24e+11Hz -0.0123718 -0.0231173
+ 2.241e+11Hz -0.0124229 -0.0231179
+ 2.242e+11Hz -0.0124739 -0.0231186
+ 2.243e+11Hz -0.0125247 -0.0231194
+ 2.244e+11Hz -0.0125754 -0.0231201
+ 2.245e+11Hz -0.0126259 -0.0231209
+ 2.246e+11Hz -0.0126763 -0.0231218
+ 2.247e+11Hz -0.0127266 -0.0231227
+ 2.248e+11Hz -0.0127768 -0.0231237
+ 2.249e+11Hz -0.0128268 -0.0231247
+ 2.25e+11Hz -0.0128768 -0.0231258
+ 2.251e+11Hz -0.0129266 -0.0231269
+ 2.252e+11Hz -0.0129763 -0.0231282
+ 2.253e+11Hz -0.013026 -0.0231294
+ 2.254e+11Hz -0.0130755 -0.0231308
+ 2.255e+11Hz -0.013125 -0.0231322
+ 2.256e+11Hz -0.0131743 -0.0231337
+ 2.257e+11Hz -0.0132236 -0.0231353
+ 2.258e+11Hz -0.0132728 -0.0231369
+ 2.259e+11Hz -0.0133219 -0.0231386
+ 2.26e+11Hz -0.013371 -0.0231405
+ 2.261e+11Hz -0.01342 -0.0231424
+ 2.262e+11Hz -0.0134689 -0.0231444
+ 2.263e+11Hz -0.0135178 -0.0231465
+ 2.264e+11Hz -0.0135667 -0.0231487
+ 2.265e+11Hz -0.0136155 -0.023151
+ 2.266e+11Hz -0.0136642 -0.0231534
+ 2.267e+11Hz -0.013713 -0.0231558
+ 2.268e+11Hz -0.0137617 -0.0231584
+ 2.269e+11Hz -0.0138104 -0.0231612
+ 2.27e+11Hz -0.0138591 -0.023164
+ 2.271e+11Hz -0.0139078 -0.0231669
+ 2.272e+11Hz -0.0139564 -0.02317
+ 2.273e+11Hz -0.0140051 -0.0231731
+ 2.274e+11Hz -0.0140538 -0.0231764
+ 2.275e+11Hz -0.0141025 -0.0231798
+ 2.276e+11Hz -0.0141513 -0.0231833
+ 2.277e+11Hz -0.0142 -0.023187
+ 2.278e+11Hz -0.0142488 -0.0231908
+ 2.279e+11Hz -0.0142977 -0.0231947
+ 2.28e+11Hz -0.0143466 -0.0231987
+ 2.281e+11Hz -0.0143956 -0.0232028
+ 2.282e+11Hz -0.0144446 -0.0232071
+ 2.283e+11Hz -0.0144937 -0.0232115
+ 2.284e+11Hz -0.0145429 -0.0232161
+ 2.285e+11Hz -0.0145922 -0.0232208
+ 2.286e+11Hz -0.0146415 -0.0232256
+ 2.287e+11Hz -0.014691 -0.0232306
+ 2.288e+11Hz -0.0147406 -0.0232356
+ 2.289e+11Hz -0.0147903 -0.0232409
+ 2.29e+11Hz -0.0148402 -0.0232462
+ 2.291e+11Hz -0.0148901 -0.0232517
+ 2.292e+11Hz -0.0149402 -0.0232573
+ 2.293e+11Hz -0.0149905 -0.0232631
+ 2.294e+11Hz -0.015041 -0.023269
+ 2.295e+11Hz -0.0150916 -0.023275
+ 2.296e+11Hz -0.0151424 -0.0232812
+ 2.297e+11Hz -0.0151933 -0.0232875
+ 2.298e+11Hz -0.0152445 -0.0232939
+ 2.299e+11Hz -0.0152959 -0.0233004
+ 2.3e+11Hz -0.0153475 -0.0233071
+ 2.301e+11Hz -0.0153993 -0.0233139
+ 2.302e+11Hz -0.0154514 -0.0233208
+ 2.303e+11Hz -0.0155037 -0.0233278
+ 2.304e+11Hz -0.0155562 -0.0233349
+ 2.305e+11Hz -0.015609 -0.0233422
+ 2.306e+11Hz -0.0156621 -0.0233495
+ 2.307e+11Hz -0.0157155 -0.0233569
+ 2.308e+11Hz -0.0157692 -0.0233645
+ 2.309e+11Hz -0.0158231 -0.0233721
+ 2.31e+11Hz -0.0158774 -0.0233799
+ 2.311e+11Hz -0.015932 -0.0233877
+ 2.312e+11Hz -0.0159869 -0.0233956
+ 2.313e+11Hz -0.0160422 -0.0234036
+ 2.314e+11Hz -0.0160978 -0.0234116
+ 2.315e+11Hz -0.0161538 -0.0234197
+ 2.316e+11Hz -0.0162102 -0.0234278
+ 2.317e+11Hz -0.0162669 -0.023436
+ 2.318e+11Hz -0.016324 -0.0234443
+ 2.319e+11Hz -0.0163815 -0.0234526
+ 2.32e+11Hz -0.0164394 -0.0234609
+ 2.321e+11Hz -0.0164978 -0.0234692
+ 2.322e+11Hz -0.0165565 -0.0234775
+ 2.323e+11Hz -0.0166157 -0.0234858
+ 2.324e+11Hz -0.0166754 -0.0234942
+ 2.325e+11Hz -0.0167355 -0.0235025
+ 2.326e+11Hz -0.016796 -0.0235107
+ 2.327e+11Hz -0.016857 -0.023519
+ 2.328e+11Hz -0.0169185 -0.0235271
+ 2.329e+11Hz -0.0169805 -0.0235353
+ 2.33e+11Hz -0.017043 -0.0235433
+ 2.331e+11Hz -0.017106 -0.0235513
+ 2.332e+11Hz -0.0171695 -0.0235592
+ 2.333e+11Hz -0.0172335 -0.023567
+ 2.334e+11Hz -0.0172981 -0.0235746
+ 2.335e+11Hz -0.0173631 -0.0235821
+ 2.336e+11Hz -0.0174288 -0.0235895
+ 2.337e+11Hz -0.0174949 -0.0235968
+ 2.338e+11Hz -0.0175616 -0.0236038
+ 2.339e+11Hz -0.0176289 -0.0236107
+ 2.34e+11Hz -0.0176968 -0.0236173
+ 2.341e+11Hz -0.0177652 -0.0236238
+ 2.342e+11Hz -0.0178341 -0.02363
+ 2.343e+11Hz -0.0179037 -0.023636
+ 2.344e+11Hz -0.0179738 -0.0236417
+ 2.345e+11Hz -0.0180446 -0.0236472
+ 2.346e+11Hz -0.0181159 -0.0236523
+ 2.347e+11Hz -0.0181878 -0.0236572
+ 2.348e+11Hz -0.0182604 -0.0236617
+ 2.349e+11Hz -0.0183335 -0.0236659
+ 2.35e+11Hz -0.0184072 -0.0236697
+ 2.351e+11Hz -0.0184815 -0.0236732
+ 2.352e+11Hz -0.0185565 -0.0236762
+ 2.353e+11Hz -0.018632 -0.0236789
+ 2.354e+11Hz -0.0187082 -0.0236811
+ 2.355e+11Hz -0.0187849 -0.0236829
+ 2.356e+11Hz -0.0188623 -0.0236842
+ 2.357e+11Hz -0.0189402 -0.023685
+ 2.358e+11Hz -0.0190188 -0.0236854
+ 2.359e+11Hz -0.019098 -0.0236852
+ 2.36e+11Hz -0.0191778 -0.0236844
+ 2.361e+11Hz -0.0192582 -0.0236832
+ 2.362e+11Hz -0.0193391 -0.0236813
+ 2.363e+11Hz -0.0194207 -0.0236788
+ 2.364e+11Hz -0.0195028 -0.0236758
+ 2.365e+11Hz -0.0195856 -0.0236721
+ 2.366e+11Hz -0.0196689 -0.0236677
+ 2.367e+11Hz -0.0197528 -0.0236627
+ 2.368e+11Hz -0.0198372 -0.023657
+ 2.369e+11Hz -0.0199222 -0.0236506
+ 2.37e+11Hz -0.0200077 -0.0236434
+ 2.371e+11Hz -0.0200938 -0.0236355
+ 2.372e+11Hz -0.0201804 -0.0236269
+ 2.373e+11Hz -0.0202676 -0.0236174
+ 2.374e+11Hz -0.0203552 -0.0236071
+ 2.375e+11Hz -0.0204434 -0.0235961
+ 2.376e+11Hz -0.020532 -0.0235841
+ 2.377e+11Hz -0.0206211 -0.0235714
+ 2.378e+11Hz -0.0207107 -0.0235577
+ 2.379e+11Hz -0.0208008 -0.0235431
+ 2.38e+11Hz -0.0208913 -0.0235277
+ 2.381e+11Hz -0.0209822 -0.0235113
+ 2.382e+11Hz -0.0210735 -0.0234939
+ 2.383e+11Hz -0.0211652 -0.0234756
+ 2.384e+11Hz -0.0212573 -0.0234563
+ 2.385e+11Hz -0.0213498 -0.023436
+ 2.386e+11Hz -0.0214426 -0.0234147
+ 2.387e+11Hz -0.0215358 -0.0233923
+ 2.388e+11Hz -0.0216293 -0.0233689
+ 2.389e+11Hz -0.021723 -0.0233444
+ 2.39e+11Hz -0.0218171 -0.0233189
+ 2.391e+11Hz -0.0219114 -0.0232922
+ 2.392e+11Hz -0.0220059 -0.0232645
+ 2.393e+11Hz -0.0221007 -0.0232356
+ 2.394e+11Hz -0.0221957 -0.0232056
+ 2.395e+11Hz -0.0222908 -0.0231744
+ 2.396e+11Hz -0.0223861 -0.0231421
+ 2.397e+11Hz -0.0224816 -0.0231086
+ 2.398e+11Hz -0.0225771 -0.0230739
+ 2.399e+11Hz -0.0226727 -0.023038
+ 2.4e+11Hz -0.0227684 -0.0230009
+ 2.401e+11Hz -0.0228642 -0.0229626
+ 2.402e+11Hz -0.02296 -0.022923
+ 2.403e+11Hz -0.0230557 -0.0228823
+ 2.404e+11Hz -0.0231514 -0.0228403
+ 2.405e+11Hz -0.0232471 -0.022797
+ 2.406e+11Hz -0.0233427 -0.0227524
+ 2.407e+11Hz -0.0234382 -0.0227067
+ 2.408e+11Hz -0.0235335 -0.0226596
+ 2.409e+11Hz -0.0236287 -0.0226112
+ 2.41e+11Hz -0.0237237 -0.0225616
+ 2.411e+11Hz -0.0238185 -0.0225107
+ 2.412e+11Hz -0.023913 -0.0224585
+ 2.413e+11Hz -0.0240073 -0.022405
+ 2.414e+11Hz -0.0241013 -0.0223502
+ 2.415e+11Hz -0.024195 -0.0222941
+ 2.416e+11Hz -0.0242883 -0.0222367
+ 2.417e+11Hz -0.0243812 -0.0221781
+ 2.418e+11Hz -0.0244737 -0.0221181
+ 2.419e+11Hz -0.0245658 -0.0220568
+ 2.42e+11Hz -0.0246574 -0.0219943
+ 2.421e+11Hz -0.0247485 -0.0219305
+ 2.422e+11Hz -0.0248391 -0.0218653
+ 2.423e+11Hz -0.0249292 -0.0217989
+ 2.424e+11Hz -0.0250186 -0.0217313
+ 2.425e+11Hz -0.0251075 -0.0216623
+ 2.426e+11Hz -0.0251957 -0.0215921
+ 2.427e+11Hz -0.0252833 -0.0215207
+ 2.428e+11Hz -0.0253702 -0.021448
+ 2.429e+11Hz -0.0254563 -0.021374
+ 2.43e+11Hz -0.0255418 -0.0212989
+ 2.431e+11Hz -0.0256264 -0.0212225
+ 2.432e+11Hz -0.0257102 -0.0211449
+ 2.433e+11Hz -0.0257932 -0.0210662
+ 2.434e+11Hz -0.0258754 -0.0209862
+ 2.435e+11Hz -0.0259566 -0.0209051
+ 2.436e+11Hz -0.026037 -0.0208228
+ 2.437e+11Hz -0.0261164 -0.0207394
+ 2.438e+11Hz -0.0261948 -0.0206549
+ 2.439e+11Hz -0.0262723 -0.0205693
+ 2.44e+11Hz -0.0263487 -0.0204826
+ 2.441e+11Hz -0.0264241 -0.0203948
+ 2.442e+11Hz -0.0264985 -0.0203059
+ 2.443e+11Hz -0.0265717 -0.0202161
+ 2.444e+11Hz -0.0266439 -0.0201252
+ 2.445e+11Hz -0.0267149 -0.0200333
+ 2.446e+11Hz -0.0267847 -0.0199405
+ 2.447e+11Hz -0.0268534 -0.0198467
+ 2.448e+11Hz -0.0269208 -0.019752
+ 2.449e+11Hz -0.0269871 -0.0196564
+ 2.45e+11Hz -0.0270521 -0.0195599
+ 2.451e+11Hz -0.0271158 -0.0194625
+ 2.452e+11Hz -0.0271782 -0.0193643
+ 2.453e+11Hz -0.0272394 -0.0192653
+ 2.454e+11Hz -0.0272992 -0.0191656
+ 2.455e+11Hz -0.0273576 -0.019065
+ 2.456e+11Hz -0.0274147 -0.0189638
+ 2.457e+11Hz -0.0274705 -0.0188618
+ 2.458e+11Hz -0.0275248 -0.0187592
+ 2.459e+11Hz -0.0275778 -0.0186559
+ 2.46e+11Hz -0.0276293 -0.0185521
+ 2.461e+11Hz -0.0276794 -0.0184476
+ 2.462e+11Hz -0.0277281 -0.0183426
+ 2.463e+11Hz -0.0277752 -0.018237
+ 2.464e+11Hz -0.027821 -0.018131
+ 2.465e+11Hz -0.0278652 -0.0180244
+ 2.466e+11Hz -0.0279079 -0.0179175
+ 2.467e+11Hz -0.0279492 -0.0178101
+ 2.468e+11Hz -0.0279889 -0.0177024
+ 2.469e+11Hz -0.0280272 -0.0175943
+ 2.47e+11Hz -0.0280639 -0.0174859
+ 2.471e+11Hz -0.028099 -0.0173773
+ 2.472e+11Hz -0.0281327 -0.0172684
+ 2.473e+11Hz -0.0281648 -0.0171592
+ 2.474e+11Hz -0.0281953 -0.0170499
+ 2.475e+11Hz -0.0282243 -0.0169405
+ 2.476e+11Hz -0.0282518 -0.0168309
+ 2.477e+11Hz -0.0282777 -0.0167212
+ 2.478e+11Hz -0.0283021 -0.0166115
+ 2.479e+11Hz -0.0283249 -0.0165017
+ 2.48e+11Hz -0.0283462 -0.016392
+ 2.481e+11Hz -0.0283659 -0.0162823
+ 2.482e+11Hz -0.0283841 -0.0161727
+ 2.483e+11Hz -0.0284008 -0.0160632
+ 2.484e+11Hz -0.0284159 -0.0159539
+ 2.485e+11Hz -0.0284295 -0.0158447
+ 2.486e+11Hz -0.0284416 -0.0157357
+ 2.487e+11Hz -0.0284522 -0.015627
+ 2.488e+11Hz -0.0284612 -0.0155185
+ 2.489e+11Hz -0.0284688 -0.0154103
+ 2.49e+11Hz -0.0284749 -0.0153025
+ 2.491e+11Hz -0.0284795 -0.015195
+ 2.492e+11Hz -0.0284826 -0.0150879
+ 2.493e+11Hz -0.0284843 -0.0149812
+ 2.494e+11Hz -0.0284846 -0.014875
+ 2.495e+11Hz -0.0284834 -0.0147692
+ 2.496e+11Hz -0.0284808 -0.014664
+ 2.497e+11Hz -0.0284768 -0.0145593
+ 2.498e+11Hz -0.0284715 -0.0144551
+ 2.499e+11Hz -0.0284648 -0.0143516
+ 2.5e+11Hz -0.0284567 -0.0142487
+ 2.501e+11Hz -0.0284473 -0.0141464
+ 2.502e+11Hz -0.0284366 -0.0140448
+ 2.503e+11Hz -0.0284245 -0.0139439
+ 2.504e+11Hz -0.0284113 -0.0138437
+ 2.505e+11Hz -0.0283967 -0.0137442
+ 2.506e+11Hz -0.028381 -0.0136456
+ 2.507e+11Hz -0.028364 -0.0135477
+ 2.508e+11Hz -0.0283458 -0.0134506
+ 2.509e+11Hz -0.0283265 -0.0133544
+ 2.51e+11Hz -0.028306 -0.013259
+ 2.511e+11Hz -0.0282844 -0.0131646
+ 2.512e+11Hz -0.0282617 -0.013071
+ 2.513e+11Hz -0.028238 -0.0129783
+ 2.514e+11Hz -0.0282132 -0.0128866
+ 2.515e+11Hz -0.0281873 -0.0127958
+ 2.516e+11Hz -0.0281605 -0.012706
+ 2.517e+11Hz -0.0281327 -0.0126172
+ 2.518e+11Hz -0.028104 -0.0125295
+ 2.519e+11Hz -0.0280743 -0.0124427
+ 2.52e+11Hz -0.0280438 -0.012357
+ 2.521e+11Hz -0.0280124 -0.0122723
+ 2.522e+11Hz -0.0279802 -0.0121886
+ 2.523e+11Hz -0.0279471 -0.0121061
+ 2.524e+11Hz -0.0279133 -0.0120246
+ 2.525e+11Hz -0.0278788 -0.0119443
+ 2.526e+11Hz -0.0278435 -0.011865
+ 2.527e+11Hz -0.0278075 -0.0117869
+ 2.528e+11Hz -0.0277709 -0.0117098
+ 2.529e+11Hz -0.0277336 -0.0116339
+ 2.53e+11Hz -0.0276957 -0.0115592
+ 2.531e+11Hz -0.0276573 -0.0114856
+ 2.532e+11Hz -0.0276183 -0.0114131
+ 2.533e+11Hz -0.0275787 -0.0113418
+ 2.534e+11Hz -0.0275387 -0.0112716
+ 2.535e+11Hz -0.0274983 -0.0112026
+ 2.536e+11Hz -0.0274574 -0.0111347
+ 2.537e+11Hz -0.0274161 -0.011068
+ 2.538e+11Hz -0.0273744 -0.0110025
+ 2.539e+11Hz -0.0273324 -0.0109381
+ 2.54e+11Hz -0.02729 -0.0108749
+ 2.541e+11Hz -0.0272474 -0.0108128
+ 2.542e+11Hz -0.0272045 -0.0107519
+ 2.543e+11Hz -0.0271614 -0.0106922
+ 2.544e+11Hz -0.0271181 -0.0106335
+ 2.545e+11Hz -0.0270746 -0.010576
+ 2.546e+11Hz -0.0270309 -0.0105197
+ 2.547e+11Hz -0.0269872 -0.0104644
+ 2.548e+11Hz -0.0269433 -0.0104103
+ 2.549e+11Hz -0.0268993 -0.0103573
+ 2.55e+11Hz -0.0268554 -0.0103054
+ 2.551e+11Hz -0.0268113 -0.0102546
+ 2.552e+11Hz -0.0267673 -0.0102049
+ 2.553e+11Hz -0.0267234 -0.0101562
+ 2.554e+11Hz -0.0266794 -0.0101086
+ 2.555e+11Hz -0.0266356 -0.0100621
+ 2.556e+11Hz -0.0265918 -0.0100166
+ 2.557e+11Hz -0.0265482 -0.00997211
+ 2.558e+11Hz -0.0265047 -0.00992863
+ 2.559e+11Hz -0.0264614 -0.00988615
+ 2.56e+11Hz -0.0264183 -0.00984465
+ 2.561e+11Hz -0.0263753 -0.00980412
+ 2.562e+11Hz -0.0263326 -0.00976454
+ 2.563e+11Hz -0.0262902 -0.0097259
+ 2.564e+11Hz -0.026248 -0.00968817
+ 2.565e+11Hz -0.0262061 -0.00965134
+ 2.566e+11Hz -0.0261645 -0.0096154
+ 2.567e+11Hz -0.0261232 -0.00958033
+ 2.568e+11Hz -0.0260822 -0.00954611
+ 2.569e+11Hz -0.0260416 -0.00951272
+ 2.57e+11Hz -0.0260014 -0.00948014
+ 2.571e+11Hz -0.0259616 -0.00944835
+ 2.572e+11Hz -0.0259221 -0.00941734
+ 2.573e+11Hz -0.025883 -0.00938708
+ 2.574e+11Hz -0.0258444 -0.00935756
+ 2.575e+11Hz -0.0258062 -0.00932876
+ 2.576e+11Hz -0.0257684 -0.00930065
+ 2.577e+11Hz -0.0257311 -0.00927321
+ 2.578e+11Hz -0.0256943 -0.00924643
+ 2.579e+11Hz -0.0256579 -0.00922029
+ 2.58e+11Hz -0.025622 -0.00919476
+ 2.581e+11Hz -0.0255866 -0.00916983
+ 2.582e+11Hz -0.0255516 -0.00914547
+ 2.583e+11Hz -0.0255172 -0.00912166
+ 2.584e+11Hz -0.0254833 -0.00909838
+ 2.585e+11Hz -0.0254499 -0.00907562
+ 2.586e+11Hz -0.025417 -0.00905334
+ 2.587e+11Hz -0.0253847 -0.00903154
+ 2.588e+11Hz -0.0253528 -0.00901018
+ 2.589e+11Hz -0.0253215 -0.00898926
+ 2.59e+11Hz -0.0252907 -0.00896874
+ 2.591e+11Hz -0.0252604 -0.00894862
+ 2.592e+11Hz -0.0252307 -0.00892886
+ 2.593e+11Hz -0.0252015 -0.00890945
+ 2.594e+11Hz -0.0251728 -0.00889037
+ 2.595e+11Hz -0.0251447 -0.0088716
+ 2.596e+11Hz -0.025117 -0.00885313
+ 2.597e+11Hz -0.0250899 -0.00883492
+ 2.598e+11Hz -0.0250633 -0.00881697
+ 2.599e+11Hz -0.0250373 -0.00879926
+ 2.6e+11Hz -0.0250117 -0.00878176
+ 2.601e+11Hz -0.0249866 -0.00876446
+ 2.602e+11Hz -0.0249621 -0.00874734
+ 2.603e+11Hz -0.024938 -0.00873039
+ 2.604e+11Hz -0.0249144 -0.00871359
+ 2.605e+11Hz -0.0248914 -0.00869692
+ 2.606e+11Hz -0.0248687 -0.00868037
+ 2.607e+11Hz -0.0248466 -0.00866392
+ 2.608e+11Hz -0.0248249 -0.00864756
+ 2.609e+11Hz -0.0248037 -0.00863126
+ 2.61e+11Hz -0.0247829 -0.00861503
+ 2.611e+11Hz -0.0247625 -0.00859884
+ 2.612e+11Hz -0.0247426 -0.00858268
+ 2.613e+11Hz -0.0247231 -0.00856654
+ 2.614e+11Hz -0.024704 -0.0085504
+ 2.615e+11Hz -0.0246852 -0.00853426
+ 2.616e+11Hz -0.0246669 -0.0085181
+ 2.617e+11Hz -0.0246489 -0.00850191
+ 2.618e+11Hz -0.0246313 -0.00848569
+ 2.619e+11Hz -0.0246141 -0.00846941
+ 2.62e+11Hz -0.0245971 -0.00845308
+ 2.621e+11Hz -0.0245805 -0.00843669
+ 2.622e+11Hz -0.0245642 -0.00842022
+ 2.623e+11Hz -0.0245483 -0.00840367
+ 2.624e+11Hz -0.0245326 -0.00838703
+ 2.625e+11Hz -0.0245171 -0.0083703
+ 2.626e+11Hz -0.024502 -0.00835347
+ 2.627e+11Hz -0.0244871 -0.00833653
+ 2.628e+11Hz -0.0244724 -0.00831948
+ 2.629e+11Hz -0.024458 -0.00830231
+ 2.63e+11Hz -0.0244437 -0.00828503
+ 2.631e+11Hz -0.0244297 -0.00826762
+ 2.632e+11Hz -0.0244159 -0.00825009
+ 2.633e+11Hz -0.0244022 -0.00823243
+ 2.634e+11Hz -0.0243887 -0.00821465
+ 2.635e+11Hz -0.0243753 -0.00819673
+ 2.636e+11Hz -0.0243621 -0.00817869
+ 2.637e+11Hz -0.024349 -0.00816051
+ 2.638e+11Hz -0.024336 -0.00814221
+ 2.639e+11Hz -0.0243231 -0.00812377
+ 2.64e+11Hz -0.0243104 -0.00810521
+ 2.641e+11Hz -0.0242976 -0.00808653
+ 2.642e+11Hz -0.024285 -0.00806772
+ 2.643e+11Hz -0.0242724 -0.00804879
+ 2.644e+11Hz -0.0242598 -0.00802974
+ 2.645e+11Hz -0.0242473 -0.00801059
+ 2.646e+11Hz -0.0242348 -0.00799132
+ 2.647e+11Hz -0.0242223 -0.00797195
+ 2.648e+11Hz -0.0242099 -0.00795248
+ 2.649e+11Hz -0.0241974 -0.00793292
+ 2.65e+11Hz -0.0241849 -0.00791326
+ 2.651e+11Hz -0.0241723 -0.00789353
+ 2.652e+11Hz -0.0241598 -0.00787372
+ 2.653e+11Hz -0.0241472 -0.00785385
+ 2.654e+11Hz -0.0241345 -0.00783391
+ 2.655e+11Hz -0.0241218 -0.00781392
+ 2.656e+11Hz -0.024109 -0.00779389
+ 2.657e+11Hz -0.0240962 -0.00777381
+ 2.658e+11Hz -0.0240833 -0.00775371
+ 2.659e+11Hz -0.0240703 -0.00773359
+ 2.66e+11Hz -0.0240572 -0.00771345
+ 2.661e+11Hz -0.024044 -0.00769331
+ 2.662e+11Hz -0.0240307 -0.00767318
+ 2.663e+11Hz -0.0240174 -0.00765307
+ 2.664e+11Hz -0.0240039 -0.00763298
+ 2.665e+11Hz -0.0239903 -0.00761293
+ 2.666e+11Hz -0.0239766 -0.00759292
+ 2.667e+11Hz -0.0239628 -0.00757297
+ 2.668e+11Hz -0.0239489 -0.00755308
+ 2.669e+11Hz -0.0239349 -0.00753327
+ 2.67e+11Hz -0.0239207 -0.00751354
+ 2.671e+11Hz -0.0239065 -0.00749391
+ 2.672e+11Hz -0.0238921 -0.00747438
+ 2.673e+11Hz -0.0238776 -0.00745497
+ 2.674e+11Hz -0.023863 -0.00743569
+ 2.675e+11Hz -0.0238483 -0.00741655
+ 2.676e+11Hz -0.0238335 -0.00739755
+ 2.677e+11Hz -0.0238186 -0.00737871
+ 2.678e+11Hz -0.0238036 -0.00736004
+ 2.679e+11Hz -0.0237885 -0.00734154
+ 2.68e+11Hz -0.0237733 -0.00732323
+ 2.681e+11Hz -0.023758 -0.00730512
+ 2.682e+11Hz -0.0237426 -0.00728721
+ 2.683e+11Hz -0.0237272 -0.00726952
+ 2.684e+11Hz -0.0237116 -0.00725205
+ 2.685e+11Hz -0.0236961 -0.00723481
+ 2.686e+11Hz -0.0236804 -0.00721782
+ 2.687e+11Hz -0.0236647 -0.00720108
+ 2.688e+11Hz -0.023649 -0.00718459
+ 2.689e+11Hz -0.0236332 -0.00716837
+ 2.69e+11Hz -0.0236174 -0.00715243
+ 2.691e+11Hz -0.0236016 -0.00713676
+ 2.692e+11Hz -0.0235858 -0.00712139
+ 2.693e+11Hz -0.02357 -0.00710631
+ 2.694e+11Hz -0.0235542 -0.00709153
+ 2.695e+11Hz -0.0235384 -0.00707705
+ 2.696e+11Hz -0.0235227 -0.00706289
+ 2.697e+11Hz -0.023507 -0.00704905
+ 2.698e+11Hz -0.0234913 -0.00703552
+ 2.699e+11Hz -0.0234758 -0.00702233
+ 2.7e+11Hz -0.0234603 -0.00700946
+ 2.701e+11Hz -0.0234449 -0.00699693
+ 2.702e+11Hz -0.0234296 -0.00698474
+ 2.703e+11Hz -0.0234144 -0.00697288
+ 2.704e+11Hz -0.0233994 -0.00696137
+ 2.705e+11Hz -0.0233845 -0.0069502
+ 2.706e+11Hz -0.0233698 -0.00693938
+ 2.707e+11Hz -0.0233552 -0.0069289
+ 2.708e+11Hz -0.0233408 -0.00691877
+ 2.709e+11Hz -0.0233267 -0.00690898
+ 2.71e+11Hz -0.0233127 -0.00689953
+ 2.711e+11Hz -0.023299 -0.00689043
+ 2.712e+11Hz -0.0232855 -0.00688167
+ 2.713e+11Hz -0.0232723 -0.00687325
+ 2.714e+11Hz -0.0232593 -0.00686517
+ 2.715e+11Hz -0.0232466 -0.00685742
+ 2.716e+11Hz -0.0232342 -0.00684999
+ 2.717e+11Hz -0.0232222 -0.00684289
+ 2.718e+11Hz -0.0232104 -0.00683611
+ 2.719e+11Hz -0.0231991 -0.00682965
+ 2.72e+11Hz -0.023188 -0.00682349
+ 2.721e+11Hz -0.0231774 -0.00681763
+ 2.722e+11Hz -0.0231671 -0.00681207
+ 2.723e+11Hz -0.0231572 -0.0068068
+ 2.724e+11Hz -0.0231477 -0.0068018
+ 2.725e+11Hz -0.0231387 -0.00679707
+ 2.726e+11Hz -0.0231301 -0.0067926
+ 2.727e+11Hz -0.023122 -0.00678839
+ 2.728e+11Hz -0.0231143 -0.00678441
+ 2.729e+11Hz -0.0231071 -0.00678066
+ 2.73e+11Hz -0.0231004 -0.00677714
+ 2.731e+11Hz -0.0230942 -0.00677381
+ 2.732e+11Hz -0.0230885 -0.00677069
+ 2.733e+11Hz -0.0230834 -0.00676774
+ 2.734e+11Hz -0.0230788 -0.00676496
+ 2.735e+11Hz -0.0230747 -0.00676234
+ 2.736e+11Hz -0.0230712 -0.00675986
+ 2.737e+11Hz -0.0230683 -0.00675751
+ 2.738e+11Hz -0.0230659 -0.00675526
+ 2.739e+11Hz -0.0230642 -0.00675311
+ 2.74e+11Hz -0.0230631 -0.00675104
+ 2.741e+11Hz -0.0230625 -0.00674904
+ 2.742e+11Hz -0.0230626 -0.00674708
+ 2.743e+11Hz -0.0230634 -0.00674515
+ 2.744e+11Hz -0.0230647 -0.00674324
+ 2.745e+11Hz -0.0230667 -0.00674131
+ 2.746e+11Hz -0.0230694 -0.00673937
+ 2.747e+11Hz -0.0230727 -0.00673738
+ 2.748e+11Hz -0.0230767 -0.00673533
+ 2.749e+11Hz -0.0230813 -0.00673321
+ 2.75e+11Hz -0.0230867 -0.00673098
+ 2.751e+11Hz -0.0230927 -0.00672863
+ 2.752e+11Hz -0.0230994 -0.00672615
+ 2.753e+11Hz -0.0231067 -0.00672351
+ 2.754e+11Hz -0.0231148 -0.00672069
+ 2.755e+11Hz -0.0231236 -0.00671766
+ 2.756e+11Hz -0.023133 -0.00671442
+ 2.757e+11Hz -0.0231432 -0.00671094
+ 2.758e+11Hz -0.023154 -0.00670719
+ 2.759e+11Hz -0.0231655 -0.00670316
+ 2.76e+11Hz -0.0231778 -0.00669883
+ 2.761e+11Hz -0.0231907 -0.00669416
+ 2.762e+11Hz -0.0232043 -0.00668915
+ 2.763e+11Hz -0.0232186 -0.00668377
+ 2.764e+11Hz -0.0232336 -0.006678
+ 2.765e+11Hz -0.0232492 -0.00667182
+ 2.766e+11Hz -0.0232656 -0.0066652
+ 2.767e+11Hz -0.0232826 -0.00665812
+ 2.768e+11Hz -0.0233003 -0.00665056
+ 2.769e+11Hz -0.0233186 -0.0066425
+ 2.77e+11Hz -0.0233376 -0.00663392
+ 2.771e+11Hz -0.0233572 -0.0066248
+ 2.772e+11Hz -0.0233775 -0.00661511
+ 2.773e+11Hz -0.0233984 -0.00660483
+ 2.774e+11Hz -0.0234199 -0.00659395
+ 2.775e+11Hz -0.0234421 -0.00658244
+ 2.776e+11Hz -0.0234648 -0.00657027
+ 2.777e+11Hz -0.0234881 -0.00655743
+ 2.778e+11Hz -0.023512 -0.00654391
+ 2.779e+11Hz -0.0235365 -0.00652966
+ 2.78e+11Hz -0.0235615 -0.00651469
+ 2.781e+11Hz -0.0235871 -0.00649896
+ 2.782e+11Hz -0.0236132 -0.00648246
+ 2.783e+11Hz -0.0236398 -0.00646517
+ 2.784e+11Hz -0.0236669 -0.00644706
+ 2.785e+11Hz -0.0236944 -0.00642812
+ 2.786e+11Hz -0.0237225 -0.00640834
+ 2.787e+11Hz -0.0237509 -0.00638769
+ 2.788e+11Hz -0.0237799 -0.00636615
+ 2.789e+11Hz -0.0238092 -0.0063437
+ 2.79e+11Hz -0.0238389 -0.00632034
+ 2.791e+11Hz -0.023869 -0.00629604
+ 2.792e+11Hz -0.0238994 -0.00627079
+ 2.793e+11Hz -0.0239302 -0.00624457
+ 2.794e+11Hz -0.0239613 -0.00621736
+ 2.795e+11Hz -0.0239926 -0.00618915
+ 2.796e+11Hz -0.0240243 -0.00615992
+ 2.797e+11Hz -0.0240562 -0.00612967
+ 2.798e+11Hz -0.0240883 -0.00609837
+ 2.799e+11Hz -0.0241206 -0.00606602
+ 2.8e+11Hz -0.0241531 -0.0060326
+ 2.801e+11Hz -0.0241858 -0.0059981
+ 2.802e+11Hz -0.0242186 -0.0059625
+ 2.803e+11Hz -0.0242515 -0.0059258
+ 2.804e+11Hz -0.0242845 -0.00588799
+ 2.805e+11Hz -0.0243176 -0.00584905
+ 2.806e+11Hz -0.0243507 -0.00580898
+ 2.807e+11Hz -0.0243838 -0.00576776
+ 2.808e+11Hz -0.0244169 -0.00572539
+ 2.809e+11Hz -0.0244499 -0.00568187
+ 2.81e+11Hz -0.0244829 -0.00563718
+ 2.811e+11Hz -0.0245158 -0.00559131
+ 2.812e+11Hz -0.0245486 -0.00554427
+ 2.813e+11Hz -0.0245812 -0.00549604
+ 2.814e+11Hz -0.0246136 -0.00544663
+ 2.815e+11Hz -0.0246459 -0.00539602
+ 2.816e+11Hz -0.0246779 -0.00534422
+ 2.817e+11Hz -0.0247096 -0.00529122
+ 2.818e+11Hz -0.024741 -0.00523701
+ 2.819e+11Hz -0.0247722 -0.00518161
+ 2.82e+11Hz -0.024803 -0.005125
+ 2.821e+11Hz -0.0248334 -0.00506719
+ 2.822e+11Hz -0.0248634 -0.00500818
+ 2.823e+11Hz -0.024893 -0.00494797
+ 2.824e+11Hz -0.0249221 -0.00488655
+ 2.825e+11Hz -0.0249508 -0.00482394
+ 2.826e+11Hz -0.0249789 -0.00476014
+ 2.827e+11Hz -0.0250065 -0.00469515
+ 2.828e+11Hz -0.0250335 -0.00462897
+ 2.829e+11Hz -0.0250599 -0.00456161
+ 2.83e+11Hz -0.0250857 -0.00449308
+ 2.831e+11Hz -0.0251108 -0.00442338
+ 2.832e+11Hz -0.0251352 -0.00435252
+ 2.833e+11Hz -0.025159 -0.0042805
+ 2.834e+11Hz -0.0251819 -0.00420735
+ 2.835e+11Hz -0.0252041 -0.00413305
+ 2.836e+11Hz -0.0252255 -0.00405764
+ 2.837e+11Hz -0.0252461 -0.0039811
+ 2.838e+11Hz -0.0252658 -0.00390347
+ 2.839e+11Hz -0.0252847 -0.00382474
+ 2.84e+11Hz -0.0253026 -0.00374494
+ 2.841e+11Hz -0.0253196 -0.00366406
+ 2.842e+11Hz -0.0253356 -0.00358214
+ 2.843e+11Hz -0.0253506 -0.00349918
+ 2.844e+11Hz -0.0253646 -0.00341519
+ 2.845e+11Hz -0.0253776 -0.0033302
+ 2.846e+11Hz -0.0253895 -0.00324421
+ 2.847e+11Hz -0.0254003 -0.00315725
+ 2.848e+11Hz -0.02541 -0.00306933
+ 2.849e+11Hz -0.0254185 -0.00298048
+ 2.85e+11Hz -0.0254259 -0.0028907
+ 2.851e+11Hz -0.0254321 -0.00280002
+ 2.852e+11Hz -0.025437 -0.00270846
+ 2.853e+11Hz -0.0254408 -0.00261604
+ 2.854e+11Hz -0.0254432 -0.00252278
+ 2.855e+11Hz -0.0254444 -0.0024287
+ 2.856e+11Hz -0.0254442 -0.00233382
+ 2.857e+11Hz -0.0254428 -0.00223816
+ 2.858e+11Hz -0.0254399 -0.00214176
+ 2.859e+11Hz -0.0254357 -0.00204462
+ 2.86e+11Hz -0.0254302 -0.00194678
+ 2.861e+11Hz -0.0254232 -0.00184826
+ 2.862e+11Hz -0.0254147 -0.00174909
+ 2.863e+11Hz -0.0254048 -0.00164928
+ 2.864e+11Hz -0.0253935 -0.00154887
+ 2.865e+11Hz -0.0253806 -0.00144788
+ 2.866e+11Hz -0.0253663 -0.00134634
+ 2.867e+11Hz -0.0253504 -0.00124428
+ 2.868e+11Hz -0.025333 -0.00114172
+ 2.869e+11Hz -0.025314 -0.00103869
+ 2.87e+11Hz -0.0252935 -0.000935225
+ 2.871e+11Hz -0.0252714 -0.000831344
+ 2.872e+11Hz -0.0252477 -0.00072708
+ 2.873e+11Hz -0.0252224 -0.000622463
+ 2.874e+11Hz -0.0251954 -0.000517523
+ 2.875e+11Hz -0.0251668 -0.000412288
+ 2.876e+11Hz -0.0251366 -0.00030679
+ 2.877e+11Hz -0.0251047 -0.00020106
+ 2.878e+11Hz -0.0250711 -9.51269e-05
+ 2.879e+11Hz -0.0250359 1.09765e-05
+ 2.88e+11Hz -0.024999 0.000117219
+ 2.881e+11Hz -0.0249603 0.00022357
+ 2.882e+11Hz -0.02492 0.000329996
+ 2.883e+11Hz -0.024878 0.000436466
+ 2.884e+11Hz -0.0248342 0.000542948
+ 2.885e+11Hz -0.0247887 0.000649409
+ 2.886e+11Hz -0.0247415 0.000755816
+ 2.887e+11Hz -0.0246926 0.000862137
+ 2.888e+11Hz -0.0246419 0.000968339
+ 2.889e+11Hz -0.0245895 0.00107439
+ 2.89e+11Hz -0.0245353 0.00118025
+ 2.891e+11Hz -0.0244794 0.0012859
+ 2.892e+11Hz -0.0244217 0.00139129
+ 2.893e+11Hz -0.0243623 0.0014964
+ 2.894e+11Hz -0.0243012 0.00160119
+ 2.895e+11Hz -0.0242383 0.00170563
+ 2.896e+11Hz -0.0241736 0.00180968
+ 2.897e+11Hz -0.0241073 0.00191331
+ 2.898e+11Hz -0.0240392 0.00201649
+ 2.899e+11Hz -0.0239693 0.00211918
+ 2.9e+11Hz -0.0238977 0.00222136
+ 2.901e+11Hz -0.0238244 0.00232298
+ 2.902e+11Hz -0.0237494 0.00242402
+ 2.903e+11Hz -0.0236727 0.00252443
+ 2.904e+11Hz -0.0235943 0.0026242
+ 2.905e+11Hz -0.0235141 0.00272327
+ 2.906e+11Hz -0.0234323 0.00282163
+ 2.907e+11Hz -0.0233488 0.00291924
+ 2.908e+11Hz -0.0232636 0.00301607
+ 2.909e+11Hz -0.0231768 0.00311207
+ 2.91e+11Hz -0.0230883 0.00320723
+ 2.911e+11Hz -0.0229982 0.00330151
+ 2.912e+11Hz -0.0229065 0.00339488
+ 2.913e+11Hz -0.0228132 0.00348731
+ 2.914e+11Hz -0.0227182 0.00357876
+ 2.915e+11Hz -0.0226217 0.0036692
+ 2.916e+11Hz -0.0225237 0.00375861
+ 2.917e+11Hz -0.022424 0.00384694
+ 2.918e+11Hz -0.0223229 0.00393419
+ 2.919e+11Hz -0.0222202 0.0040203
+ 2.92e+11Hz -0.022116 0.00410526
+ 2.921e+11Hz -0.0220104 0.00418903
+ 2.922e+11Hz -0.0219033 0.00427158
+ 2.923e+11Hz -0.0217947 0.00435289
+ 2.924e+11Hz -0.0216847 0.00443293
+ 2.925e+11Hz -0.0215734 0.00451167
+ 2.926e+11Hz -0.0214606 0.00458908
+ 2.927e+11Hz -0.0213465 0.00466514
+ 2.928e+11Hz -0.0212311 0.00473982
+ 2.929e+11Hz -0.0211143 0.00481309
+ 2.93e+11Hz -0.0209963 0.00488493
+ 2.931e+11Hz -0.020877 0.00495531
+ 2.932e+11Hz -0.0207564 0.00502421
+ 2.933e+11Hz -0.0206347 0.0050916
+ 2.934e+11Hz -0.0205117 0.00515746
+ 2.935e+11Hz -0.0203876 0.00522177
+ 2.936e+11Hz -0.0202624 0.0052845
+ 2.937e+11Hz -0.0201361 0.00534563
+ 2.938e+11Hz -0.0200086 0.00540515
+ 2.939e+11Hz -0.0198802 0.00546302
+ 2.94e+11Hz -0.0197507 0.00551923
+ 2.941e+11Hz -0.0196202 0.00557376
+ 2.942e+11Hz -0.0194887 0.00562659
+ 2.943e+11Hz -0.0193563 0.0056777
+ 2.944e+11Hz -0.019223 0.00572707
+ 2.945e+11Hz -0.0190888 0.00577469
+ 2.946e+11Hz -0.0189538 0.00582053
+ 2.947e+11Hz -0.018818 0.00586458
+ 2.948e+11Hz -0.0186813 0.00590683
+ 2.949e+11Hz -0.018544 0.00594726
+ 2.95e+11Hz -0.0184059 0.00598586
+ 2.951e+11Hz -0.0182671 0.0060226
+ 2.952e+11Hz -0.0181277 0.00605749
+ 2.953e+11Hz -0.0179877 0.0060905
+ 2.954e+11Hz -0.017847 0.00612163
+ 2.955e+11Hz -0.0177058 0.00615086
+ 2.956e+11Hz -0.0175641 0.00617818
+ 2.957e+11Hz -0.017422 0.00620358
+ 2.958e+11Hz -0.0172793 0.00622706
+ 2.959e+11Hz -0.0171363 0.0062486
+ 2.96e+11Hz -0.0169929 0.0062682
+ 2.961e+11Hz -0.0168491 0.00628586
+ 2.962e+11Hz -0.016705 0.00630155
+ 2.963e+11Hz -0.0165606 0.00631529
+ 2.964e+11Hz -0.016416 0.00632705
+ 2.965e+11Hz -0.0162712 0.00633685
+ 2.966e+11Hz -0.0161262 0.00634468
+ 2.967e+11Hz -0.0159811 0.00635052
+ 2.968e+11Hz -0.0158359 0.00635439
+ 2.969e+11Hz -0.0156906 0.00635628
+ 2.97e+11Hz -0.0155453 0.00635619
+ 2.971e+11Hz -0.0154 0.00635411
+ 2.972e+11Hz -0.0152547 0.00635006
+ 2.973e+11Hz -0.0151095 0.00634403
+ 2.974e+11Hz -0.0149645 0.00633603
+ 2.975e+11Hz -0.0148195 0.00632605
+ 2.976e+11Hz -0.0146748 0.0063141
+ 2.977e+11Hz -0.0145303 0.00630019
+ 2.978e+11Hz -0.014386 0.00628432
+ 2.979e+11Hz -0.014242 0.0062665
+ 2.98e+11Hz -0.0140984 0.00624673
+ 2.981e+11Hz -0.0139551 0.00622503
+ 2.982e+11Hz -0.0138121 0.00620139
+ 2.983e+11Hz -0.0136697 0.00617583
+ 2.984e+11Hz -0.0135276 0.00614836
+ 2.985e+11Hz -0.0133861 0.00611898
+ 2.986e+11Hz -0.0132451 0.00608772
+ 2.987e+11Hz -0.0131047 0.00605458
+ 2.988e+11Hz -0.0129648 0.00601957
+ 2.989e+11Hz -0.0128256 0.0059827
+ 2.99e+11Hz -0.0126871 0.00594399
+ 2.991e+11Hz -0.0125492 0.00590346
+ 2.992e+11Hz -0.0124121 0.00586112
+ 2.993e+11Hz -0.0122757 0.00581698
+ 2.994e+11Hz -0.0121401 0.00577107
+ 2.995e+11Hz -0.0120054 0.00572339
+ 2.996e+11Hz -0.0118714 0.00567396
+ 2.997e+11Hz -0.0117384 0.00562281
+ 2.998e+11Hz -0.0116063 0.00556996
+ 2.999e+11Hz -0.0114751 0.00551541
+ 3e+11Hz -0.0113448 0.0054592
+ ]

.ENDS
.SUBCKT Sub_SPfile_X5 1 2 3
R1N 1 10 -50
R1P 10 11 100
R2N 2 20 -50
R2P 20 21 100

A11 %vd(10 3) %vd(11, 12) xfer1
.model xfer1 xfer R_I=true table=[
+ 0Hz 0.00291081 0
+ 1e+08Hz 0.00291087 7.06655e-05
+ 2e+08Hz 0.00291105 0.000141329
+ 3e+08Hz 0.00291135 0.000211989
+ 4e+08Hz 0.00291177 0.000282643
+ 5e+08Hz 0.00291231 0.00035329
+ 6e+08Hz 0.00291298 0.000423928
+ 7e+08Hz 0.00291376 0.000494555
+ 8e+08Hz 0.00291466 0.000565169
+ 9e+08Hz 0.00291568 0.000635768
+ 1e+09Hz 0.00291682 0.00070635
+ 1.1e+09Hz 0.00291808 0.000776915
+ 1.2e+09Hz 0.00291946 0.000847459
+ 1.3e+09Hz 0.00292095 0.000917981
+ 1.4e+09Hz 0.00292256 0.00098848
+ 1.5e+09Hz 0.00292429 0.00105895
+ 1.6e+09Hz 0.00292613 0.0011294
+ 1.7e+09Hz 0.00292809 0.00119982
+ 1.8e+09Hz 0.00293017 0.0012702
+ 1.9e+09Hz 0.00293236 0.00134056
+ 2e+09Hz 0.00293466 0.00141088
+ 2.1e+09Hz 0.00293708 0.00148116
+ 2.2e+09Hz 0.0029396 0.00155141
+ 2.3e+09Hz 0.00294224 0.00162162
+ 2.4e+09Hz 0.00294499 0.00169179
+ 2.5e+09Hz 0.00294785 0.00176191
+ 2.6e+09Hz 0.00295082 0.001832
+ 2.7e+09Hz 0.00295389 0.00190203
+ 2.8e+09Hz 0.00295707 0.00197202
+ 2.9e+09Hz 0.00296036 0.00204197
+ 3e+09Hz 0.00296375 0.00211186
+ 3.1e+09Hz 0.00296724 0.0021817
+ 3.2e+09Hz 0.00297084 0.00225149
+ 3.3e+09Hz 0.00297454 0.00232123
+ 3.4e+09Hz 0.00297834 0.00239091
+ 3.5e+09Hz 0.00298223 0.00246053
+ 3.6e+09Hz 0.00298623 0.0025301
+ 3.7e+09Hz 0.00299032 0.00259961
+ 3.8e+09Hz 0.00299451 0.00266906
+ 3.9e+09Hz 0.00299879 0.00273844
+ 4e+09Hz 0.00300316 0.00280777
+ 4.1e+09Hz 0.00300763 0.00287703
+ 4.2e+09Hz 0.00301219 0.00294622
+ 4.3e+09Hz 0.00301683 0.00301535
+ 4.4e+09Hz 0.00302156 0.00308442
+ 4.5e+09Hz 0.00302638 0.00315341
+ 4.6e+09Hz 0.00303128 0.00322234
+ 4.7e+09Hz 0.00303627 0.0032912
+ 4.8e+09Hz 0.00304134 0.00335999
+ 4.9e+09Hz 0.00304648 0.0034287
+ 5e+09Hz 0.00305171 0.00349734
+ 5.1e+09Hz 0.00305702 0.00356592
+ 5.2e+09Hz 0.0030624 0.00363441
+ 5.3e+09Hz 0.00306785 0.00370283
+ 5.4e+09Hz 0.00307338 0.00377118
+ 5.5e+09Hz 0.00307898 0.00383945
+ 5.6e+09Hz 0.00308465 0.00390765
+ 5.7e+09Hz 0.00309039 0.00397577
+ 5.8e+09Hz 0.00309619 0.00404381
+ 5.9e+09Hz 0.00310207 0.00411177
+ 6e+09Hz 0.003108 0.00417966
+ 6.1e+09Hz 0.003114 0.00424746
+ 6.2e+09Hz 0.00312006 0.00431519
+ 6.3e+09Hz 0.00312617 0.00438284
+ 6.4e+09Hz 0.00313235 0.00445041
+ 6.5e+09Hz 0.00313858 0.00451789
+ 6.6e+09Hz 0.00314487 0.0045853
+ 6.7e+09Hz 0.00315121 0.00465263
+ 6.8e+09Hz 0.0031576 0.00471987
+ 6.9e+09Hz 0.00316404 0.00478704
+ 7e+09Hz 0.00317053 0.00485412
+ 7.1e+09Hz 0.00317707 0.00492112
+ 7.2e+09Hz 0.00318365 0.00498804
+ 7.3e+09Hz 0.00319028 0.00505489
+ 7.4e+09Hz 0.00319695 0.00512164
+ 7.5e+09Hz 0.00320366 0.00518832
+ 7.6e+09Hz 0.00321042 0.00525492
+ 7.7e+09Hz 0.00321721 0.00532144
+ 7.8e+09Hz 0.00322403 0.00538787
+ 7.9e+09Hz 0.0032309 0.00545423
+ 8e+09Hz 0.00323779 0.0055205
+ 8.1e+09Hz 0.00324472 0.0055867
+ 8.2e+09Hz 0.00325168 0.00565281
+ 8.3e+09Hz 0.00325867 0.00571885
+ 8.4e+09Hz 0.00326569 0.0057848
+ 8.5e+09Hz 0.00327274 0.00585068
+ 8.6e+09Hz 0.00327981 0.00591648
+ 8.7e+09Hz 0.00328691 0.0059822
+ 8.8e+09Hz 0.00329402 0.00604785
+ 8.9e+09Hz 0.00330117 0.00611341
+ 9e+09Hz 0.00330833 0.0061789
+ 9.1e+09Hz 0.00331551 0.00624432
+ 9.2e+09Hz 0.00332271 0.00630965
+ 9.3e+09Hz 0.00332993 0.00637492
+ 9.4e+09Hz 0.00333716 0.00644011
+ 9.5e+09Hz 0.00334441 0.00650522
+ 9.6e+09Hz 0.00335167 0.00657026
+ 9.7e+09Hz 0.00335894 0.00663523
+ 9.8e+09Hz 0.00336623 0.00670013
+ 9.9e+09Hz 0.00337352 0.00676496
+ 1e+10Hz 0.00338082 0.00682971
+ 1.01e+10Hz 0.00338814 0.0068944
+ 1.02e+10Hz 0.00339545 0.00695902
+ 1.03e+10Hz 0.00340278 0.00702356
+ 1.04e+10Hz 0.00341011 0.00708805
+ 1.05e+10Hz 0.00341744 0.00715246
+ 1.06e+10Hz 0.00342478 0.00721681
+ 1.07e+10Hz 0.00343212 0.00728109
+ 1.08e+10Hz 0.00343946 0.00734531
+ 1.09e+10Hz 0.0034468 0.00740947
+ 1.1e+10Hz 0.00345415 0.00747356
+ 1.11e+10Hz 0.00346149 0.00753759
+ 1.12e+10Hz 0.00346882 0.00760157
+ 1.13e+10Hz 0.00347616 0.00766548
+ 1.14e+10Hz 0.00348349 0.00772933
+ 1.15e+10Hz 0.00349082 0.00779312
+ 1.16e+10Hz 0.00349815 0.00785686
+ 1.17e+10Hz 0.00350547 0.00792054
+ 1.18e+10Hz 0.00351278 0.00798416
+ 1.19e+10Hz 0.00352009 0.00804773
+ 1.2e+10Hz 0.00352738 0.00811125
+ 1.21e+10Hz 0.00353468 0.00817472
+ 1.22e+10Hz 0.00354196 0.00823813
+ 1.23e+10Hz 0.00354923 0.00830149
+ 1.24e+10Hz 0.0035565 0.0083648
+ 1.25e+10Hz 0.00356375 0.00842807
+ 1.26e+10Hz 0.003571 0.00849129
+ 1.27e+10Hz 0.00357823 0.00855446
+ 1.28e+10Hz 0.00358545 0.00861758
+ 1.29e+10Hz 0.00359267 0.00868066
+ 1.3e+10Hz 0.00359987 0.00874369
+ 1.31e+10Hz 0.00360706 0.00880669
+ 1.32e+10Hz 0.00361423 0.00886964
+ 1.33e+10Hz 0.00362139 0.00893255
+ 1.34e+10Hz 0.00362854 0.00899542
+ 1.35e+10Hz 0.00363568 0.00905825
+ 1.36e+10Hz 0.00364281 0.00912104
+ 1.37e+10Hz 0.00364992 0.0091838
+ 1.38e+10Hz 0.00365701 0.00924652
+ 1.39e+10Hz 0.0036641 0.0093092
+ 1.4e+10Hz 0.00367116 0.00937185
+ 1.41e+10Hz 0.00367822 0.00943447
+ 1.42e+10Hz 0.00368526 0.00949705
+ 1.43e+10Hz 0.00369229 0.0095596
+ 1.44e+10Hz 0.0036993 0.00962213
+ 1.45e+10Hz 0.00370629 0.00968462
+ 1.46e+10Hz 0.00371328 0.00974708
+ 1.47e+10Hz 0.00372025 0.00980952
+ 1.48e+10Hz 0.0037272 0.00987193
+ 1.49e+10Hz 0.00373414 0.00993431
+ 1.5e+10Hz 0.00374107 0.00999667
+ 1.51e+10Hz 0.00374798 0.010059
+ 1.52e+10Hz 0.00375488 0.0101213
+ 1.53e+10Hz 0.00376176 0.0101836
+ 1.54e+10Hz 0.00376863 0.0102459
+ 1.55e+10Hz 0.00377549 0.0103081
+ 1.56e+10Hz 0.00378233 0.0103703
+ 1.57e+10Hz 0.00378916 0.0104326
+ 1.58e+10Hz 0.00379598 0.0104947
+ 1.59e+10Hz 0.00380278 0.0105569
+ 1.6e+10Hz 0.00380957 0.0106191
+ 1.61e+10Hz 0.00381635 0.0106812
+ 1.62e+10Hz 0.00382312 0.0107433
+ 1.63e+10Hz 0.00382987 0.0108054
+ 1.64e+10Hz 0.00383661 0.0108675
+ 1.65e+10Hz 0.00384334 0.0109296
+ 1.66e+10Hz 0.00385006 0.0109917
+ 1.67e+10Hz 0.00385677 0.0110537
+ 1.68e+10Hz 0.00386347 0.0111158
+ 1.69e+10Hz 0.00387016 0.0111778
+ 1.7e+10Hz 0.00387684 0.0112398
+ 1.71e+10Hz 0.00388351 0.0113018
+ 1.72e+10Hz 0.00389017 0.0113638
+ 1.73e+10Hz 0.00389682 0.0114258
+ 1.74e+10Hz 0.00390346 0.0114878
+ 1.75e+10Hz 0.00391009 0.0115498
+ 1.76e+10Hz 0.00391672 0.0116118
+ 1.77e+10Hz 0.00392334 0.0116737
+ 1.78e+10Hz 0.00392995 0.0117357
+ 1.79e+10Hz 0.00393656 0.0117977
+ 1.8e+10Hz 0.00394316 0.0118596
+ 1.81e+10Hz 0.00394976 0.0119216
+ 1.82e+10Hz 0.00395635 0.0119835
+ 1.83e+10Hz 0.00396293 0.0120454
+ 1.84e+10Hz 0.00396951 0.0121074
+ 1.85e+10Hz 0.00397609 0.0121693
+ 1.86e+10Hz 0.00398266 0.0122313
+ 1.87e+10Hz 0.00398924 0.0122932
+ 1.88e+10Hz 0.0039958 0.0123552
+ 1.89e+10Hz 0.00400237 0.0124171
+ 1.9e+10Hz 0.00400893 0.012479
+ 1.91e+10Hz 0.0040155 0.012541
+ 1.92e+10Hz 0.00402206 0.0126029
+ 1.93e+10Hz 0.00402862 0.0126648
+ 1.94e+10Hz 0.00403519 0.0127268
+ 1.95e+10Hz 0.00404175 0.0127887
+ 1.96e+10Hz 0.00404832 0.0128506
+ 1.97e+10Hz 0.00405488 0.0129126
+ 1.98e+10Hz 0.00406145 0.0129745
+ 1.99e+10Hz 0.00406802 0.0130365
+ 2e+10Hz 0.0040746 0.0130984
+ 2.01e+10Hz 0.00408118 0.0131604
+ 2.02e+10Hz 0.00408776 0.0132223
+ 2.03e+10Hz 0.00409435 0.0132843
+ 2.04e+10Hz 0.00410094 0.0133463
+ 2.05e+10Hz 0.00410753 0.0134082
+ 2.06e+10Hz 0.00411414 0.0134702
+ 2.07e+10Hz 0.00412075 0.0135322
+ 2.08e+10Hz 0.00412736 0.0135942
+ 2.09e+10Hz 0.00413398 0.0136561
+ 2.1e+10Hz 0.00414062 0.0137181
+ 2.11e+10Hz 0.00414725 0.0137801
+ 2.12e+10Hz 0.0041539 0.0138421
+ 2.13e+10Hz 0.00416056 0.0139041
+ 2.14e+10Hz 0.00416723 0.0139661
+ 2.15e+10Hz 0.0041739 0.0140281
+ 2.16e+10Hz 0.00418059 0.0140901
+ 2.17e+10Hz 0.00418728 0.0141522
+ 2.18e+10Hz 0.00419399 0.0142142
+ 2.19e+10Hz 0.00420071 0.0142762
+ 2.2e+10Hz 0.00420744 0.0143383
+ 2.21e+10Hz 0.00421419 0.0144003
+ 2.22e+10Hz 0.00422094 0.0144623
+ 2.23e+10Hz 0.00422771 0.0145244
+ 2.24e+10Hz 0.0042345 0.0145864
+ 2.25e+10Hz 0.00424129 0.0146485
+ 2.26e+10Hz 0.0042481 0.0147106
+ 2.27e+10Hz 0.00425493 0.0147726
+ 2.28e+10Hz 0.00426177 0.0148347
+ 2.29e+10Hz 0.00426863 0.0148968
+ 2.3e+10Hz 0.0042755 0.0149588
+ 2.31e+10Hz 0.00428238 0.0150209
+ 2.32e+10Hz 0.00428929 0.015083
+ 2.33e+10Hz 0.00429621 0.0151451
+ 2.34e+10Hz 0.00430315 0.0152072
+ 2.35e+10Hz 0.0043101 0.0152693
+ 2.36e+10Hz 0.00431707 0.0153314
+ 2.37e+10Hz 0.00432406 0.0153935
+ 2.38e+10Hz 0.00433107 0.0154556
+ 2.39e+10Hz 0.0043381 0.0155177
+ 2.4e+10Hz 0.00434514 0.0155798
+ 2.41e+10Hz 0.00435221 0.015642
+ 2.42e+10Hz 0.00435929 0.0157041
+ 2.43e+10Hz 0.0043664 0.0157662
+ 2.44e+10Hz 0.00437352 0.0158283
+ 2.45e+10Hz 0.00438066 0.0158905
+ 2.46e+10Hz 0.00438782 0.0159526
+ 2.47e+10Hz 0.00439501 0.0160147
+ 2.48e+10Hz 0.00440221 0.0160769
+ 2.49e+10Hz 0.00440944 0.016139
+ 2.5e+10Hz 0.00441668 0.0162011
+ 2.51e+10Hz 0.00442395 0.0162633
+ 2.52e+10Hz 0.00443124 0.0163254
+ 2.53e+10Hz 0.00443855 0.0163875
+ 2.54e+10Hz 0.00444588 0.0164497
+ 2.55e+10Hz 0.00445323 0.0165118
+ 2.56e+10Hz 0.00446061 0.016574
+ 2.57e+10Hz 0.004468 0.0166361
+ 2.58e+10Hz 0.00447542 0.0166982
+ 2.59e+10Hz 0.00448287 0.0167604
+ 2.6e+10Hz 0.00449033 0.0168225
+ 2.61e+10Hz 0.00449782 0.0168847
+ 2.62e+10Hz 0.00450533 0.0169468
+ 2.63e+10Hz 0.00451286 0.0170089
+ 2.64e+10Hz 0.00452042 0.0170711
+ 2.65e+10Hz 0.004528 0.0171332
+ 2.66e+10Hz 0.0045356 0.0171953
+ 2.67e+10Hz 0.00454323 0.0172574
+ 2.68e+10Hz 0.00455088 0.0173195
+ 2.69e+10Hz 0.00455855 0.0173817
+ 2.7e+10Hz 0.00456624 0.0174438
+ 2.71e+10Hz 0.00457396 0.0175059
+ 2.72e+10Hz 0.00458171 0.017568
+ 2.73e+10Hz 0.00458947 0.0176301
+ 2.74e+10Hz 0.00459726 0.0176922
+ 2.75e+10Hz 0.00460507 0.0177543
+ 2.76e+10Hz 0.00461291 0.0178164
+ 2.77e+10Hz 0.00462077 0.0178785
+ 2.78e+10Hz 0.00462865 0.0179406
+ 2.79e+10Hz 0.00463656 0.0180027
+ 2.8e+10Hz 0.00464449 0.0180648
+ 2.81e+10Hz 0.00465245 0.0181268
+ 2.82e+10Hz 0.00466043 0.0181889
+ 2.83e+10Hz 0.00466843 0.018251
+ 2.84e+10Hz 0.00467645 0.018313
+ 2.85e+10Hz 0.0046845 0.0183751
+ 2.86e+10Hz 0.00469257 0.0184371
+ 2.87e+10Hz 0.00470066 0.0184992
+ 2.88e+10Hz 0.00470878 0.0185612
+ 2.89e+10Hz 0.00471693 0.0186232
+ 2.9e+10Hz 0.00472509 0.0186852
+ 2.91e+10Hz 0.00473328 0.0187473
+ 2.92e+10Hz 0.00474149 0.0188093
+ 2.93e+10Hz 0.00474972 0.0188712
+ 2.94e+10Hz 0.00475798 0.0189332
+ 2.95e+10Hz 0.00476626 0.0189952
+ 2.96e+10Hz 0.00477456 0.0190572
+ 2.97e+10Hz 0.00478288 0.0191192
+ 2.98e+10Hz 0.00479123 0.0191811
+ 2.99e+10Hz 0.0047996 0.0192431
+ 3e+10Hz 0.00480799 0.019305
+ 3.01e+10Hz 0.0048164 0.019367
+ 3.02e+10Hz 0.00482484 0.0194289
+ 3.03e+10Hz 0.0048333 0.0194908
+ 3.04e+10Hz 0.00484178 0.0195527
+ 3.05e+10Hz 0.00485028 0.0196146
+ 3.06e+10Hz 0.0048588 0.0196765
+ 3.07e+10Hz 0.00486735 0.0197384
+ 3.08e+10Hz 0.00487591 0.0198003
+ 3.09e+10Hz 0.0048845 0.0198621
+ 3.1e+10Hz 0.00489311 0.019924
+ 3.11e+10Hz 0.00490174 0.0199858
+ 3.12e+10Hz 0.00491039 0.0200477
+ 3.13e+10Hz 0.00491906 0.0201095
+ 3.14e+10Hz 0.00492775 0.0201713
+ 3.15e+10Hz 0.00493646 0.0202331
+ 3.16e+10Hz 0.00494519 0.0202949
+ 3.17e+10Hz 0.00495395 0.0203567
+ 3.18e+10Hz 0.00496272 0.0204185
+ 3.19e+10Hz 0.00497151 0.0204802
+ 3.2e+10Hz 0.00498032 0.020542
+ 3.21e+10Hz 0.00498916 0.0206038
+ 3.22e+10Hz 0.00499801 0.0206655
+ 3.23e+10Hz 0.00500688 0.0207272
+ 3.24e+10Hz 0.00501577 0.0207889
+ 3.25e+10Hz 0.00502468 0.0208506
+ 3.26e+10Hz 0.00503361 0.0209123
+ 3.27e+10Hz 0.00504255 0.020974
+ 3.28e+10Hz 0.00505152 0.0210357
+ 3.29e+10Hz 0.0050605 0.0210974
+ 3.3e+10Hz 0.00506951 0.021159
+ 3.31e+10Hz 0.00507853 0.0212207
+ 3.32e+10Hz 0.00508756 0.0212823
+ 3.33e+10Hz 0.00509662 0.0213439
+ 3.34e+10Hz 0.0051057 0.0214055
+ 3.35e+10Hz 0.00511479 0.0214672
+ 3.36e+10Hz 0.0051239 0.0215287
+ 3.37e+10Hz 0.00513303 0.0215903
+ 3.38e+10Hz 0.00514217 0.0216519
+ 3.39e+10Hz 0.00515133 0.0217135
+ 3.4e+10Hz 0.00516051 0.021775
+ 3.41e+10Hz 0.00516971 0.0218366
+ 3.42e+10Hz 0.00517892 0.0218981
+ 3.43e+10Hz 0.00518815 0.0219596
+ 3.44e+10Hz 0.00519739 0.0220211
+ 3.45e+10Hz 0.00520666 0.0220827
+ 3.46e+10Hz 0.00521593 0.0221442
+ 3.47e+10Hz 0.00522523 0.0222056
+ 3.48e+10Hz 0.00523454 0.0222671
+ 3.49e+10Hz 0.00524387 0.0223286
+ 3.5e+10Hz 0.00525321 0.02239
+ 3.51e+10Hz 0.00526257 0.0224515
+ 3.52e+10Hz 0.00527194 0.0225129
+ 3.53e+10Hz 0.00528133 0.0225743
+ 3.54e+10Hz 0.00529073 0.0226358
+ 3.55e+10Hz 0.00530015 0.0226972
+ 3.56e+10Hz 0.00530959 0.0227586
+ 3.57e+10Hz 0.00531904 0.02282
+ 3.58e+10Hz 0.0053285 0.0228814
+ 3.59e+10Hz 0.00533798 0.0229427
+ 3.6e+10Hz 0.00534747 0.0230041
+ 3.61e+10Hz 0.00535698 0.0230654
+ 3.62e+10Hz 0.00536651 0.0231268
+ 3.63e+10Hz 0.00537605 0.0231881
+ 3.64e+10Hz 0.0053856 0.0232495
+ 3.65e+10Hz 0.00539517 0.0233108
+ 3.66e+10Hz 0.00540475 0.0233721
+ 3.67e+10Hz 0.00541434 0.0234334
+ 3.68e+10Hz 0.00542395 0.0234947
+ 3.69e+10Hz 0.00543358 0.023556
+ 3.7e+10Hz 0.00544321 0.0236173
+ 3.71e+10Hz 0.00545287 0.0236785
+ 3.72e+10Hz 0.00546253 0.0237398
+ 3.73e+10Hz 0.00547221 0.0238011
+ 3.74e+10Hz 0.0054819 0.0238623
+ 3.75e+10Hz 0.00549161 0.0239235
+ 3.76e+10Hz 0.00550133 0.0239848
+ 3.77e+10Hz 0.00551107 0.024046
+ 3.78e+10Hz 0.00552082 0.0241072
+ 3.79e+10Hz 0.00553058 0.0241684
+ 3.8e+10Hz 0.00554036 0.0242296
+ 3.81e+10Hz 0.00555014 0.0242908
+ 3.82e+10Hz 0.00555995 0.024352
+ 3.83e+10Hz 0.00556976 0.0244132
+ 3.84e+10Hz 0.00557959 0.0244744
+ 3.85e+10Hz 0.00558944 0.0245356
+ 3.86e+10Hz 0.00559929 0.0245968
+ 3.87e+10Hz 0.00560916 0.0246579
+ 3.88e+10Hz 0.00561905 0.0247191
+ 3.89e+10Hz 0.00562894 0.0247802
+ 3.9e+10Hz 0.00563885 0.0248414
+ 3.91e+10Hz 0.00564878 0.0249025
+ 3.92e+10Hz 0.00565871 0.0249636
+ 3.93e+10Hz 0.00566867 0.0250248
+ 3.94e+10Hz 0.00567863 0.0250859
+ 3.95e+10Hz 0.00568861 0.025147
+ 3.96e+10Hz 0.0056986 0.0252081
+ 3.97e+10Hz 0.0057086 0.0252692
+ 3.98e+10Hz 0.00571862 0.0253303
+ 3.99e+10Hz 0.00572865 0.0253914
+ 4e+10Hz 0.0057387 0.0254525
+ 4.01e+10Hz 0.00574876 0.0255136
+ 4.02e+10Hz 0.00575883 0.0255747
+ 4.03e+10Hz 0.00576892 0.0256358
+ 4.04e+10Hz 0.00577902 0.0256968
+ 4.05e+10Hz 0.00578913 0.0257579
+ 4.06e+10Hz 0.00579926 0.025819
+ 4.07e+10Hz 0.0058094 0.02588
+ 4.08e+10Hz 0.00581955 0.0259411
+ 4.09e+10Hz 0.00582972 0.0260021
+ 4.1e+10Hz 0.0058399 0.0260632
+ 4.11e+10Hz 0.0058501 0.0261242
+ 4.12e+10Hz 0.00586031 0.0261853
+ 4.13e+10Hz 0.00587054 0.0262463
+ 4.14e+10Hz 0.00588078 0.0263074
+ 4.15e+10Hz 0.00589103 0.0263684
+ 4.16e+10Hz 0.0059013 0.0264294
+ 4.17e+10Hz 0.00591158 0.0264904
+ 4.18e+10Hz 0.00592188 0.0265515
+ 4.19e+10Hz 0.00593219 0.0266125
+ 4.2e+10Hz 0.00594251 0.0266735
+ 4.21e+10Hz 0.00595285 0.0267345
+ 4.22e+10Hz 0.00596321 0.0267955
+ 4.23e+10Hz 0.00597357 0.0268565
+ 4.24e+10Hz 0.00598396 0.0269175
+ 4.25e+10Hz 0.00599436 0.0269786
+ 4.26e+10Hz 0.00600477 0.0270395
+ 4.27e+10Hz 0.0060152 0.0271005
+ 4.28e+10Hz 0.00602564 0.0271615
+ 4.29e+10Hz 0.0060361 0.0272225
+ 4.3e+10Hz 0.00604658 0.0272835
+ 4.31e+10Hz 0.00605707 0.0273445
+ 4.32e+10Hz 0.00606758 0.0274055
+ 4.33e+10Hz 0.0060781 0.0274665
+ 4.34e+10Hz 0.00608863 0.0275275
+ 4.35e+10Hz 0.00609919 0.0275884
+ 4.36e+10Hz 0.00610975 0.0276494
+ 4.37e+10Hz 0.00612034 0.0277104
+ 4.38e+10Hz 0.00613094 0.0277714
+ 4.39e+10Hz 0.00614155 0.0278323
+ 4.4e+10Hz 0.00615219 0.0278933
+ 4.41e+10Hz 0.00616284 0.0279543
+ 4.42e+10Hz 0.0061735 0.0280152
+ 4.43e+10Hz 0.00618418 0.0280762
+ 4.44e+10Hz 0.00619488 0.0281372
+ 4.45e+10Hz 0.0062056 0.0281981
+ 4.46e+10Hz 0.00621633 0.0282591
+ 4.47e+10Hz 0.00622708 0.02832
+ 4.48e+10Hz 0.00623784 0.028381
+ 4.49e+10Hz 0.00624862 0.028442
+ 4.5e+10Hz 0.00625942 0.0285029
+ 4.51e+10Hz 0.00627024 0.0285639
+ 4.52e+10Hz 0.00628107 0.0286248
+ 4.53e+10Hz 0.00629193 0.0286857
+ 4.54e+10Hz 0.00630279 0.0287467
+ 4.55e+10Hz 0.00631368 0.0288076
+ 4.56e+10Hz 0.00632458 0.0288686
+ 4.57e+10Hz 0.0063355 0.0289295
+ 4.58e+10Hz 0.00634645 0.0289905
+ 4.59e+10Hz 0.0063574 0.0290514
+ 4.6e+10Hz 0.00636838 0.0291123
+ 4.61e+10Hz 0.00637937 0.0291733
+ 4.62e+10Hz 0.00639038 0.0292342
+ 4.63e+10Hz 0.00640141 0.0292951
+ 4.64e+10Hz 0.00641246 0.029356
+ 4.65e+10Hz 0.00642353 0.029417
+ 4.66e+10Hz 0.00643461 0.0294779
+ 4.67e+10Hz 0.00644572 0.0295388
+ 4.68e+10Hz 0.00645684 0.0295997
+ 4.69e+10Hz 0.00646798 0.0296606
+ 4.7e+10Hz 0.00647914 0.0297215
+ 4.71e+10Hz 0.00649032 0.0297824
+ 4.72e+10Hz 0.00650152 0.0298434
+ 4.73e+10Hz 0.00651274 0.0299043
+ 4.74e+10Hz 0.00652397 0.0299652
+ 4.75e+10Hz 0.00653523 0.0300261
+ 4.76e+10Hz 0.00654651 0.030087
+ 4.77e+10Hz 0.0065578 0.0301479
+ 4.78e+10Hz 0.00656912 0.0302088
+ 4.79e+10Hz 0.00658045 0.0302696
+ 4.8e+10Hz 0.0065918 0.0303305
+ 4.81e+10Hz 0.00660318 0.0303914
+ 4.82e+10Hz 0.00661457 0.0304523
+ 4.83e+10Hz 0.00662598 0.0305132
+ 4.84e+10Hz 0.00663741 0.0305741
+ 4.85e+10Hz 0.00664887 0.030635
+ 4.86e+10Hz 0.00666034 0.0306958
+ 4.87e+10Hz 0.00667183 0.0307567
+ 4.88e+10Hz 0.00668335 0.0308176
+ 4.89e+10Hz 0.00669488 0.0308784
+ 4.9e+10Hz 0.00670643 0.0309393
+ 4.91e+10Hz 0.006718 0.0310001
+ 4.92e+10Hz 0.0067296 0.031061
+ 4.93e+10Hz 0.00674121 0.0311218
+ 4.94e+10Hz 0.00675285 0.0311827
+ 4.95e+10Hz 0.0067645 0.0312435
+ 4.96e+10Hz 0.00677618 0.0313044
+ 4.97e+10Hz 0.00678788 0.0313652
+ 4.98e+10Hz 0.0067996 0.031426
+ 4.99e+10Hz 0.00681133 0.0314869
+ 5e+10Hz 0.00682309 0.0315477
+ 5.01e+10Hz 0.00683487 0.0316085
+ 5.02e+10Hz 0.00684667 0.0316693
+ 5.03e+10Hz 0.00685849 0.0317301
+ 5.04e+10Hz 0.00687034 0.0317909
+ 5.05e+10Hz 0.0068822 0.0318518
+ 5.06e+10Hz 0.00689408 0.0319126
+ 5.07e+10Hz 0.00690599 0.0319733
+ 5.08e+10Hz 0.00691791 0.0320341
+ 5.09e+10Hz 0.00692986 0.0320949
+ 5.1e+10Hz 0.00694183 0.0321557
+ 5.11e+10Hz 0.00695382 0.0322165
+ 5.12e+10Hz 0.00696583 0.0322773
+ 5.13e+10Hz 0.00697786 0.032338
+ 5.14e+10Hz 0.00698991 0.0323988
+ 5.15e+10Hz 0.00700198 0.0324595
+ 5.16e+10Hz 0.00701408 0.0325203
+ 5.17e+10Hz 0.0070262 0.0325811
+ 5.18e+10Hz 0.00703833 0.0326418
+ 5.19e+10Hz 0.00705049 0.0327025
+ 5.2e+10Hz 0.00706267 0.0327633
+ 5.21e+10Hz 0.00707487 0.032824
+ 5.22e+10Hz 0.00708709 0.0328847
+ 5.23e+10Hz 0.00709934 0.0329454
+ 5.24e+10Hz 0.0071116 0.0330061
+ 5.25e+10Hz 0.00712388 0.0330668
+ 5.26e+10Hz 0.00713619 0.0331275
+ 5.27e+10Hz 0.00714852 0.0331882
+ 5.28e+10Hz 0.00716087 0.0332489
+ 5.29e+10Hz 0.00717324 0.0333096
+ 5.3e+10Hz 0.00718563 0.0333703
+ 5.31e+10Hz 0.00719804 0.0334309
+ 5.32e+10Hz 0.00721047 0.0334916
+ 5.33e+10Hz 0.00722292 0.0335522
+ 5.34e+10Hz 0.0072354 0.0336129
+ 5.35e+10Hz 0.0072479 0.0336735
+ 5.36e+10Hz 0.00726041 0.0337342
+ 5.37e+10Hz 0.00727295 0.0337948
+ 5.38e+10Hz 0.00728551 0.0338554
+ 5.39e+10Hz 0.00729809 0.033916
+ 5.4e+10Hz 0.00731069 0.0339766
+ 5.41e+10Hz 0.00732331 0.0340372
+ 5.42e+10Hz 0.00733596 0.0340978
+ 5.43e+10Hz 0.00734862 0.0341584
+ 5.44e+10Hz 0.00736131 0.034219
+ 5.45e+10Hz 0.00737401 0.0342796
+ 5.46e+10Hz 0.00738674 0.0343401
+ 5.47e+10Hz 0.00739948 0.0344007
+ 5.48e+10Hz 0.00741225 0.0344612
+ 5.49e+10Hz 0.00742504 0.0345218
+ 5.5e+10Hz 0.00743785 0.0345823
+ 5.51e+10Hz 0.00745068 0.0346429
+ 5.52e+10Hz 0.00746353 0.0347034
+ 5.53e+10Hz 0.0074764 0.0347639
+ 5.54e+10Hz 0.00748929 0.0348244
+ 5.55e+10Hz 0.0075022 0.0348849
+ 5.56e+10Hz 0.00751513 0.0349454
+ 5.57e+10Hz 0.00752808 0.0350059
+ 5.58e+10Hz 0.00754105 0.0350664
+ 5.59e+10Hz 0.00755405 0.0351268
+ 5.6e+10Hz 0.00756706 0.0351873
+ 5.61e+10Hz 0.00758009 0.0352477
+ 5.62e+10Hz 0.00759315 0.0353082
+ 5.63e+10Hz 0.00760622 0.0353686
+ 5.64e+10Hz 0.00761931 0.035429
+ 5.65e+10Hz 0.00763242 0.0354894
+ 5.66e+10Hz 0.00764556 0.0355499
+ 5.67e+10Hz 0.00765871 0.0356103
+ 5.68e+10Hz 0.00767188 0.0356707
+ 5.69e+10Hz 0.00768508 0.0357311
+ 5.7e+10Hz 0.00769829 0.0357914
+ 5.71e+10Hz 0.00771152 0.0358518
+ 5.72e+10Hz 0.00772477 0.0359122
+ 5.73e+10Hz 0.00773804 0.0359725
+ 5.74e+10Hz 0.00775133 0.0360329
+ 5.75e+10Hz 0.00776464 0.0360932
+ 5.76e+10Hz 0.00777797 0.0361535
+ 5.77e+10Hz 0.00779132 0.0362138
+ 5.78e+10Hz 0.00780469 0.0362742
+ 5.79e+10Hz 0.00781808 0.0363345
+ 5.8e+10Hz 0.00783148 0.0363948
+ 5.81e+10Hz 0.00784491 0.0364551
+ 5.82e+10Hz 0.00785836 0.0365153
+ 5.83e+10Hz 0.00787182 0.0365756
+ 5.84e+10Hz 0.0078853 0.0366359
+ 5.85e+10Hz 0.00789881 0.0366961
+ 5.86e+10Hz 0.00791233 0.0367564
+ 5.87e+10Hz 0.00792587 0.0368166
+ 5.88e+10Hz 0.00793943 0.0368768
+ 5.89e+10Hz 0.007953 0.036937
+ 5.9e+10Hz 0.0079666 0.0369973
+ 5.91e+10Hz 0.00798022 0.0370575
+ 5.92e+10Hz 0.00799385 0.0371177
+ 5.93e+10Hz 0.0080075 0.0371778
+ 5.94e+10Hz 0.00802117 0.037238
+ 5.95e+10Hz 0.00803486 0.0372982
+ 5.96e+10Hz 0.00804857 0.0373583
+ 5.97e+10Hz 0.0080623 0.0374185
+ 5.98e+10Hz 0.00807604 0.0374787
+ 5.99e+10Hz 0.00808981 0.0375388
+ 6e+10Hz 0.00810359 0.0375989
+ 6.01e+10Hz 0.00811739 0.037659
+ 6.02e+10Hz 0.00813121 0.0377191
+ 6.03e+10Hz 0.00814504 0.0377793
+ 6.04e+10Hz 0.0081589 0.0378393
+ 6.05e+10Hz 0.00817277 0.0378994
+ 6.06e+10Hz 0.00818666 0.0379595
+ 6.07e+10Hz 0.00820057 0.0380196
+ 6.08e+10Hz 0.0082145 0.0380796
+ 6.09e+10Hz 0.00822844 0.0381397
+ 6.1e+10Hz 0.0082424 0.0381997
+ 6.11e+10Hz 0.00825638 0.0382598
+ 6.12e+10Hz 0.00827038 0.0383198
+ 6.13e+10Hz 0.0082844 0.0383798
+ 6.14e+10Hz 0.00829843 0.0384398
+ 6.15e+10Hz 0.00831248 0.0384998
+ 6.16e+10Hz 0.00832655 0.0385598
+ 6.17e+10Hz 0.00834064 0.0386198
+ 6.18e+10Hz 0.00835475 0.0386798
+ 6.19e+10Hz 0.00836887 0.0387398
+ 6.2e+10Hz 0.00838301 0.0387997
+ 6.21e+10Hz 0.00839717 0.0388597
+ 6.22e+10Hz 0.00841135 0.0389196
+ 6.23e+10Hz 0.00842554 0.0389796
+ 6.24e+10Hz 0.00843975 0.0390395
+ 6.25e+10Hz 0.00845398 0.0390994
+ 6.26e+10Hz 0.00846822 0.0391594
+ 6.27e+10Hz 0.00848249 0.0392193
+ 6.28e+10Hz 0.00849677 0.0392792
+ 6.29e+10Hz 0.00851107 0.0393391
+ 6.3e+10Hz 0.00852538 0.039399
+ 6.31e+10Hz 0.00853972 0.0394588
+ 6.32e+10Hz 0.00855407 0.0395187
+ 6.33e+10Hz 0.00856843 0.0395786
+ 6.34e+10Hz 0.00858282 0.0396384
+ 6.35e+10Hz 0.00859722 0.0396983
+ 6.36e+10Hz 0.00861164 0.0397581
+ 6.37e+10Hz 0.00862608 0.0398179
+ 6.38e+10Hz 0.00864054 0.0398778
+ 6.39e+10Hz 0.00865501 0.0399376
+ 6.4e+10Hz 0.0086695 0.0399974
+ 6.41e+10Hz 0.00868401 0.0400572
+ 6.42e+10Hz 0.00869854 0.040117
+ 6.43e+10Hz 0.00871308 0.0401768
+ 6.44e+10Hz 0.00872764 0.0402366
+ 6.45e+10Hz 0.00874221 0.0402964
+ 6.46e+10Hz 0.00875681 0.0403561
+ 6.47e+10Hz 0.00877142 0.0404159
+ 6.48e+10Hz 0.00878605 0.0404757
+ 6.49e+10Hz 0.0088007 0.0405354
+ 6.5e+10Hz 0.00881536 0.0405951
+ 6.51e+10Hz 0.00883005 0.0406549
+ 6.52e+10Hz 0.00884474 0.0407146
+ 6.53e+10Hz 0.00885946 0.0407743
+ 6.54e+10Hz 0.0088742 0.040834
+ 6.55e+10Hz 0.00888895 0.0408937
+ 6.56e+10Hz 0.00890372 0.0409535
+ 6.57e+10Hz 0.00891851 0.0410131
+ 6.58e+10Hz 0.00893331 0.0410728
+ 6.59e+10Hz 0.00894813 0.0411325
+ 6.6e+10Hz 0.00896297 0.0411922
+ 6.61e+10Hz 0.00897783 0.0412519
+ 6.62e+10Hz 0.00899271 0.0413115
+ 6.63e+10Hz 0.0090076 0.0413712
+ 6.64e+10Hz 0.00902251 0.0414308
+ 6.65e+10Hz 0.00903744 0.0414905
+ 6.66e+10Hz 0.00905239 0.0415501
+ 6.67e+10Hz 0.00906735 0.0416098
+ 6.68e+10Hz 0.00908233 0.0416694
+ 6.69e+10Hz 0.00909733 0.041729
+ 6.7e+10Hz 0.00911235 0.0417886
+ 6.71e+10Hz 0.00912739 0.0418482
+ 6.72e+10Hz 0.00914244 0.0419078
+ 6.73e+10Hz 0.00915751 0.0419674
+ 6.74e+10Hz 0.0091726 0.042027
+ 6.75e+10Hz 0.00918771 0.0420866
+ 6.76e+10Hz 0.00920283 0.0421462
+ 6.77e+10Hz 0.00921798 0.0422057
+ 6.78e+10Hz 0.00923314 0.0422653
+ 6.79e+10Hz 0.00924832 0.0423248
+ 6.8e+10Hz 0.00926352 0.0423844
+ 6.81e+10Hz 0.00927873 0.0424439
+ 6.82e+10Hz 0.00929397 0.0425035
+ 6.83e+10Hz 0.00930922 0.042563
+ 6.84e+10Hz 0.00932449 0.0426225
+ 6.85e+10Hz 0.00933978 0.042682
+ 6.86e+10Hz 0.00935509 0.0427416
+ 6.87e+10Hz 0.00937042 0.0428011
+ 6.88e+10Hz 0.00938576 0.0428606
+ 6.89e+10Hz 0.00940113 0.0429201
+ 6.9e+10Hz 0.00941651 0.0429796
+ 6.91e+10Hz 0.00943191 0.0430391
+ 6.92e+10Hz 0.00944733 0.0430985
+ 6.93e+10Hz 0.00946277 0.043158
+ 6.94e+10Hz 0.00947823 0.0432175
+ 6.95e+10Hz 0.0094937 0.0432769
+ 6.96e+10Hz 0.0095092 0.0433364
+ 6.97e+10Hz 0.00952471 0.0433958
+ 6.98e+10Hz 0.00954024 0.0434553
+ 6.99e+10Hz 0.0095558 0.0435147
+ 7e+10Hz 0.00957137 0.0435742
+ 7.01e+10Hz 0.00958696 0.0436336
+ 7.02e+10Hz 0.00960257 0.043693
+ 7.03e+10Hz 0.00961819 0.0437524
+ 7.04e+10Hz 0.00963384 0.0438118
+ 7.05e+10Hz 0.00964951 0.0438712
+ 7.06e+10Hz 0.00966519 0.0439306
+ 7.07e+10Hz 0.0096809 0.04399
+ 7.08e+10Hz 0.00969662 0.0440494
+ 7.09e+10Hz 0.00971237 0.0441088
+ 7.1e+10Hz 0.00972813 0.0441682
+ 7.11e+10Hz 0.00974391 0.0442275
+ 7.12e+10Hz 0.00975971 0.0442869
+ 7.13e+10Hz 0.00977554 0.0443462
+ 7.14e+10Hz 0.00979138 0.0444056
+ 7.15e+10Hz 0.00980724 0.0444649
+ 7.16e+10Hz 0.00982312 0.0445243
+ 7.17e+10Hz 0.00983902 0.0445836
+ 7.18e+10Hz 0.00985494 0.0446429
+ 7.19e+10Hz 0.00987088 0.0447022
+ 7.2e+10Hz 0.00988684 0.0447616
+ 7.21e+10Hz 0.00990282 0.0448209
+ 7.22e+10Hz 0.00991882 0.0448802
+ 7.23e+10Hz 0.00993484 0.0449395
+ 7.24e+10Hz 0.00995088 0.0449987
+ 7.25e+10Hz 0.00996694 0.045058
+ 7.26e+10Hz 0.00998302 0.0451173
+ 7.27e+10Hz 0.00999912 0.0451766
+ 7.28e+10Hz 0.0100152 0.0452358
+ 7.29e+10Hz 0.0100314 0.0452951
+ 7.3e+10Hz 0.0100475 0.0453544
+ 7.31e+10Hz 0.0100637 0.0454136
+ 7.32e+10Hz 0.0100799 0.0454728
+ 7.33e+10Hz 0.0100961 0.0455321
+ 7.34e+10Hz 0.0101124 0.0455913
+ 7.35e+10Hz 0.0101286 0.0456505
+ 7.36e+10Hz 0.0101449 0.0457097
+ 7.37e+10Hz 0.0101612 0.0457689
+ 7.38e+10Hz 0.0101776 0.0458281
+ 7.39e+10Hz 0.0101939 0.0458873
+ 7.4e+10Hz 0.0102103 0.0459465
+ 7.41e+10Hz 0.0102266 0.0460057
+ 7.42e+10Hz 0.0102431 0.0460648
+ 7.43e+10Hz 0.0102595 0.046124
+ 7.44e+10Hz 0.0102759 0.0461832
+ 7.45e+10Hz 0.0102924 0.0462423
+ 7.46e+10Hz 0.0103089 0.0463015
+ 7.47e+10Hz 0.0103254 0.0463606
+ 7.48e+10Hz 0.0103419 0.0464197
+ 7.49e+10Hz 0.0103585 0.0464789
+ 7.5e+10Hz 0.010375 0.046538
+ 7.51e+10Hz 0.0103916 0.0465971
+ 7.52e+10Hz 0.0104082 0.0466562
+ 7.53e+10Hz 0.0104249 0.0467153
+ 7.54e+10Hz 0.0104415 0.0467743
+ 7.55e+10Hz 0.0104582 0.0468334
+ 7.56e+10Hz 0.0104749 0.0468925
+ 7.57e+10Hz 0.0104916 0.0469516
+ 7.58e+10Hz 0.0105083 0.0470106
+ 7.59e+10Hz 0.0105251 0.0470697
+ 7.6e+10Hz 0.0105419 0.0471287
+ 7.61e+10Hz 0.0105587 0.0471877
+ 7.62e+10Hz 0.0105755 0.0472468
+ 7.63e+10Hz 0.0105923 0.0473058
+ 7.64e+10Hz 0.0106092 0.0473648
+ 7.65e+10Hz 0.0106261 0.0474238
+ 7.66e+10Hz 0.010643 0.0474828
+ 7.67e+10Hz 0.0106599 0.0475418
+ 7.68e+10Hz 0.0106768 0.0476008
+ 7.69e+10Hz 0.0106938 0.0476597
+ 7.7e+10Hz 0.0107108 0.0477187
+ 7.71e+10Hz 0.0107278 0.0477776
+ 7.72e+10Hz 0.0107448 0.0478366
+ 7.73e+10Hz 0.0107619 0.0478955
+ 7.74e+10Hz 0.010779 0.0479545
+ 7.75e+10Hz 0.010796 0.0480134
+ 7.76e+10Hz 0.0108132 0.0480723
+ 7.77e+10Hz 0.0108303 0.0481312
+ 7.78e+10Hz 0.0108474 0.0481901
+ 7.79e+10Hz 0.0108646 0.048249
+ 7.8e+10Hz 0.0108818 0.0483079
+ 7.81e+10Hz 0.010899 0.0483668
+ 7.82e+10Hz 0.0109163 0.0484256
+ 7.83e+10Hz 0.0109335 0.0484845
+ 7.84e+10Hz 0.0109508 0.0485433
+ 7.85e+10Hz 0.0109681 0.0486021
+ 7.86e+10Hz 0.0109854 0.048661
+ 7.87e+10Hz 0.0110028 0.0487198
+ 7.88e+10Hz 0.0110201 0.0487786
+ 7.89e+10Hz 0.0110375 0.0488374
+ 7.9e+10Hz 0.0110549 0.0488962
+ 7.91e+10Hz 0.0110723 0.048955
+ 7.92e+10Hz 0.0110898 0.0490138
+ 7.93e+10Hz 0.0111072 0.0490725
+ 7.94e+10Hz 0.0111247 0.0491313
+ 7.95e+10Hz 0.0111422 0.04919
+ 7.96e+10Hz 0.0111597 0.0492488
+ 7.97e+10Hz 0.0111773 0.0493075
+ 7.98e+10Hz 0.0111948 0.0493662
+ 7.99e+10Hz 0.0112124 0.049425
+ 8e+10Hz 0.01123 0.0494837
+ 8.01e+10Hz 0.0112477 0.0495423
+ 8.02e+10Hz 0.0112653 0.049601
+ 8.03e+10Hz 0.011283 0.0496597
+ 8.04e+10Hz 0.0113007 0.0497184
+ 8.05e+10Hz 0.0113184 0.049777
+ 8.06e+10Hz 0.0113361 0.0498357
+ 8.07e+10Hz 0.0113538 0.0498943
+ 8.08e+10Hz 0.0113716 0.049953
+ 8.09e+10Hz 0.0113894 0.0500116
+ 8.1e+10Hz 0.0114072 0.0500702
+ 8.11e+10Hz 0.011425 0.0501288
+ 8.12e+10Hz 0.0114429 0.0501874
+ 8.13e+10Hz 0.0114608 0.050246
+ 8.14e+10Hz 0.0114786 0.0503045
+ 8.15e+10Hz 0.0114965 0.0503631
+ 8.16e+10Hz 0.0115145 0.0504216
+ 8.17e+10Hz 0.0115324 0.0504802
+ 8.18e+10Hz 0.0115504 0.0505387
+ 8.19e+10Hz 0.0115684 0.0505973
+ 8.2e+10Hz 0.0115864 0.0506558
+ 8.21e+10Hz 0.0116044 0.0507143
+ 8.22e+10Hz 0.0116224 0.0507728
+ 8.23e+10Hz 0.0116405 0.0508313
+ 8.24e+10Hz 0.0116586 0.0508897
+ 8.25e+10Hz 0.0116767 0.0509482
+ 8.26e+10Hz 0.0116948 0.0510067
+ 8.27e+10Hz 0.011713 0.0510651
+ 8.28e+10Hz 0.0117311 0.0511235
+ 8.29e+10Hz 0.0117493 0.051182
+ 8.3e+10Hz 0.0117675 0.0512404
+ 8.31e+10Hz 0.0117857 0.0512988
+ 8.32e+10Hz 0.011804 0.0513572
+ 8.33e+10Hz 0.0118222 0.0514156
+ 8.34e+10Hz 0.0118405 0.0514739
+ 8.35e+10Hz 0.0118588 0.0515323
+ 8.36e+10Hz 0.0118771 0.0515907
+ 8.37e+10Hz 0.0118955 0.051649
+ 8.38e+10Hz 0.0119138 0.0517074
+ 8.39e+10Hz 0.0119322 0.0517657
+ 8.4e+10Hz 0.0119506 0.051824
+ 8.41e+10Hz 0.011969 0.0518823
+ 8.42e+10Hz 0.0119874 0.0519406
+ 8.43e+10Hz 0.0120059 0.0519989
+ 8.44e+10Hz 0.0120243 0.0520572
+ 8.45e+10Hz 0.0120428 0.0521155
+ 8.46e+10Hz 0.0120613 0.0521737
+ 8.47e+10Hz 0.0120798 0.052232
+ 8.48e+10Hz 0.0120984 0.0522902
+ 8.49e+10Hz 0.0121169 0.0523485
+ 8.5e+10Hz 0.0121355 0.0524067
+ 8.51e+10Hz 0.0121541 0.0524649
+ 8.52e+10Hz 0.0121727 0.0525231
+ 8.53e+10Hz 0.0121914 0.0525813
+ 8.54e+10Hz 0.01221 0.0526395
+ 8.55e+10Hz 0.0122287 0.0526977
+ 8.56e+10Hz 0.0122474 0.0527558
+ 8.57e+10Hz 0.0122661 0.052814
+ 8.58e+10Hz 0.0122848 0.0528721
+ 8.59e+10Hz 0.0123035 0.0529303
+ 8.6e+10Hz 0.0123223 0.0529884
+ 8.61e+10Hz 0.0123411 0.0530465
+ 8.62e+10Hz 0.0123599 0.0531046
+ 8.63e+10Hz 0.0123787 0.0531627
+ 8.64e+10Hz 0.0123976 0.0532208
+ 8.65e+10Hz 0.0124164 0.0532789
+ 8.66e+10Hz 0.0124353 0.053337
+ 8.67e+10Hz 0.0124542 0.053395
+ 8.68e+10Hz 0.0124731 0.0534531
+ 8.69e+10Hz 0.012492 0.0535111
+ 8.7e+10Hz 0.0125109 0.0535692
+ 8.71e+10Hz 0.0125299 0.0536272
+ 8.72e+10Hz 0.0125489 0.0536852
+ 8.73e+10Hz 0.0125679 0.0537432
+ 8.74e+10Hz 0.0125869 0.0538012
+ 8.75e+10Hz 0.0126059 0.0538592
+ 8.76e+10Hz 0.012625 0.0539172
+ 8.77e+10Hz 0.012644 0.0539751
+ 8.78e+10Hz 0.0126631 0.0540331
+ 8.79e+10Hz 0.0126822 0.0540911
+ 8.8e+10Hz 0.0127014 0.054149
+ 8.81e+10Hz 0.0127205 0.0542069
+ 8.82e+10Hz 0.0127397 0.0542649
+ 8.83e+10Hz 0.0127588 0.0543228
+ 8.84e+10Hz 0.012778 0.0543807
+ 8.85e+10Hz 0.0127972 0.0544386
+ 8.86e+10Hz 0.0128165 0.0544965
+ 8.87e+10Hz 0.0128357 0.0545544
+ 8.88e+10Hz 0.012855 0.0546122
+ 8.89e+10Hz 0.0128743 0.0546701
+ 8.9e+10Hz 0.0128936 0.0547279
+ 8.91e+10Hz 0.0129129 0.0547858
+ 8.92e+10Hz 0.0129322 0.0548436
+ 8.93e+10Hz 0.0129516 0.0549014
+ 8.94e+10Hz 0.0129709 0.0549593
+ 8.95e+10Hz 0.0129903 0.0550171
+ 8.96e+10Hz 0.0130097 0.0550749
+ 8.97e+10Hz 0.0130292 0.0551327
+ 8.98e+10Hz 0.0130486 0.0551905
+ 8.99e+10Hz 0.0130681 0.0552482
+ 9e+10Hz 0.0130875 0.055306
+ 9.01e+10Hz 0.013107 0.0553638
+ 9.02e+10Hz 0.0131265 0.0554215
+ 9.03e+10Hz 0.0131461 0.0554793
+ 9.04e+10Hz 0.0131656 0.055537
+ 9.05e+10Hz 0.0131852 0.0555947
+ 9.06e+10Hz 0.0132048 0.0556525
+ 9.07e+10Hz 0.0132244 0.0557102
+ 9.08e+10Hz 0.013244 0.0557679
+ 9.09e+10Hz 0.0132636 0.0558256
+ 9.1e+10Hz 0.0132833 0.0558833
+ 9.11e+10Hz 0.013303 0.055941
+ 9.12e+10Hz 0.0133227 0.0559986
+ 9.13e+10Hz 0.0133424 0.0560563
+ 9.14e+10Hz 0.0133621 0.056114
+ 9.15e+10Hz 0.0133818 0.0561716
+ 9.16e+10Hz 0.0134016 0.0562292
+ 9.17e+10Hz 0.0134214 0.0562869
+ 9.18e+10Hz 0.0134412 0.0563445
+ 9.19e+10Hz 0.013461 0.0564021
+ 9.2e+10Hz 0.0134808 0.0564597
+ 9.21e+10Hz 0.0135007 0.0565173
+ 9.22e+10Hz 0.0135205 0.0565749
+ 9.23e+10Hz 0.0135404 0.0566325
+ 9.24e+10Hz 0.0135604 0.0566901
+ 9.25e+10Hz 0.0135803 0.0567476
+ 9.26e+10Hz 0.0136002 0.0568052
+ 9.27e+10Hz 0.0136202 0.0568628
+ 9.28e+10Hz 0.0136402 0.0569203
+ 9.29e+10Hz 0.0136602 0.0569778
+ 9.3e+10Hz 0.0136802 0.0570354
+ 9.31e+10Hz 0.0137002 0.0570929
+ 9.32e+10Hz 0.0137203 0.0571504
+ 9.33e+10Hz 0.0137403 0.0572079
+ 9.34e+10Hz 0.0137604 0.0572654
+ 9.35e+10Hz 0.0137805 0.0573229
+ 9.36e+10Hz 0.0138006 0.0573804
+ 9.37e+10Hz 0.0138208 0.0574379
+ 9.38e+10Hz 0.013841 0.0574954
+ 9.39e+10Hz 0.0138611 0.0575528
+ 9.4e+10Hz 0.0138814 0.0576103
+ 9.41e+10Hz 0.0139016 0.0576677
+ 9.42e+10Hz 0.0139218 0.0577252
+ 9.43e+10Hz 0.0139421 0.0577826
+ 9.44e+10Hz 0.0139623 0.05784
+ 9.45e+10Hz 0.0139826 0.0578974
+ 9.46e+10Hz 0.0140029 0.0579549
+ 9.47e+10Hz 0.0140233 0.0580123
+ 9.48e+10Hz 0.0140436 0.0580696
+ 9.49e+10Hz 0.014064 0.058127
+ 9.5e+10Hz 0.0140844 0.0581844
+ 9.51e+10Hz 0.0141048 0.0582418
+ 9.52e+10Hz 0.0141252 0.0582992
+ 9.53e+10Hz 0.0141457 0.0583565
+ 9.54e+10Hz 0.0141661 0.0584139
+ 9.55e+10Hz 0.0141866 0.0584712
+ 9.56e+10Hz 0.0142071 0.0585285
+ 9.57e+10Hz 0.0142276 0.0585859
+ 9.58e+10Hz 0.0142482 0.0586432
+ 9.59e+10Hz 0.0142687 0.0587005
+ 9.6e+10Hz 0.0142893 0.0587578
+ 9.61e+10Hz 0.0143099 0.0588151
+ 9.62e+10Hz 0.0143305 0.0588724
+ 9.63e+10Hz 0.0143512 0.0589297
+ 9.64e+10Hz 0.0143718 0.0589869
+ 9.65e+10Hz 0.0143925 0.0590442
+ 9.66e+10Hz 0.0144132 0.0591014
+ 9.67e+10Hz 0.0144339 0.0591587
+ 9.68e+10Hz 0.0144546 0.0592159
+ 9.69e+10Hz 0.0144754 0.0592732
+ 9.7e+10Hz 0.0144961 0.0593304
+ 9.71e+10Hz 0.014517 0.0593876
+ 9.72e+10Hz 0.0145378 0.0594448
+ 9.73e+10Hz 0.0145586 0.059502
+ 9.74e+10Hz 0.0145794 0.0595592
+ 9.75e+10Hz 0.0146003 0.0596164
+ 9.76e+10Hz 0.0146212 0.0596736
+ 9.77e+10Hz 0.0146421 0.0597307
+ 9.78e+10Hz 0.014663 0.0597879
+ 9.79e+10Hz 0.014684 0.059845
+ 9.8e+10Hz 0.014705 0.0599022
+ 9.81e+10Hz 0.0147259 0.0599593
+ 9.82e+10Hz 0.014747 0.0600165
+ 9.83e+10Hz 0.014768 0.0600736
+ 9.84e+10Hz 0.014789 0.0601307
+ 9.85e+10Hz 0.0148101 0.0601878
+ 9.86e+10Hz 0.0148312 0.0602449
+ 9.87e+10Hz 0.0148523 0.060302
+ 9.88e+10Hz 0.0148734 0.060359
+ 9.89e+10Hz 0.0148946 0.0604161
+ 9.9e+10Hz 0.0149157 0.0604732
+ 9.91e+10Hz 0.0149369 0.0605302
+ 9.92e+10Hz 0.0149581 0.0605873
+ 9.93e+10Hz 0.0149794 0.0606443
+ 9.94e+10Hz 0.0150006 0.0607013
+ 9.95e+10Hz 0.0150219 0.0607583
+ 9.96e+10Hz 0.0150432 0.0608153
+ 9.97e+10Hz 0.0150645 0.0608723
+ 9.98e+10Hz 0.0150858 0.0609293
+ 9.99e+10Hz 0.0151072 0.0609863
+ 1e+11Hz 0.0151285 0.0610433
+ 1.001e+11Hz 0.0151499 0.0611003
+ 1.002e+11Hz 0.0151713 0.0611572
+ 1.003e+11Hz 0.0151927 0.0612141
+ 1.004e+11Hz 0.0152142 0.0612711
+ 1.005e+11Hz 0.0152357 0.061328
+ 1.006e+11Hz 0.0152572 0.0613849
+ 1.007e+11Hz 0.0152787 0.0614418
+ 1.008e+11Hz 0.0153002 0.0614987
+ 1.009e+11Hz 0.0153218 0.0615556
+ 1.01e+11Hz 0.0153433 0.0616125
+ 1.011e+11Hz 0.0153649 0.0616693
+ 1.012e+11Hz 0.0153865 0.0617262
+ 1.013e+11Hz 0.0154081 0.0617831
+ 1.014e+11Hz 0.0154298 0.0618399
+ 1.015e+11Hz 0.0154515 0.0618967
+ 1.016e+11Hz 0.0154731 0.0619536
+ 1.017e+11Hz 0.0154949 0.0620104
+ 1.018e+11Hz 0.0155166 0.0620672
+ 1.019e+11Hz 0.0155383 0.0621239
+ 1.02e+11Hz 0.0155601 0.0621807
+ 1.021e+11Hz 0.0155819 0.0622375
+ 1.022e+11Hz 0.0156037 0.0622943
+ 1.023e+11Hz 0.0156255 0.062351
+ 1.024e+11Hz 0.0156474 0.0624077
+ 1.025e+11Hz 0.0156693 0.0624645
+ 1.026e+11Hz 0.0156912 0.0625212
+ 1.027e+11Hz 0.0157131 0.0625779
+ 1.028e+11Hz 0.015735 0.0626346
+ 1.029e+11Hz 0.0157569 0.0626913
+ 1.03e+11Hz 0.0157789 0.0627479
+ 1.031e+11Hz 0.0158009 0.0628046
+ 1.032e+11Hz 0.0158229 0.0628613
+ 1.033e+11Hz 0.0158449 0.0629179
+ 1.034e+11Hz 0.015867 0.0629745
+ 1.035e+11Hz 0.015889 0.0630312
+ 1.036e+11Hz 0.0159111 0.0630878
+ 1.037e+11Hz 0.0159332 0.0631444
+ 1.038e+11Hz 0.0159554 0.063201
+ 1.039e+11Hz 0.0159775 0.0632575
+ 1.04e+11Hz 0.0159997 0.0633141
+ 1.041e+11Hz 0.0160219 0.0633707
+ 1.042e+11Hz 0.0160441 0.0634272
+ 1.043e+11Hz 0.0160663 0.0634837
+ 1.044e+11Hz 0.0160885 0.0635403
+ 1.045e+11Hz 0.0161108 0.0635968
+ 1.046e+11Hz 0.0161331 0.0636533
+ 1.047e+11Hz 0.0161554 0.0637098
+ 1.048e+11Hz 0.0161777 0.0637662
+ 1.049e+11Hz 0.0162 0.0638227
+ 1.05e+11Hz 0.0162224 0.0638791
+ 1.051e+11Hz 0.0162447 0.0639356
+ 1.052e+11Hz 0.0162671 0.063992
+ 1.053e+11Hz 0.0162896 0.0640484
+ 1.054e+11Hz 0.016312 0.0641049
+ 1.055e+11Hz 0.0163344 0.0641613
+ 1.056e+11Hz 0.0163569 0.0642176
+ 1.057e+11Hz 0.0163794 0.064274
+ 1.058e+11Hz 0.0164019 0.0643304
+ 1.059e+11Hz 0.0164244 0.0643867
+ 1.06e+11Hz 0.016447 0.0644431
+ 1.061e+11Hz 0.0164695 0.0644994
+ 1.062e+11Hz 0.0164921 0.0645557
+ 1.063e+11Hz 0.0165147 0.064612
+ 1.064e+11Hz 0.0165373 0.0646683
+ 1.065e+11Hz 0.01656 0.0647246
+ 1.066e+11Hz 0.0165826 0.0647808
+ 1.067e+11Hz 0.0166053 0.0648371
+ 1.068e+11Hz 0.016628 0.0648933
+ 1.069e+11Hz 0.0166507 0.0649495
+ 1.07e+11Hz 0.0166734 0.0650058
+ 1.071e+11Hz 0.0166961 0.065062
+ 1.072e+11Hz 0.0167189 0.0651182
+ 1.073e+11Hz 0.0167417 0.0651743
+ 1.074e+11Hz 0.0167645 0.0652305
+ 1.075e+11Hz 0.0167873 0.0652867
+ 1.076e+11Hz 0.0168101 0.0653428
+ 1.077e+11Hz 0.016833 0.0653989
+ 1.078e+11Hz 0.0168558 0.0654551
+ 1.079e+11Hz 0.0168787 0.0655112
+ 1.08e+11Hz 0.0169016 0.0655673
+ 1.081e+11Hz 0.0169246 0.0656234
+ 1.082e+11Hz 0.0169475 0.0656794
+ 1.083e+11Hz 0.0169704 0.0657355
+ 1.084e+11Hz 0.0169934 0.0657915
+ 1.085e+11Hz 0.0170164 0.0658476
+ 1.086e+11Hz 0.0170394 0.0659036
+ 1.087e+11Hz 0.0170624 0.0659596
+ 1.088e+11Hz 0.0170855 0.0660156
+ 1.089e+11Hz 0.0171085 0.0660716
+ 1.09e+11Hz 0.0171316 0.0661276
+ 1.091e+11Hz 0.0171547 0.0661835
+ 1.092e+11Hz 0.0171778 0.0662395
+ 1.093e+11Hz 0.0172009 0.0662954
+ 1.094e+11Hz 0.017224 0.0663514
+ 1.095e+11Hz 0.0172472 0.0664073
+ 1.096e+11Hz 0.0172704 0.0664632
+ 1.097e+11Hz 0.0172936 0.0665191
+ 1.098e+11Hz 0.0173167 0.0665749
+ 1.099e+11Hz 0.01734 0.0666308
+ 1.1e+11Hz 0.0173632 0.0666867
+ 1.101e+11Hz 0.0173865 0.0667425
+ 1.102e+11Hz 0.0174097 0.0667984
+ 1.103e+11Hz 0.017433 0.0668542
+ 1.104e+11Hz 0.0174563 0.06691
+ 1.105e+11Hz 0.0174796 0.0669658
+ 1.106e+11Hz 0.017503 0.0670216
+ 1.107e+11Hz 0.0175263 0.0670773
+ 1.108e+11Hz 0.0175497 0.0671331
+ 1.109e+11Hz 0.017573 0.0671888
+ 1.11e+11Hz 0.0175964 0.0672446
+ 1.111e+11Hz 0.0176198 0.0673003
+ 1.112e+11Hz 0.0176433 0.067356
+ 1.113e+11Hz 0.0176667 0.0674117
+ 1.114e+11Hz 0.0176902 0.0674674
+ 1.115e+11Hz 0.0177137 0.0675231
+ 1.116e+11Hz 0.0177371 0.0675788
+ 1.117e+11Hz 0.0177606 0.0676344
+ 1.118e+11Hz 0.0177842 0.0676901
+ 1.119e+11Hz 0.0178077 0.0677457
+ 1.12e+11Hz 0.0178312 0.0678013
+ 1.121e+11Hz 0.0178548 0.0678569
+ 1.122e+11Hz 0.0178784 0.0679125
+ 1.123e+11Hz 0.017902 0.0679681
+ 1.124e+11Hz 0.0179256 0.0680237
+ 1.125e+11Hz 0.0179492 0.0680793
+ 1.126e+11Hz 0.0179729 0.0681348
+ 1.127e+11Hz 0.0179965 0.0681904
+ 1.128e+11Hz 0.0180202 0.0682459
+ 1.129e+11Hz 0.0180439 0.0683014
+ 1.13e+11Hz 0.0180676 0.0683569
+ 1.131e+11Hz 0.0180913 0.0684124
+ 1.132e+11Hz 0.018115 0.0684679
+ 1.133e+11Hz 0.0181388 0.0685234
+ 1.134e+11Hz 0.0181625 0.0685789
+ 1.135e+11Hz 0.0181863 0.0686344
+ 1.136e+11Hz 0.0182101 0.0686898
+ 1.137e+11Hz 0.0182339 0.0687452
+ 1.138e+11Hz 0.0182577 0.0688007
+ 1.139e+11Hz 0.0182816 0.0688561
+ 1.14e+11Hz 0.0183054 0.0689115
+ 1.141e+11Hz 0.0183293 0.0689669
+ 1.142e+11Hz 0.0183531 0.0690223
+ 1.143e+11Hz 0.018377 0.0690777
+ 1.144e+11Hz 0.018401 0.069133
+ 1.145e+11Hz 0.0184249 0.0691884
+ 1.146e+11Hz 0.0184488 0.0692437
+ 1.147e+11Hz 0.0184728 0.0692991
+ 1.148e+11Hz 0.0184967 0.0693544
+ 1.149e+11Hz 0.0185207 0.0694097
+ 1.15e+11Hz 0.0185447 0.069465
+ 1.151e+11Hz 0.0185687 0.0695203
+ 1.152e+11Hz 0.0185928 0.0695756
+ 1.153e+11Hz 0.0186168 0.0696309
+ 1.154e+11Hz 0.0186409 0.0696862
+ 1.155e+11Hz 0.018665 0.0697414
+ 1.156e+11Hz 0.0186891 0.0697967
+ 1.157e+11Hz 0.0187132 0.0698519
+ 1.158e+11Hz 0.0187373 0.0699071
+ 1.159e+11Hz 0.0187614 0.0699624
+ 1.16e+11Hz 0.0187856 0.0700176
+ 1.161e+11Hz 0.0188097 0.0700728
+ 1.162e+11Hz 0.0188339 0.070128
+ 1.163e+11Hz 0.0188581 0.0701831
+ 1.164e+11Hz 0.0188823 0.0702383
+ 1.165e+11Hz 0.0189066 0.0702935
+ 1.166e+11Hz 0.0189308 0.0703486
+ 1.167e+11Hz 0.0189551 0.0704038
+ 1.168e+11Hz 0.0189793 0.0704589
+ 1.169e+11Hz 0.0190036 0.070514
+ 1.17e+11Hz 0.0190279 0.0705692
+ 1.171e+11Hz 0.0190523 0.0706243
+ 1.172e+11Hz 0.0190766 0.0706794
+ 1.173e+11Hz 0.0191009 0.0707345
+ 1.174e+11Hz 0.0191253 0.0707896
+ 1.175e+11Hz 0.0191497 0.0708446
+ 1.176e+11Hz 0.0191741 0.0708997
+ 1.177e+11Hz 0.0191985 0.0709548
+ 1.178e+11Hz 0.0192229 0.0710098
+ 1.179e+11Hz 0.0192474 0.0710648
+ 1.18e+11Hz 0.0192719 0.0711199
+ 1.181e+11Hz 0.0192964 0.0711749
+ 1.182e+11Hz 0.0193208 0.0712299
+ 1.183e+11Hz 0.0193454 0.0712849
+ 1.184e+11Hz 0.0193699 0.0713399
+ 1.185e+11Hz 0.0193944 0.0713949
+ 1.186e+11Hz 0.019419 0.0714499
+ 1.187e+11Hz 0.0194436 0.0715048
+ 1.188e+11Hz 0.0194682 0.0715598
+ 1.189e+11Hz 0.0194928 0.0716148
+ 1.19e+11Hz 0.0195174 0.0716697
+ 1.191e+11Hz 0.0195421 0.0717247
+ 1.192e+11Hz 0.0195667 0.0717796
+ 1.193e+11Hz 0.0195914 0.0718345
+ 1.194e+11Hz 0.0196161 0.0718894
+ 1.195e+11Hz 0.0196408 0.0719443
+ 1.196e+11Hz 0.0196655 0.0719992
+ 1.197e+11Hz 0.0196903 0.0720541
+ 1.198e+11Hz 0.0197151 0.072109
+ 1.199e+11Hz 0.0197398 0.0721638
+ 1.2e+11Hz 0.0197646 0.0722187
+ 1.201e+11Hz 0.0197895 0.0722735
+ 1.202e+11Hz 0.0198143 0.0723284
+ 1.203e+11Hz 0.0198391 0.0723832
+ 1.204e+11Hz 0.019864 0.072438
+ 1.205e+11Hz 0.0198889 0.0724928
+ 1.206e+11Hz 0.0199138 0.0725477
+ 1.207e+11Hz 0.0199387 0.0726024
+ 1.208e+11Hz 0.0199637 0.0726572
+ 1.209e+11Hz 0.0199886 0.072712
+ 1.21e+11Hz 0.0200136 0.0727668
+ 1.211e+11Hz 0.0200386 0.0728215
+ 1.212e+11Hz 0.0200636 0.0728763
+ 1.213e+11Hz 0.0200887 0.072931
+ 1.214e+11Hz 0.0201137 0.0729858
+ 1.215e+11Hz 0.0201388 0.0730405
+ 1.216e+11Hz 0.0201639 0.0730952
+ 1.217e+11Hz 0.020189 0.0731499
+ 1.218e+11Hz 0.0202141 0.0732046
+ 1.219e+11Hz 0.0202393 0.0732593
+ 1.22e+11Hz 0.0202644 0.073314
+ 1.221e+11Hz 0.0202896 0.0733687
+ 1.222e+11Hz 0.0203148 0.0734233
+ 1.223e+11Hz 0.02034 0.073478
+ 1.224e+11Hz 0.0203653 0.0735326
+ 1.225e+11Hz 0.0203905 0.0735872
+ 1.226e+11Hz 0.0204158 0.0736419
+ 1.227e+11Hz 0.0204411 0.0736965
+ 1.228e+11Hz 0.0204664 0.0737511
+ 1.229e+11Hz 0.0204917 0.0738057
+ 1.23e+11Hz 0.0205171 0.0738603
+ 1.231e+11Hz 0.0205425 0.0739148
+ 1.232e+11Hz 0.0205679 0.0739694
+ 1.233e+11Hz 0.0205933 0.0740239
+ 1.234e+11Hz 0.0206187 0.0740785
+ 1.235e+11Hz 0.0206442 0.074133
+ 1.236e+11Hz 0.0206697 0.0741875
+ 1.237e+11Hz 0.0206952 0.074242
+ 1.238e+11Hz 0.0207207 0.0742965
+ 1.239e+11Hz 0.0207462 0.074351
+ 1.24e+11Hz 0.0207718 0.0744055
+ 1.241e+11Hz 0.0207973 0.07446
+ 1.242e+11Hz 0.0208229 0.0745144
+ 1.243e+11Hz 0.0208486 0.0745689
+ 1.244e+11Hz 0.0208742 0.0746233
+ 1.245e+11Hz 0.0208998 0.0746777
+ 1.246e+11Hz 0.0209255 0.0747321
+ 1.247e+11Hz 0.0209512 0.0747865
+ 1.248e+11Hz 0.0209769 0.0748409
+ 1.249e+11Hz 0.0210027 0.0748953
+ 1.25e+11Hz 0.0210284 0.0749496
+ 1.251e+11Hz 0.0210542 0.075004
+ 1.252e+11Hz 0.02108 0.0750583
+ 1.253e+11Hz 0.0211058 0.0751127
+ 1.254e+11Hz 0.0211317 0.075167
+ 1.255e+11Hz 0.0211575 0.0752213
+ 1.256e+11Hz 0.0211834 0.0752755
+ 1.257e+11Hz 0.0212093 0.0753298
+ 1.258e+11Hz 0.0212352 0.0753841
+ 1.259e+11Hz 0.0212612 0.0754383
+ 1.26e+11Hz 0.0212871 0.0754926
+ 1.261e+11Hz 0.0213131 0.0755468
+ 1.262e+11Hz 0.0213391 0.075601
+ 1.263e+11Hz 0.0213651 0.0756552
+ 1.264e+11Hz 0.0213912 0.0757094
+ 1.265e+11Hz 0.0214173 0.0757636
+ 1.266e+11Hz 0.0214433 0.0758177
+ 1.267e+11Hz 0.0214695 0.0758719
+ 1.268e+11Hz 0.0214956 0.075926
+ 1.269e+11Hz 0.0215217 0.0759801
+ 1.27e+11Hz 0.0215479 0.0760342
+ 1.271e+11Hz 0.0215741 0.0760883
+ 1.272e+11Hz 0.0216003 0.0761423
+ 1.273e+11Hz 0.0216265 0.0761964
+ 1.274e+11Hz 0.0216528 0.0762504
+ 1.275e+11Hz 0.0216791 0.0763045
+ 1.276e+11Hz 0.0217054 0.0763585
+ 1.277e+11Hz 0.0217317 0.0764125
+ 1.278e+11Hz 0.021758 0.0764665
+ 1.279e+11Hz 0.0217844 0.0765204
+ 1.28e+11Hz 0.0218107 0.0765744
+ 1.281e+11Hz 0.0218371 0.0766283
+ 1.282e+11Hz 0.0218635 0.0766822
+ 1.283e+11Hz 0.02189 0.0767362
+ 1.284e+11Hz 0.0219164 0.07679
+ 1.285e+11Hz 0.0219429 0.0768439
+ 1.286e+11Hz 0.0219694 0.0768978
+ 1.287e+11Hz 0.0219959 0.0769516
+ 1.288e+11Hz 0.0220224 0.0770054
+ 1.289e+11Hz 0.022049 0.0770592
+ 1.29e+11Hz 0.0220756 0.077113
+ 1.291e+11Hz 0.0221022 0.0771668
+ 1.292e+11Hz 0.0221288 0.0772206
+ 1.293e+11Hz 0.0221554 0.0772743
+ 1.294e+11Hz 0.022182 0.077328
+ 1.295e+11Hz 0.0222087 0.0773817
+ 1.296e+11Hz 0.0222354 0.0774354
+ 1.297e+11Hz 0.0222621 0.0774891
+ 1.298e+11Hz 0.0222888 0.0775428
+ 1.299e+11Hz 0.0223156 0.0775964
+ 1.3e+11Hz 0.0223424 0.07765
+ 1.301e+11Hz 0.0223691 0.0777036
+ 1.302e+11Hz 0.0223959 0.0777572
+ 1.303e+11Hz 0.0224228 0.0778108
+ 1.304e+11Hz 0.0224496 0.0778643
+ 1.305e+11Hz 0.0224765 0.0779179
+ 1.306e+11Hz 0.0225033 0.0779714
+ 1.307e+11Hz 0.0225302 0.0780249
+ 1.308e+11Hz 0.0225571 0.0780783
+ 1.309e+11Hz 0.0225841 0.0781318
+ 1.31e+11Hz 0.022611 0.0781852
+ 1.311e+11Hz 0.022638 0.0782387
+ 1.312e+11Hz 0.022665 0.0782921
+ 1.313e+11Hz 0.022692 0.0783455
+ 1.314e+11Hz 0.022719 0.0783988
+ 1.315e+11Hz 0.022746 0.0784522
+ 1.316e+11Hz 0.0227731 0.0785055
+ 1.317e+11Hz 0.0228001 0.0785588
+ 1.318e+11Hz 0.0228272 0.0786121
+ 1.319e+11Hz 0.0228543 0.0786654
+ 1.32e+11Hz 0.0228815 0.0787186
+ 1.321e+11Hz 0.0229086 0.0787719
+ 1.322e+11Hz 0.0229357 0.0788251
+ 1.323e+11Hz 0.0229629 0.0788783
+ 1.324e+11Hz 0.0229901 0.0789315
+ 1.325e+11Hz 0.0230173 0.0789846
+ 1.326e+11Hz 0.0230445 0.0790378
+ 1.327e+11Hz 0.0230717 0.0790909
+ 1.328e+11Hz 0.023099 0.079144
+ 1.329e+11Hz 0.0231263 0.0791971
+ 1.33e+11Hz 0.0231535 0.0792502
+ 1.331e+11Hz 0.0231808 0.0793032
+ 1.332e+11Hz 0.0232081 0.0793562
+ 1.333e+11Hz 0.0232355 0.0794093
+ 1.334e+11Hz 0.0232628 0.0794622
+ 1.335e+11Hz 0.0232901 0.0795152
+ 1.336e+11Hz 0.0233175 0.0795682
+ 1.337e+11Hz 0.0233449 0.0796211
+ 1.338e+11Hz 0.0233723 0.079674
+ 1.339e+11Hz 0.0233997 0.0797269
+ 1.34e+11Hz 0.0234271 0.0797798
+ 1.341e+11Hz 0.0234546 0.0798326
+ 1.342e+11Hz 0.023482 0.0798855
+ 1.343e+11Hz 0.0235095 0.0799383
+ 1.344e+11Hz 0.023537 0.0799911
+ 1.345e+11Hz 0.0235645 0.0800439
+ 1.346e+11Hz 0.023592 0.0800967
+ 1.347e+11Hz 0.0236195 0.0801494
+ 1.348e+11Hz 0.023647 0.0802021
+ 1.349e+11Hz 0.0236745 0.0802548
+ 1.35e+11Hz 0.0237021 0.0803075
+ 1.351e+11Hz 0.0237297 0.0803602
+ 1.352e+11Hz 0.0237573 0.0804129
+ 1.353e+11Hz 0.0237848 0.0804655
+ 1.354e+11Hz 0.0238125 0.0805181
+ 1.355e+11Hz 0.0238401 0.0805707
+ 1.356e+11Hz 0.0238677 0.0806233
+ 1.357e+11Hz 0.0238953 0.0806759
+ 1.358e+11Hz 0.023923 0.0807284
+ 1.359e+11Hz 0.0239507 0.0807809
+ 1.36e+11Hz 0.0239783 0.0808335
+ 1.361e+11Hz 0.024006 0.0808859
+ 1.362e+11Hz 0.0240337 0.0809384
+ 1.363e+11Hz 0.0240614 0.0809909
+ 1.364e+11Hz 0.0240892 0.0810433
+ 1.365e+11Hz 0.0241169 0.0810958
+ 1.366e+11Hz 0.0241446 0.0811482
+ 1.367e+11Hz 0.0241724 0.0812006
+ 1.368e+11Hz 0.0242002 0.0812529
+ 1.369e+11Hz 0.0242279 0.0813053
+ 1.37e+11Hz 0.0242557 0.0813576
+ 1.371e+11Hz 0.0242835 0.08141
+ 1.372e+11Hz 0.0243113 0.0814623
+ 1.373e+11Hz 0.0243391 0.0815146
+ 1.374e+11Hz 0.024367 0.0815669
+ 1.375e+11Hz 0.0243948 0.0816191
+ 1.376e+11Hz 0.0244227 0.0816714
+ 1.377e+11Hz 0.0244505 0.0817236
+ 1.378e+11Hz 0.0244784 0.0817758
+ 1.379e+11Hz 0.0245063 0.081828
+ 1.38e+11Hz 0.0245342 0.0818802
+ 1.381e+11Hz 0.0245621 0.0819324
+ 1.382e+11Hz 0.02459 0.0819846
+ 1.383e+11Hz 0.0246179 0.0820367
+ 1.384e+11Hz 0.0246458 0.0820888
+ 1.385e+11Hz 0.0246738 0.082141
+ 1.386e+11Hz 0.0247017 0.0821931
+ 1.387e+11Hz 0.0247297 0.0822452
+ 1.388e+11Hz 0.0247576 0.0822972
+ 1.389e+11Hz 0.0247856 0.0823493
+ 1.39e+11Hz 0.0248136 0.0824013
+ 1.391e+11Hz 0.0248416 0.0824534
+ 1.392e+11Hz 0.0248696 0.0825054
+ 1.393e+11Hz 0.0248976 0.0825574
+ 1.394e+11Hz 0.0249257 0.0826094
+ 1.395e+11Hz 0.0249537 0.0826614
+ 1.396e+11Hz 0.0249817 0.0827134
+ 1.397e+11Hz 0.0250098 0.0827653
+ 1.398e+11Hz 0.0250379 0.0828173
+ 1.399e+11Hz 0.025066 0.0828692
+ 1.4e+11Hz 0.025094 0.0829212
+ 1.401e+11Hz 0.0251221 0.0829731
+ 1.402e+11Hz 0.0251502 0.083025
+ 1.403e+11Hz 0.0251784 0.0830769
+ 1.404e+11Hz 0.0252065 0.0831288
+ 1.405e+11Hz 0.0252346 0.0831806
+ 1.406e+11Hz 0.0252628 0.0832325
+ 1.407e+11Hz 0.0252909 0.0832844
+ 1.408e+11Hz 0.0253191 0.0833362
+ 1.409e+11Hz 0.0253473 0.0833881
+ 1.41e+11Hz 0.0253755 0.0834399
+ 1.411e+11Hz 0.0254037 0.0834917
+ 1.412e+11Hz 0.0254319 0.0835435
+ 1.413e+11Hz 0.0254601 0.0835953
+ 1.414e+11Hz 0.0254884 0.0836471
+ 1.415e+11Hz 0.0255166 0.0836989
+ 1.416e+11Hz 0.0255449 0.0837507
+ 1.417e+11Hz 0.0255732 0.0838024
+ 1.418e+11Hz 0.0256015 0.0838542
+ 1.419e+11Hz 0.0256297 0.0839059
+ 1.42e+11Hz 0.0256581 0.0839577
+ 1.421e+11Hz 0.0256864 0.0840094
+ 1.422e+11Hz 0.0257147 0.0840611
+ 1.423e+11Hz 0.0257431 0.0841129
+ 1.424e+11Hz 0.0257714 0.0841646
+ 1.425e+11Hz 0.0257998 0.0842163
+ 1.426e+11Hz 0.0258282 0.084268
+ 1.427e+11Hz 0.0258566 0.0843197
+ 1.428e+11Hz 0.025885 0.0843713
+ 1.429e+11Hz 0.0259134 0.084423
+ 1.43e+11Hz 0.0259418 0.0844747
+ 1.431e+11Hz 0.0259703 0.0845264
+ 1.432e+11Hz 0.0259988 0.084578
+ 1.433e+11Hz 0.0260273 0.0846297
+ 1.434e+11Hz 0.0260558 0.0846813
+ 1.435e+11Hz 0.0260843 0.084733
+ 1.436e+11Hz 0.0261128 0.0847846
+ 1.437e+11Hz 0.0261413 0.0848363
+ 1.438e+11Hz 0.0261699 0.0848879
+ 1.439e+11Hz 0.0261985 0.0849395
+ 1.44e+11Hz 0.0262271 0.0849911
+ 1.441e+11Hz 0.0262557 0.0850427
+ 1.442e+11Hz 0.0262843 0.0850943
+ 1.443e+11Hz 0.0263129 0.0851459
+ 1.444e+11Hz 0.0263416 0.0851975
+ 1.445e+11Hz 0.0263703 0.0852491
+ 1.446e+11Hz 0.026399 0.0853007
+ 1.447e+11Hz 0.0264277 0.0853523
+ 1.448e+11Hz 0.0264564 0.0854039
+ 1.449e+11Hz 0.0264851 0.0854555
+ 1.45e+11Hz 0.0265139 0.085507
+ 1.451e+11Hz 0.0265427 0.0855586
+ 1.452e+11Hz 0.0265715 0.0856101
+ 1.453e+11Hz 0.0266003 0.0856617
+ 1.454e+11Hz 0.0266292 0.0857133
+ 1.455e+11Hz 0.026658 0.0857648
+ 1.456e+11Hz 0.0266869 0.0858163
+ 1.457e+11Hz 0.0267158 0.0858679
+ 1.458e+11Hz 0.0267447 0.0859194
+ 1.459e+11Hz 0.0267737 0.0859709
+ 1.46e+11Hz 0.0268026 0.0860225
+ 1.461e+11Hz 0.0268316 0.086074
+ 1.462e+11Hz 0.0268606 0.0861255
+ 1.463e+11Hz 0.0268897 0.086177
+ 1.464e+11Hz 0.0269187 0.0862285
+ 1.465e+11Hz 0.0269478 0.08628
+ 1.466e+11Hz 0.0269769 0.0863315
+ 1.467e+11Hz 0.027006 0.086383
+ 1.468e+11Hz 0.0270351 0.0864345
+ 1.469e+11Hz 0.0270643 0.086486
+ 1.47e+11Hz 0.0270935 0.0865375
+ 1.471e+11Hz 0.0271227 0.0865889
+ 1.472e+11Hz 0.027152 0.0866404
+ 1.473e+11Hz 0.0271812 0.0866918
+ 1.474e+11Hz 0.0272105 0.0867433
+ 1.475e+11Hz 0.0272398 0.0867948
+ 1.476e+11Hz 0.0272692 0.0868462
+ 1.477e+11Hz 0.0272985 0.0868976
+ 1.478e+11Hz 0.0273279 0.0869491
+ 1.479e+11Hz 0.0273574 0.0870005
+ 1.48e+11Hz 0.0273868 0.0870519
+ 1.481e+11Hz 0.0274163 0.0871033
+ 1.482e+11Hz 0.0274458 0.0871547
+ 1.483e+11Hz 0.0274753 0.0872061
+ 1.484e+11Hz 0.0275049 0.0872575
+ 1.485e+11Hz 0.0275344 0.0873089
+ 1.486e+11Hz 0.0275641 0.0873603
+ 1.487e+11Hz 0.0275937 0.0874116
+ 1.488e+11Hz 0.0276234 0.087463
+ 1.489e+11Hz 0.0276531 0.0875144
+ 1.49e+11Hz 0.0276828 0.0875657
+ 1.491e+11Hz 0.0277125 0.087617
+ 1.492e+11Hz 0.0277423 0.0876684
+ 1.493e+11Hz 0.0277721 0.0877197
+ 1.494e+11Hz 0.027802 0.087771
+ 1.495e+11Hz 0.0278319 0.0878223
+ 1.496e+11Hz 0.0278618 0.0878736
+ 1.497e+11Hz 0.0278917 0.0879249
+ 1.498e+11Hz 0.0279217 0.0879761
+ 1.499e+11Hz 0.0279517 0.0880274
+ 1.5e+11Hz 0.0279817 0.0880786
+ ]

A12 %vd(20 3) %vd(12, 3) xfer2
.model xfer2 xfer R_I=true table=[
+ 0Hz 0.997077 0
+ 1e+08Hz 0.997077 -0.0002216
+ 2e+08Hz 0.997076 -0.000443198
+ 3e+08Hz 0.997076 -0.000664791
+ 4e+08Hz 0.997076 -0.000886377
+ 5e+08Hz 0.997075 -0.00110795
+ 6e+08Hz 0.997074 -0.00132952
+ 7e+08Hz 0.997073 -0.00155107
+ 8e+08Hz 0.997072 -0.0017726
+ 9e+08Hz 0.99707 -0.00199412
+ 1e+09Hz 0.997069 -0.00221561
+ 1.1e+09Hz 0.997067 -0.00243708
+ 1.2e+09Hz 0.997066 -0.00265853
+ 1.3e+09Hz 0.997063 -0.00287994
+ 1.4e+09Hz 0.997061 -0.00310133
+ 1.5e+09Hz 0.997059 -0.00332268
+ 1.6e+09Hz 0.997057 -0.003544
+ 1.7e+09Hz 0.997054 -0.00376528
+ 1.8e+09Hz 0.997051 -0.00398652
+ 1.9e+09Hz 0.997049 -0.00420772
+ 2e+09Hz 0.997046 -0.00442888
+ 2.1e+09Hz 0.997043 -0.00464999
+ 2.2e+09Hz 0.997039 -0.00487106
+ 2.3e+09Hz 0.997036 -0.00509207
+ 2.4e+09Hz 0.997032 -0.00531304
+ 2.5e+09Hz 0.997028 -0.00553395
+ 2.6e+09Hz 0.997025 -0.0057548
+ 2.7e+09Hz 0.99702 -0.00597559
+ 2.8e+09Hz 0.997016 -0.00619633
+ 2.9e+09Hz 0.997012 -0.006417
+ 3e+09Hz 0.997008 -0.00663762
+ 3.1e+09Hz 0.997003 -0.00685816
+ 3.2e+09Hz 0.996998 -0.00707864
+ 3.3e+09Hz 0.996994 -0.00729905
+ 3.4e+09Hz 0.996989 -0.0075194
+ 3.5e+09Hz 0.996984 -0.00773967
+ 3.6e+09Hz 0.996978 -0.00795986
+ 3.7e+09Hz 0.996973 -0.00817999
+ 3.8e+09Hz 0.996968 -0.00840003
+ 3.9e+09Hz 0.996962 -0.00862
+ 4e+09Hz 0.996956 -0.00883989
+ 4.1e+09Hz 0.99695 -0.0090597
+ 4.2e+09Hz 0.996944 -0.00927942
+ 4.3e+09Hz 0.996938 -0.00949907
+ 4.4e+09Hz 0.996932 -0.00971862
+ 4.5e+09Hz 0.996926 -0.0099381
+ 4.6e+09Hz 0.996919 -0.0101575
+ 4.7e+09Hz 0.996913 -0.0103768
+ 4.8e+09Hz 0.996906 -0.010596
+ 4.9e+09Hz 0.9969 -0.0108151
+ 5e+09Hz 0.996893 -0.0110341
+ 5.1e+09Hz 0.996886 -0.0112531
+ 5.2e+09Hz 0.996879 -0.0114719
+ 5.3e+09Hz 0.996872 -0.0116907
+ 5.4e+09Hz 0.996864 -0.0119093
+ 5.5e+09Hz 0.996857 -0.0121279
+ 5.6e+09Hz 0.99685 -0.0123464
+ 5.7e+09Hz 0.996842 -0.0125647
+ 5.8e+09Hz 0.996834 -0.012783
+ 5.9e+09Hz 0.996827 -0.0130012
+ 6e+09Hz 0.996819 -0.0132193
+ 6.1e+09Hz 0.996811 -0.0134373
+ 6.2e+09Hz 0.996803 -0.0136551
+ 6.3e+09Hz 0.996795 -0.0138729
+ 6.4e+09Hz 0.996787 -0.0140906
+ 6.5e+09Hz 0.996779 -0.0143082
+ 6.6e+09Hz 0.99677 -0.0145257
+ 6.7e+09Hz 0.996762 -0.0147431
+ 6.8e+09Hz 0.996754 -0.0149604
+ 6.9e+09Hz 0.996745 -0.0151776
+ 7e+09Hz 0.996737 -0.0153947
+ 7.1e+09Hz 0.996728 -0.0156117
+ 7.2e+09Hz 0.996719 -0.0158286
+ 7.3e+09Hz 0.996711 -0.0160453
+ 7.4e+09Hz 0.996702 -0.0162621
+ 7.5e+09Hz 0.996693 -0.0164787
+ 7.6e+09Hz 0.996684 -0.0166951
+ 7.7e+09Hz 0.996675 -0.0169116
+ 7.8e+09Hz 0.996666 -0.0171279
+ 7.9e+09Hz 0.996657 -0.0173441
+ 8e+09Hz 0.996648 -0.0175602
+ 8.1e+09Hz 0.996639 -0.0177762
+ 8.2e+09Hz 0.996629 -0.0179921
+ 8.3e+09Hz 0.99662 -0.0182079
+ 8.4e+09Hz 0.996611 -0.0184236
+ 8.5e+09Hz 0.996601 -0.0186393
+ 8.6e+09Hz 0.996592 -0.0188548
+ 8.7e+09Hz 0.996583 -0.0190703
+ 8.8e+09Hz 0.996573 -0.0192856
+ 8.9e+09Hz 0.996564 -0.0195009
+ 9e+09Hz 0.996554 -0.0197161
+ 9.1e+09Hz 0.996545 -0.0199312
+ 9.2e+09Hz 0.996535 -0.0201462
+ 9.3e+09Hz 0.996525 -0.0203611
+ 9.4e+09Hz 0.996515 -0.0205759
+ 9.5e+09Hz 0.996506 -0.0207906
+ 9.6e+09Hz 0.996496 -0.0210053
+ 9.7e+09Hz 0.996486 -0.0212198
+ 9.8e+09Hz 0.996476 -0.0214343
+ 9.9e+09Hz 0.996467 -0.0216487
+ 1e+10Hz 0.996457 -0.021863
+ 1.01e+10Hz 0.996447 -0.0220773
+ 1.02e+10Hz 0.996437 -0.0222915
+ 1.03e+10Hz 0.996427 -0.0225055
+ 1.04e+10Hz 0.996417 -0.0227196
+ 1.05e+10Hz 0.996407 -0.0229335
+ 1.06e+10Hz 0.996398 -0.0231473
+ 1.07e+10Hz 0.996387 -0.0233611
+ 1.08e+10Hz 0.996378 -0.0235749
+ 1.09e+10Hz 0.996367 -0.0237885
+ 1.1e+10Hz 0.996358 -0.0240021
+ 1.11e+10Hz 0.996348 -0.0242156
+ 1.12e+10Hz 0.996337 -0.024429
+ 1.13e+10Hz 0.996327 -0.0246424
+ 1.14e+10Hz 0.996317 -0.0248557
+ 1.15e+10Hz 0.996307 -0.025069
+ 1.16e+10Hz 0.996297 -0.0252821
+ 1.17e+10Hz 0.996287 -0.0254953
+ 1.18e+10Hz 0.996277 -0.0257084
+ 1.19e+10Hz 0.996267 -0.0259214
+ 1.2e+10Hz 0.996257 -0.0261343
+ 1.21e+10Hz 0.996247 -0.0263472
+ 1.22e+10Hz 0.996237 -0.0265601
+ 1.23e+10Hz 0.996227 -0.0267729
+ 1.24e+10Hz 0.996216 -0.0269856
+ 1.25e+10Hz 0.996206 -0.0271983
+ 1.26e+10Hz 0.996196 -0.0274109
+ 1.27e+10Hz 0.996186 -0.0276235
+ 1.28e+10Hz 0.996176 -0.0278361
+ 1.29e+10Hz 0.996166 -0.0280486
+ 1.3e+10Hz 0.996155 -0.0282611
+ 1.31e+10Hz 0.996145 -0.0284735
+ 1.32e+10Hz 0.996135 -0.0286859
+ 1.33e+10Hz 0.996125 -0.0288982
+ 1.34e+10Hz 0.996115 -0.0291105
+ 1.35e+10Hz 0.996105 -0.0293228
+ 1.36e+10Hz 0.996094 -0.029535
+ 1.37e+10Hz 0.996084 -0.0297472
+ 1.38e+10Hz 0.996074 -0.0299594
+ 1.39e+10Hz 0.996064 -0.0301715
+ 1.4e+10Hz 0.996054 -0.0303836
+ 1.41e+10Hz 0.996043 -0.0305957
+ 1.42e+10Hz 0.996033 -0.0308077
+ 1.43e+10Hz 0.996023 -0.0310197
+ 1.44e+10Hz 0.996013 -0.0312317
+ 1.45e+10Hz 0.996003 -0.0314437
+ 1.46e+10Hz 0.995992 -0.0316557
+ 1.47e+10Hz 0.995982 -0.0318676
+ 1.48e+10Hz 0.995972 -0.0320795
+ 1.49e+10Hz 0.995962 -0.0322914
+ 1.5e+10Hz 0.995951 -0.0325032
+ 1.51e+10Hz 0.995941 -0.0327151
+ 1.52e+10Hz 0.995931 -0.0329269
+ 1.53e+10Hz 0.99592 -0.0331387
+ 1.54e+10Hz 0.99591 -0.0333505
+ 1.55e+10Hz 0.9959 -0.0335623
+ 1.56e+10Hz 0.995889 -0.033774
+ 1.57e+10Hz 0.995879 -0.0339858
+ 1.58e+10Hz 0.995869 -0.0341975
+ 1.59e+10Hz 0.995858 -0.0344093
+ 1.6e+10Hz 0.995848 -0.034621
+ 1.61e+10Hz 0.995838 -0.0348327
+ 1.62e+10Hz 0.995827 -0.0350444
+ 1.63e+10Hz 0.995817 -0.0352561
+ 1.64e+10Hz 0.995806 -0.0354678
+ 1.65e+10Hz 0.995796 -0.0356795
+ 1.66e+10Hz 0.995785 -0.0358912
+ 1.67e+10Hz 0.995775 -0.0361029
+ 1.68e+10Hz 0.995765 -0.0363146
+ 1.69e+10Hz 0.995754 -0.0365263
+ 1.7e+10Hz 0.995744 -0.0367379
+ 1.71e+10Hz 0.995733 -0.0369496
+ 1.72e+10Hz 0.995722 -0.0371613
+ 1.73e+10Hz 0.995712 -0.037373
+ 1.74e+10Hz 0.995701 -0.0375846
+ 1.75e+10Hz 0.995691 -0.0377963
+ 1.76e+10Hz 0.99568 -0.038008
+ 1.77e+10Hz 0.995669 -0.0382197
+ 1.78e+10Hz 0.995659 -0.0384314
+ 1.79e+10Hz 0.995648 -0.0386431
+ 1.8e+10Hz 0.995637 -0.0388548
+ 1.81e+10Hz 0.995626 -0.0390665
+ 1.82e+10Hz 0.995616 -0.0392782
+ 1.83e+10Hz 0.995605 -0.0394899
+ 1.84e+10Hz 0.995594 -0.0397016
+ 1.85e+10Hz 0.995583 -0.0399133
+ 1.86e+10Hz 0.995572 -0.0401251
+ 1.87e+10Hz 0.995561 -0.0403368
+ 1.88e+10Hz 0.99555 -0.0405485
+ 1.89e+10Hz 0.995539 -0.0407603
+ 1.9e+10Hz 0.995528 -0.0409721
+ 1.91e+10Hz 0.995517 -0.0411838
+ 1.92e+10Hz 0.995506 -0.0413956
+ 1.93e+10Hz 0.995495 -0.0416074
+ 1.94e+10Hz 0.995484 -0.0418192
+ 1.95e+10Hz 0.995472 -0.042031
+ 1.96e+10Hz 0.995461 -0.0422428
+ 1.97e+10Hz 0.99545 -0.0424546
+ 1.98e+10Hz 0.995439 -0.0426664
+ 1.99e+10Hz 0.995427 -0.0428783
+ 2e+10Hz 0.995416 -0.0430901
+ 2.01e+10Hz 0.995404 -0.043302
+ 2.02e+10Hz 0.995393 -0.0435139
+ 2.03e+10Hz 0.995382 -0.0437257
+ 2.04e+10Hz 0.99537 -0.0439376
+ 2.05e+10Hz 0.995358 -0.0441495
+ 2.06e+10Hz 0.995347 -0.0443614
+ 2.07e+10Hz 0.995335 -0.0445733
+ 2.08e+10Hz 0.995323 -0.0447853
+ 2.09e+10Hz 0.995311 -0.0449972
+ 2.1e+10Hz 0.9953 -0.0452091
+ 2.11e+10Hz 0.995288 -0.0454211
+ 2.12e+10Hz 0.995276 -0.0456331
+ 2.13e+10Hz 0.995264 -0.045845
+ 2.14e+10Hz 0.995252 -0.046057
+ 2.15e+10Hz 0.99524 -0.046269
+ 2.16e+10Hz 0.995228 -0.046481
+ 2.17e+10Hz 0.995216 -0.046693
+ 2.18e+10Hz 0.995203 -0.046905
+ 2.19e+10Hz 0.995191 -0.0471171
+ 2.2e+10Hz 0.995179 -0.0473291
+ 2.21e+10Hz 0.995166 -0.0475411
+ 2.22e+10Hz 0.995154 -0.0477532
+ 2.23e+10Hz 0.995142 -0.0479652
+ 2.24e+10Hz 0.995129 -0.0481773
+ 2.25e+10Hz 0.995116 -0.0483893
+ 2.26e+10Hz 0.995104 -0.0486014
+ 2.27e+10Hz 0.995091 -0.0488135
+ 2.28e+10Hz 0.995078 -0.0490256
+ 2.29e+10Hz 0.995066 -0.0492377
+ 2.3e+10Hz 0.995053 -0.0494498
+ 2.31e+10Hz 0.99504 -0.0496619
+ 2.32e+10Hz 0.995027 -0.049874
+ 2.33e+10Hz 0.995014 -0.0500861
+ 2.34e+10Hz 0.995001 -0.0502982
+ 2.35e+10Hz 0.994988 -0.0505103
+ 2.36e+10Hz 0.994975 -0.0507225
+ 2.37e+10Hz 0.994962 -0.0509346
+ 2.38e+10Hz 0.994948 -0.0511467
+ 2.39e+10Hz 0.994935 -0.0513588
+ 2.4e+10Hz 0.994922 -0.051571
+ 2.41e+10Hz 0.994908 -0.0517831
+ 2.42e+10Hz 0.994895 -0.0519952
+ 2.43e+10Hz 0.994881 -0.0522074
+ 2.44e+10Hz 0.994867 -0.0524195
+ 2.45e+10Hz 0.994854 -0.0526316
+ 2.46e+10Hz 0.99484 -0.0528438
+ 2.47e+10Hz 0.994826 -0.0530559
+ 2.48e+10Hz 0.994812 -0.053268
+ 2.49e+10Hz 0.994798 -0.0534802
+ 2.5e+10Hz 0.994784 -0.0536923
+ 2.51e+10Hz 0.99477 -0.0539044
+ 2.52e+10Hz 0.994756 -0.0541166
+ 2.53e+10Hz 0.994742 -0.0543287
+ 2.54e+10Hz 0.994728 -0.0545408
+ 2.55e+10Hz 0.994714 -0.0547529
+ 2.56e+10Hz 0.994699 -0.054965
+ 2.57e+10Hz 0.994685 -0.0551772
+ 2.58e+10Hz 0.99467 -0.0553893
+ 2.59e+10Hz 0.994656 -0.0556014
+ 2.6e+10Hz 0.994641 -0.0558135
+ 2.61e+10Hz 0.994627 -0.0560256
+ 2.62e+10Hz 0.994612 -0.0562376
+ 2.63e+10Hz 0.994597 -0.0564497
+ 2.64e+10Hz 0.994583 -0.0566618
+ 2.65e+10Hz 0.994568 -0.0568738
+ 2.66e+10Hz 0.994553 -0.0570859
+ 2.67e+10Hz 0.994538 -0.057298
+ 2.68e+10Hz 0.994523 -0.05751
+ 2.69e+10Hz 0.994508 -0.057722
+ 2.7e+10Hz 0.994493 -0.0579341
+ 2.71e+10Hz 0.994477 -0.0581461
+ 2.72e+10Hz 0.994462 -0.0583581
+ 2.73e+10Hz 0.994447 -0.0585701
+ 2.74e+10Hz 0.994431 -0.0587821
+ 2.75e+10Hz 0.994416 -0.058994
+ 2.76e+10Hz 0.994401 -0.059206
+ 2.77e+10Hz 0.994385 -0.059418
+ 2.78e+10Hz 0.994369 -0.0596299
+ 2.79e+10Hz 0.994354 -0.0598419
+ 2.8e+10Hz 0.994338 -0.0600538
+ 2.81e+10Hz 0.994322 -0.0602657
+ 2.82e+10Hz 0.994306 -0.0604776
+ 2.83e+10Hz 0.994291 -0.0606895
+ 2.84e+10Hz 0.994275 -0.0609014
+ 2.85e+10Hz 0.994259 -0.0611132
+ 2.86e+10Hz 0.994243 -0.0613251
+ 2.87e+10Hz 0.994227 -0.0615369
+ 2.88e+10Hz 0.99421 -0.0617487
+ 2.89e+10Hz 0.994194 -0.0619606
+ 2.9e+10Hz 0.994178 -0.0621724
+ 2.91e+10Hz 0.994162 -0.0623841
+ 2.92e+10Hz 0.994145 -0.0625959
+ 2.93e+10Hz 0.994129 -0.0628077
+ 2.94e+10Hz 0.994112 -0.0630194
+ 2.95e+10Hz 0.994096 -0.0632311
+ 2.96e+10Hz 0.994079 -0.0634429
+ 2.97e+10Hz 0.994063 -0.0636546
+ 2.98e+10Hz 0.994046 -0.0638663
+ 2.99e+10Hz 0.994029 -0.0640779
+ 3e+10Hz 0.994013 -0.0642896
+ 3.01e+10Hz 0.993996 -0.0645012
+ 3.02e+10Hz 0.993979 -0.0647129
+ 3.03e+10Hz 0.993962 -0.0649245
+ 3.04e+10Hz 0.993945 -0.0651361
+ 3.05e+10Hz 0.993928 -0.0653477
+ 3.06e+10Hz 0.993911 -0.0655592
+ 3.07e+10Hz 0.993894 -0.0657708
+ 3.08e+10Hz 0.993877 -0.0659823
+ 3.09e+10Hz 0.993859 -0.0661938
+ 3.1e+10Hz 0.993842 -0.0664054
+ 3.11e+10Hz 0.993825 -0.0666169
+ 3.12e+10Hz 0.993807 -0.0668283
+ 3.13e+10Hz 0.99379 -0.0670398
+ 3.14e+10Hz 0.993773 -0.0672512
+ 3.15e+10Hz 0.993755 -0.0674627
+ 3.16e+10Hz 0.993738 -0.0676741
+ 3.17e+10Hz 0.99372 -0.0678855
+ 3.18e+10Hz 0.993703 -0.0680969
+ 3.19e+10Hz 0.993685 -0.0683083
+ 3.2e+10Hz 0.993667 -0.0685196
+ 3.21e+10Hz 0.993649 -0.0687309
+ 3.22e+10Hz 0.993632 -0.0689423
+ 3.23e+10Hz 0.993614 -0.0691536
+ 3.24e+10Hz 0.993596 -0.0693649
+ 3.25e+10Hz 0.993578 -0.0695762
+ 3.26e+10Hz 0.99356 -0.0697874
+ 3.27e+10Hz 0.993542 -0.0699987
+ 3.28e+10Hz 0.993524 -0.0702099
+ 3.29e+10Hz 0.993506 -0.0704212
+ 3.3e+10Hz 0.993488 -0.0706324
+ 3.31e+10Hz 0.99347 -0.0708436
+ 3.32e+10Hz 0.993451 -0.0710547
+ 3.33e+10Hz 0.993433 -0.0712659
+ 3.34e+10Hz 0.993415 -0.0714771
+ 3.35e+10Hz 0.993397 -0.0716882
+ 3.36e+10Hz 0.993378 -0.0718994
+ 3.37e+10Hz 0.99336 -0.0721105
+ 3.38e+10Hz 0.993341 -0.0723216
+ 3.39e+10Hz 0.993323 -0.0725327
+ 3.4e+10Hz 0.993304 -0.0727437
+ 3.41e+10Hz 0.993286 -0.0729548
+ 3.42e+10Hz 0.993267 -0.0731659
+ 3.43e+10Hz 0.993248 -0.0733769
+ 3.44e+10Hz 0.99323 -0.0735879
+ 3.45e+10Hz 0.993211 -0.073799
+ 3.46e+10Hz 0.993192 -0.07401
+ 3.47e+10Hz 0.993174 -0.074221
+ 3.48e+10Hz 0.993155 -0.074432
+ 3.49e+10Hz 0.993136 -0.0746429
+ 3.5e+10Hz 0.993117 -0.0748539
+ 3.51e+10Hz 0.993098 -0.0750649
+ 3.52e+10Hz 0.993079 -0.0752758
+ 3.53e+10Hz 0.99306 -0.0754867
+ 3.54e+10Hz 0.993041 -0.0756977
+ 3.55e+10Hz 0.993022 -0.0759086
+ 3.56e+10Hz 0.993003 -0.0761195
+ 3.57e+10Hz 0.992984 -0.0763304
+ 3.58e+10Hz 0.992964 -0.0765413
+ 3.59e+10Hz 0.992945 -0.0767522
+ 3.6e+10Hz 0.992926 -0.076963
+ 3.61e+10Hz 0.992907 -0.0771739
+ 3.62e+10Hz 0.992887 -0.0773848
+ 3.63e+10Hz 0.992868 -0.0775956
+ 3.64e+10Hz 0.992848 -0.0778064
+ 3.65e+10Hz 0.992829 -0.0780173
+ 3.66e+10Hz 0.99281 -0.0782281
+ 3.67e+10Hz 0.99279 -0.0784389
+ 3.68e+10Hz 0.99277 -0.0786497
+ 3.69e+10Hz 0.992751 -0.0788605
+ 3.7e+10Hz 0.992731 -0.0790713
+ 3.71e+10Hz 0.992712 -0.0792821
+ 3.72e+10Hz 0.992692 -0.0794929
+ 3.73e+10Hz 0.992672 -0.0797037
+ 3.74e+10Hz 0.992652 -0.0799145
+ 3.75e+10Hz 0.992633 -0.0801253
+ 3.76e+10Hz 0.992613 -0.080336
+ 3.77e+10Hz 0.992593 -0.0805468
+ 3.78e+10Hz 0.992573 -0.0807576
+ 3.79e+10Hz 0.992553 -0.0809683
+ 3.8e+10Hz 0.992533 -0.0811791
+ 3.81e+10Hz 0.992513 -0.0813898
+ 3.82e+10Hz 0.992493 -0.0816006
+ 3.83e+10Hz 0.992473 -0.0818113
+ 3.84e+10Hz 0.992453 -0.082022
+ 3.85e+10Hz 0.992433 -0.0822328
+ 3.86e+10Hz 0.992413 -0.0824435
+ 3.87e+10Hz 0.992392 -0.0826543
+ 3.88e+10Hz 0.992372 -0.082865
+ 3.89e+10Hz 0.992352 -0.0830757
+ 3.9e+10Hz 0.992332 -0.0832864
+ 3.91e+10Hz 0.992311 -0.0834972
+ 3.92e+10Hz 0.992291 -0.0837079
+ 3.93e+10Hz 0.99227 -0.0839186
+ 3.94e+10Hz 0.99225 -0.0841293
+ 3.95e+10Hz 0.992229 -0.0843401
+ 3.96e+10Hz 0.992209 -0.0845508
+ 3.97e+10Hz 0.992188 -0.0847615
+ 3.98e+10Hz 0.992168 -0.0849722
+ 3.99e+10Hz 0.992147 -0.0851829
+ 4e+10Hz 0.992126 -0.0853937
+ 4.01e+10Hz 0.992106 -0.0856044
+ 4.02e+10Hz 0.992085 -0.0858151
+ 4.03e+10Hz 0.992064 -0.0860258
+ 4.04e+10Hz 0.992043 -0.0862365
+ 4.05e+10Hz 0.992022 -0.0864473
+ 4.06e+10Hz 0.992001 -0.086658
+ 4.07e+10Hz 0.991981 -0.0868687
+ 4.08e+10Hz 0.99196 -0.0870794
+ 4.09e+10Hz 0.991938 -0.0872901
+ 4.1e+10Hz 0.991918 -0.0875009
+ 4.11e+10Hz 0.991896 -0.0877116
+ 4.12e+10Hz 0.991875 -0.0879223
+ 4.13e+10Hz 0.991854 -0.0881331
+ 4.14e+10Hz 0.991833 -0.0883438
+ 4.15e+10Hz 0.991812 -0.0885545
+ 4.16e+10Hz 0.99179 -0.0887653
+ 4.17e+10Hz 0.991769 -0.088976
+ 4.18e+10Hz 0.991748 -0.0891867
+ 4.19e+10Hz 0.991726 -0.0893975
+ 4.2e+10Hz 0.991705 -0.0896082
+ 4.21e+10Hz 0.991683 -0.089819
+ 4.22e+10Hz 0.991662 -0.0900297
+ 4.23e+10Hz 0.99164 -0.0902405
+ 4.24e+10Hz 0.991619 -0.0904512
+ 4.25e+10Hz 0.991597 -0.090662
+ 4.26e+10Hz 0.991575 -0.0908727
+ 4.27e+10Hz 0.991553 -0.0910835
+ 4.28e+10Hz 0.991532 -0.0912942
+ 4.29e+10Hz 0.99151 -0.091505
+ 4.3e+10Hz 0.991488 -0.0917158
+ 4.31e+10Hz 0.991466 -0.0919265
+ 4.32e+10Hz 0.991444 -0.0921373
+ 4.33e+10Hz 0.991422 -0.0923481
+ 4.34e+10Hz 0.9914 -0.0925589
+ 4.35e+10Hz 0.991378 -0.0927696
+ 4.36e+10Hz 0.991356 -0.0929804
+ 4.37e+10Hz 0.991334 -0.0931912
+ 4.38e+10Hz 0.991312 -0.093402
+ 4.39e+10Hz 0.99129 -0.0936128
+ 4.4e+10Hz 0.991267 -0.0938236
+ 4.41e+10Hz 0.991245 -0.0940344
+ 4.42e+10Hz 0.991223 -0.0942451
+ 4.43e+10Hz 0.9912 -0.0944559
+ 4.44e+10Hz 0.991178 -0.0946667
+ 4.45e+10Hz 0.991155 -0.0948776
+ 4.46e+10Hz 0.991132 -0.0950884
+ 4.47e+10Hz 0.99111 -0.0952991
+ 4.48e+10Hz 0.991087 -0.09551
+ 4.49e+10Hz 0.991065 -0.0957208
+ 4.5e+10Hz 0.991042 -0.0959316
+ 4.51e+10Hz 0.991019 -0.0961424
+ 4.52e+10Hz 0.990996 -0.0963532
+ 4.53e+10Hz 0.990973 -0.096564
+ 4.54e+10Hz 0.99095 -0.0967748
+ 4.55e+10Hz 0.990927 -0.0969856
+ 4.56e+10Hz 0.990904 -0.0971964
+ 4.57e+10Hz 0.990881 -0.0974073
+ 4.58e+10Hz 0.990858 -0.0976181
+ 4.59e+10Hz 0.990835 -0.0978289
+ 4.6e+10Hz 0.990812 -0.0980397
+ 4.61e+10Hz 0.990789 -0.0982505
+ 4.62e+10Hz 0.990765 -0.0984613
+ 4.63e+10Hz 0.990742 -0.0986722
+ 4.64e+10Hz 0.990719 -0.098883
+ 4.65e+10Hz 0.990695 -0.0990938
+ 4.66e+10Hz 0.990672 -0.0993046
+ 4.67e+10Hz 0.990648 -0.0995154
+ 4.68e+10Hz 0.990625 -0.0997263
+ 4.69e+10Hz 0.990601 -0.0999371
+ 4.7e+10Hz 0.990577 -0.100148
+ 4.71e+10Hz 0.990554 -0.100359
+ 4.72e+10Hz 0.99053 -0.10057
+ 4.73e+10Hz 0.990506 -0.10078
+ 4.74e+10Hz 0.990482 -0.100991
+ 4.75e+10Hz 0.990458 -0.101202
+ 4.76e+10Hz 0.990434 -0.101413
+ 4.77e+10Hz 0.99041 -0.101624
+ 4.78e+10Hz 0.990386 -0.101834
+ 4.79e+10Hz 0.990362 -0.102045
+ 4.8e+10Hz 0.990338 -0.102256
+ 4.81e+10Hz 0.990314 -0.102467
+ 4.82e+10Hz 0.99029 -0.102678
+ 4.83e+10Hz 0.990265 -0.102888
+ 4.84e+10Hz 0.990241 -0.103099
+ 4.85e+10Hz 0.990216 -0.10331
+ 4.86e+10Hz 0.990192 -0.103521
+ 4.87e+10Hz 0.990167 -0.103731
+ 4.88e+10Hz 0.990143 -0.103942
+ 4.89e+10Hz 0.990118 -0.104153
+ 4.9e+10Hz 0.990094 -0.104364
+ 4.91e+10Hz 0.990069 -0.104574
+ 4.92e+10Hz 0.990044 -0.104785
+ 4.93e+10Hz 0.990019 -0.104996
+ 4.94e+10Hz 0.989994 -0.105207
+ 4.95e+10Hz 0.989969 -0.105417
+ 4.96e+10Hz 0.989945 -0.105628
+ 4.97e+10Hz 0.989919 -0.105839
+ 4.98e+10Hz 0.989894 -0.10605
+ 4.99e+10Hz 0.989869 -0.10626
+ 5e+10Hz 0.989844 -0.106471
+ 5.01e+10Hz 0.989819 -0.106682
+ 5.02e+10Hz 0.989794 -0.106892
+ 5.03e+10Hz 0.989768 -0.107103
+ 5.04e+10Hz 0.989743 -0.107314
+ 5.05e+10Hz 0.989718 -0.107524
+ 5.06e+10Hz 0.989692 -0.107735
+ 5.07e+10Hz 0.989667 -0.107946
+ 5.08e+10Hz 0.989641 -0.108156
+ 5.09e+10Hz 0.989615 -0.108367
+ 5.1e+10Hz 0.98959 -0.108578
+ 5.11e+10Hz 0.989564 -0.108788
+ 5.12e+10Hz 0.989538 -0.108999
+ 5.13e+10Hz 0.989512 -0.10921
+ 5.14e+10Hz 0.989487 -0.10942
+ 5.15e+10Hz 0.989461 -0.109631
+ 5.16e+10Hz 0.989435 -0.109841
+ 5.17e+10Hz 0.989409 -0.110052
+ 5.18e+10Hz 0.989383 -0.110262
+ 5.19e+10Hz 0.989356 -0.110473
+ 5.2e+10Hz 0.98933 -0.110683
+ 5.21e+10Hz 0.989304 -0.110894
+ 5.22e+10Hz 0.989278 -0.111104
+ 5.23e+10Hz 0.989251 -0.111315
+ 5.24e+10Hz 0.989225 -0.111525
+ 5.25e+10Hz 0.989199 -0.111736
+ 5.26e+10Hz 0.989172 -0.111947
+ 5.27e+10Hz 0.989146 -0.112157
+ 5.28e+10Hz 0.989119 -0.112367
+ 5.29e+10Hz 0.989093 -0.112578
+ 5.3e+10Hz 0.989066 -0.112788
+ 5.31e+10Hz 0.989039 -0.112999
+ 5.32e+10Hz 0.989012 -0.113209
+ 5.33e+10Hz 0.988986 -0.11342
+ 5.34e+10Hz 0.988959 -0.11363
+ 5.35e+10Hz 0.988932 -0.11384
+ 5.36e+10Hz 0.988905 -0.114051
+ 5.37e+10Hz 0.988878 -0.114261
+ 5.38e+10Hz 0.988851 -0.114471
+ 5.39e+10Hz 0.988824 -0.114682
+ 5.4e+10Hz 0.988797 -0.114892
+ 5.41e+10Hz 0.98877 -0.115102
+ 5.42e+10Hz 0.988742 -0.115313
+ 5.43e+10Hz 0.988715 -0.115523
+ 5.44e+10Hz 0.988688 -0.115733
+ 5.45e+10Hz 0.98866 -0.115943
+ 5.46e+10Hz 0.988633 -0.116154
+ 5.47e+10Hz 0.988606 -0.116364
+ 5.48e+10Hz 0.988578 -0.116574
+ 5.49e+10Hz 0.98855 -0.116784
+ 5.5e+10Hz 0.988523 -0.116994
+ 5.51e+10Hz 0.988495 -0.117205
+ 5.52e+10Hz 0.988468 -0.117415
+ 5.53e+10Hz 0.98844 -0.117625
+ 5.54e+10Hz 0.988412 -0.117835
+ 5.55e+10Hz 0.988384 -0.118045
+ 5.56e+10Hz 0.988356 -0.118255
+ 5.57e+10Hz 0.988328 -0.118465
+ 5.58e+10Hz 0.9883 -0.118676
+ 5.59e+10Hz 0.988272 -0.118886
+ 5.6e+10Hz 0.988244 -0.119096
+ 5.61e+10Hz 0.988216 -0.119306
+ 5.62e+10Hz 0.988188 -0.119516
+ 5.63e+10Hz 0.98816 -0.119726
+ 5.64e+10Hz 0.988132 -0.119936
+ 5.65e+10Hz 0.988103 -0.120146
+ 5.66e+10Hz 0.988075 -0.120356
+ 5.67e+10Hz 0.988047 -0.120566
+ 5.68e+10Hz 0.988018 -0.120776
+ 5.69e+10Hz 0.98799 -0.120985
+ 5.7e+10Hz 0.987961 -0.121195
+ 5.71e+10Hz 0.987933 -0.121405
+ 5.72e+10Hz 0.987904 -0.121615
+ 5.73e+10Hz 0.987876 -0.121825
+ 5.74e+10Hz 0.987847 -0.122035
+ 5.75e+10Hz 0.987818 -0.122245
+ 5.76e+10Hz 0.987789 -0.122455
+ 5.77e+10Hz 0.987761 -0.122664
+ 5.78e+10Hz 0.987732 -0.122874
+ 5.79e+10Hz 0.987703 -0.123084
+ 5.8e+10Hz 0.987674 -0.123294
+ 5.81e+10Hz 0.987645 -0.123504
+ 5.82e+10Hz 0.987616 -0.123714
+ 5.83e+10Hz 0.987587 -0.123923
+ 5.84e+10Hz 0.987558 -0.124133
+ 5.85e+10Hz 0.987529 -0.124343
+ 5.86e+10Hz 0.987499 -0.124552
+ 5.87e+10Hz 0.98747 -0.124762
+ 5.88e+10Hz 0.987441 -0.124972
+ 5.89e+10Hz 0.987412 -0.125181
+ 5.9e+10Hz 0.987382 -0.125391
+ 5.91e+10Hz 0.987353 -0.125601
+ 5.92e+10Hz 0.987324 -0.12581
+ 5.93e+10Hz 0.987294 -0.12602
+ 5.94e+10Hz 0.987264 -0.12623
+ 5.95e+10Hz 0.987235 -0.126439
+ 5.96e+10Hz 0.987205 -0.126649
+ 5.97e+10Hz 0.987176 -0.126858
+ 5.98e+10Hz 0.987146 -0.127068
+ 5.99e+10Hz 0.987116 -0.127277
+ 6e+10Hz 0.987086 -0.127487
+ 6.01e+10Hz 0.987057 -0.127697
+ 6.02e+10Hz 0.987027 -0.127906
+ 6.03e+10Hz 0.986997 -0.128116
+ 6.04e+10Hz 0.986967 -0.128325
+ 6.05e+10Hz 0.986937 -0.128534
+ 6.06e+10Hz 0.986907 -0.128744
+ 6.07e+10Hz 0.986877 -0.128953
+ 6.08e+10Hz 0.986847 -0.129163
+ 6.09e+10Hz 0.986817 -0.129372
+ 6.1e+10Hz 0.986787 -0.129582
+ 6.11e+10Hz 0.986756 -0.129791
+ 6.12e+10Hz 0.986726 -0.130001
+ 6.13e+10Hz 0.986696 -0.13021
+ 6.14e+10Hz 0.986665 -0.130419
+ 6.15e+10Hz 0.986635 -0.130629
+ 6.16e+10Hz 0.986605 -0.130838
+ 6.17e+10Hz 0.986574 -0.131048
+ 6.18e+10Hz 0.986544 -0.131257
+ 6.19e+10Hz 0.986513 -0.131466
+ 6.2e+10Hz 0.986483 -0.131676
+ 6.21e+10Hz 0.986452 -0.131885
+ 6.22e+10Hz 0.986421 -0.132094
+ 6.23e+10Hz 0.986391 -0.132303
+ 6.24e+10Hz 0.98636 -0.132513
+ 6.25e+10Hz 0.986329 -0.132722
+ 6.26e+10Hz 0.986298 -0.132931
+ 6.27e+10Hz 0.986267 -0.13314
+ 6.28e+10Hz 0.986237 -0.13335
+ 6.29e+10Hz 0.986206 -0.133559
+ 6.3e+10Hz 0.986175 -0.133768
+ 6.31e+10Hz 0.986144 -0.133977
+ 6.32e+10Hz 0.986112 -0.134187
+ 6.33e+10Hz 0.986081 -0.134396
+ 6.34e+10Hz 0.98605 -0.134605
+ 6.35e+10Hz 0.986019 -0.134814
+ 6.36e+10Hz 0.985988 -0.135023
+ 6.37e+10Hz 0.985957 -0.135233
+ 6.38e+10Hz 0.985925 -0.135442
+ 6.39e+10Hz 0.985894 -0.135651
+ 6.4e+10Hz 0.985863 -0.13586
+ 6.41e+10Hz 0.985831 -0.136069
+ 6.42e+10Hz 0.9858 -0.136278
+ 6.43e+10Hz 0.985768 -0.136488
+ 6.44e+10Hz 0.985737 -0.136697
+ 6.45e+10Hz 0.985705 -0.136906
+ 6.46e+10Hz 0.985673 -0.137115
+ 6.47e+10Hz 0.985642 -0.137324
+ 6.48e+10Hz 0.98561 -0.137533
+ 6.49e+10Hz 0.985578 -0.137742
+ 6.5e+10Hz 0.985546 -0.137951
+ 6.51e+10Hz 0.985514 -0.13816
+ 6.52e+10Hz 0.985483 -0.138369
+ 6.53e+10Hz 0.985451 -0.138578
+ 6.54e+10Hz 0.985419 -0.138788
+ 6.55e+10Hz 0.985387 -0.138996
+ 6.56e+10Hz 0.985355 -0.139206
+ 6.57e+10Hz 0.985322 -0.139415
+ 6.58e+10Hz 0.98529 -0.139624
+ 6.59e+10Hz 0.985258 -0.139833
+ 6.6e+10Hz 0.985226 -0.140042
+ 6.61e+10Hz 0.985194 -0.140251
+ 6.62e+10Hz 0.985161 -0.14046
+ 6.63e+10Hz 0.985129 -0.140669
+ 6.64e+10Hz 0.985097 -0.140878
+ 6.65e+10Hz 0.985064 -0.141087
+ 6.66e+10Hz 0.985032 -0.141296
+ 6.67e+10Hz 0.984999 -0.141505
+ 6.68e+10Hz 0.984966 -0.141714
+ 6.69e+10Hz 0.984934 -0.141923
+ 6.7e+10Hz 0.984901 -0.142131
+ 6.71e+10Hz 0.984869 -0.142341
+ 6.72e+10Hz 0.984836 -0.142549
+ 6.73e+10Hz 0.984803 -0.142758
+ 6.74e+10Hz 0.98477 -0.142967
+ 6.75e+10Hz 0.984737 -0.143176
+ 6.76e+10Hz 0.984704 -0.143385
+ 6.77e+10Hz 0.984671 -0.143594
+ 6.78e+10Hz 0.984638 -0.143803
+ 6.79e+10Hz 0.984605 -0.144012
+ 6.8e+10Hz 0.984572 -0.144221
+ 6.81e+10Hz 0.984539 -0.14443
+ 6.82e+10Hz 0.984506 -0.144639
+ 6.83e+10Hz 0.984472 -0.144847
+ 6.84e+10Hz 0.984439 -0.145056
+ 6.85e+10Hz 0.984406 -0.145265
+ 6.86e+10Hz 0.984372 -0.145474
+ 6.87e+10Hz 0.984339 -0.145683
+ 6.88e+10Hz 0.984306 -0.145892
+ 6.89e+10Hz 0.984272 -0.146101
+ 6.9e+10Hz 0.984238 -0.14631
+ 6.91e+10Hz 0.984205 -0.146518
+ 6.92e+10Hz 0.984171 -0.146727
+ 6.93e+10Hz 0.984137 -0.146936
+ 6.94e+10Hz 0.984104 -0.147145
+ 6.95e+10Hz 0.98407 -0.147354
+ 6.96e+10Hz 0.984036 -0.147563
+ 6.97e+10Hz 0.984002 -0.147771
+ 6.98e+10Hz 0.983968 -0.14798
+ 6.99e+10Hz 0.983934 -0.148189
+ 7e+10Hz 0.9839 -0.148398
+ 7.01e+10Hz 0.983866 -0.148607
+ 7.02e+10Hz 0.983832 -0.148815
+ 7.03e+10Hz 0.983798 -0.149024
+ 7.04e+10Hz 0.983763 -0.149233
+ 7.05e+10Hz 0.983729 -0.149442
+ 7.06e+10Hz 0.983695 -0.14965
+ 7.07e+10Hz 0.98366 -0.149859
+ 7.08e+10Hz 0.983626 -0.150068
+ 7.09e+10Hz 0.983591 -0.150277
+ 7.1e+10Hz 0.983557 -0.150485
+ 7.11e+10Hz 0.983522 -0.150694
+ 7.12e+10Hz 0.983488 -0.150903
+ 7.13e+10Hz 0.983453 -0.151112
+ 7.14e+10Hz 0.983418 -0.15132
+ 7.15e+10Hz 0.983383 -0.151529
+ 7.16e+10Hz 0.983349 -0.151738
+ 7.17e+10Hz 0.983314 -0.151947
+ 7.18e+10Hz 0.983279 -0.152155
+ 7.19e+10Hz 0.983244 -0.152364
+ 7.2e+10Hz 0.983209 -0.152572
+ 7.21e+10Hz 0.983174 -0.152781
+ 7.22e+10Hz 0.983139 -0.15299
+ 7.23e+10Hz 0.983104 -0.153198
+ 7.24e+10Hz 0.983068 -0.153407
+ 7.25e+10Hz 0.983033 -0.153616
+ 7.26e+10Hz 0.982998 -0.153824
+ 7.27e+10Hz 0.982962 -0.154033
+ 7.28e+10Hz 0.982927 -0.154242
+ 7.29e+10Hz 0.982891 -0.15445
+ 7.3e+10Hz 0.982856 -0.154659
+ 7.31e+10Hz 0.98282 -0.154867
+ 7.32e+10Hz 0.982785 -0.155076
+ 7.33e+10Hz 0.982749 -0.155284
+ 7.34e+10Hz 0.982713 -0.155493
+ 7.35e+10Hz 0.982677 -0.155702
+ 7.36e+10Hz 0.982641 -0.15591
+ 7.37e+10Hz 0.982606 -0.156119
+ 7.38e+10Hz 0.98257 -0.156327
+ 7.39e+10Hz 0.982534 -0.156536
+ 7.4e+10Hz 0.982498 -0.156744
+ 7.41e+10Hz 0.982462 -0.156953
+ 7.42e+10Hz 0.982425 -0.157161
+ 7.43e+10Hz 0.982389 -0.15737
+ 7.44e+10Hz 0.982353 -0.157578
+ 7.45e+10Hz 0.982317 -0.157786
+ 7.46e+10Hz 0.98228 -0.157995
+ 7.47e+10Hz 0.982244 -0.158203
+ 7.48e+10Hz 0.982208 -0.158412
+ 7.49e+10Hz 0.982171 -0.15862
+ 7.5e+10Hz 0.982134 -0.158829
+ 7.51e+10Hz 0.982098 -0.159037
+ 7.52e+10Hz 0.982061 -0.159245
+ 7.53e+10Hz 0.982024 -0.159454
+ 7.54e+10Hz 0.981988 -0.159662
+ 7.55e+10Hz 0.981951 -0.15987
+ 7.56e+10Hz 0.981914 -0.160079
+ 7.57e+10Hz 0.981877 -0.160287
+ 7.58e+10Hz 0.98184 -0.160495
+ 7.59e+10Hz 0.981803 -0.160704
+ 7.6e+10Hz 0.981766 -0.160912
+ 7.61e+10Hz 0.981729 -0.16112
+ 7.62e+10Hz 0.981692 -0.161329
+ 7.63e+10Hz 0.981654 -0.161537
+ 7.64e+10Hz 0.981617 -0.161745
+ 7.65e+10Hz 0.98158 -0.161953
+ 7.66e+10Hz 0.981542 -0.162161
+ 7.67e+10Hz 0.981505 -0.16237
+ 7.68e+10Hz 0.981468 -0.162578
+ 7.69e+10Hz 0.98143 -0.162786
+ 7.7e+10Hz 0.981393 -0.162994
+ 7.71e+10Hz 0.981355 -0.163202
+ 7.72e+10Hz 0.981317 -0.16341
+ 7.73e+10Hz 0.981279 -0.163619
+ 7.74e+10Hz 0.981242 -0.163827
+ 7.75e+10Hz 0.981204 -0.164035
+ 7.76e+10Hz 0.981166 -0.164243
+ 7.77e+10Hz 0.981128 -0.164451
+ 7.78e+10Hz 0.98109 -0.164659
+ 7.79e+10Hz 0.981052 -0.164867
+ 7.8e+10Hz 0.981014 -0.165075
+ 7.81e+10Hz 0.980976 -0.165283
+ 7.82e+10Hz 0.980938 -0.165491
+ 7.83e+10Hz 0.980899 -0.165699
+ 7.84e+10Hz 0.980861 -0.165907
+ 7.85e+10Hz 0.980823 -0.166115
+ 7.86e+10Hz 0.980784 -0.166323
+ 7.87e+10Hz 0.980746 -0.166531
+ 7.88e+10Hz 0.980707 -0.166739
+ 7.89e+10Hz 0.980669 -0.166947
+ 7.9e+10Hz 0.98063 -0.167155
+ 7.91e+10Hz 0.980592 -0.167362
+ 7.92e+10Hz 0.980553 -0.16757
+ 7.93e+10Hz 0.980514 -0.167778
+ 7.94e+10Hz 0.980476 -0.167986
+ 7.95e+10Hz 0.980437 -0.168194
+ 7.96e+10Hz 0.980398 -0.168402
+ 7.97e+10Hz 0.980359 -0.168609
+ 7.98e+10Hz 0.98032 -0.168817
+ 7.99e+10Hz 0.980281 -0.169025
+ 8e+10Hz 0.980242 -0.169233
+ 8.01e+10Hz 0.980203 -0.16944
+ 8.02e+10Hz 0.980163 -0.169648
+ 8.03e+10Hz 0.980124 -0.169856
+ 8.04e+10Hz 0.980085 -0.170064
+ 8.05e+10Hz 0.980046 -0.170271
+ 8.06e+10Hz 0.980006 -0.170479
+ 8.07e+10Hz 0.979967 -0.170686
+ 8.08e+10Hz 0.979928 -0.170894
+ 8.09e+10Hz 0.979888 -0.171102
+ 8.1e+10Hz 0.979849 -0.171309
+ 8.11e+10Hz 0.979809 -0.171517
+ 8.12e+10Hz 0.979769 -0.171724
+ 8.13e+10Hz 0.97973 -0.171932
+ 8.14e+10Hz 0.97969 -0.17214
+ 8.15e+10Hz 0.97965 -0.172347
+ 8.16e+10Hz 0.97961 -0.172554
+ 8.17e+10Hz 0.97957 -0.172762
+ 8.18e+10Hz 0.97953 -0.172969
+ 8.19e+10Hz 0.979491 -0.173177
+ 8.2e+10Hz 0.979451 -0.173384
+ 8.21e+10Hz 0.97941 -0.173592
+ 8.22e+10Hz 0.97937 -0.173799
+ 8.23e+10Hz 0.97933 -0.174007
+ 8.24e+10Hz 0.97929 -0.174214
+ 8.25e+10Hz 0.97925 -0.174421
+ 8.26e+10Hz 0.979209 -0.174629
+ 8.27e+10Hz 0.979169 -0.174836
+ 8.28e+10Hz 0.979129 -0.175043
+ 8.29e+10Hz 0.979088 -0.175251
+ 8.3e+10Hz 0.979048 -0.175458
+ 8.31e+10Hz 0.979007 -0.175665
+ 8.32e+10Hz 0.978967 -0.175872
+ 8.33e+10Hz 0.978926 -0.17608
+ 8.34e+10Hz 0.978886 -0.176287
+ 8.35e+10Hz 0.978845 -0.176494
+ 8.36e+10Hz 0.978804 -0.176701
+ 8.37e+10Hz 0.978763 -0.176908
+ 8.38e+10Hz 0.978723 -0.177116
+ 8.39e+10Hz 0.978682 -0.177323
+ 8.4e+10Hz 0.978641 -0.17753
+ 8.41e+10Hz 0.9786 -0.177737
+ 8.42e+10Hz 0.978559 -0.177944
+ 8.43e+10Hz 0.978518 -0.178151
+ 8.44e+10Hz 0.978477 -0.178358
+ 8.45e+10Hz 0.978436 -0.178565
+ 8.46e+10Hz 0.978394 -0.178773
+ 8.47e+10Hz 0.978353 -0.17898
+ 8.48e+10Hz 0.978312 -0.179187
+ 8.49e+10Hz 0.978271 -0.179394
+ 8.5e+10Hz 0.978229 -0.179601
+ 8.51e+10Hz 0.978188 -0.179808
+ 8.52e+10Hz 0.978147 -0.180015
+ 8.53e+10Hz 0.978105 -0.180222
+ 8.54e+10Hz 0.978064 -0.180428
+ 8.55e+10Hz 0.978022 -0.180636
+ 8.56e+10Hz 0.97798 -0.180842
+ 8.57e+10Hz 0.977939 -0.181049
+ 8.58e+10Hz 0.977897 -0.181256
+ 8.59e+10Hz 0.977855 -0.181463
+ 8.6e+10Hz 0.977814 -0.18167
+ 8.61e+10Hz 0.977772 -0.181877
+ 8.62e+10Hz 0.97773 -0.182084
+ 8.63e+10Hz 0.977688 -0.182291
+ 8.64e+10Hz 0.977646 -0.182497
+ 8.65e+10Hz 0.977604 -0.182704
+ 8.66e+10Hz 0.977562 -0.182911
+ 8.67e+10Hz 0.97752 -0.183118
+ 8.68e+10Hz 0.977478 -0.183325
+ 8.69e+10Hz 0.977436 -0.183531
+ 8.7e+10Hz 0.977394 -0.183738
+ 8.71e+10Hz 0.977351 -0.183945
+ 8.72e+10Hz 0.977309 -0.184152
+ 8.73e+10Hz 0.977267 -0.184358
+ 8.74e+10Hz 0.977224 -0.184565
+ 8.75e+10Hz 0.977182 -0.184772
+ 8.76e+10Hz 0.97714 -0.184978
+ 8.77e+10Hz 0.977097 -0.185185
+ 8.78e+10Hz 0.977055 -0.185392
+ 8.79e+10Hz 0.977012 -0.185598
+ 8.8e+10Hz 0.976969 -0.185805
+ 8.81e+10Hz 0.976927 -0.186012
+ 8.82e+10Hz 0.976884 -0.186218
+ 8.83e+10Hz 0.976841 -0.186425
+ 8.84e+10Hz 0.976799 -0.186632
+ 8.85e+10Hz 0.976756 -0.186838
+ 8.86e+10Hz 0.976713 -0.187045
+ 8.87e+10Hz 0.97667 -0.187251
+ 8.88e+10Hz 0.976627 -0.187458
+ 8.89e+10Hz 0.976584 -0.187665
+ 8.9e+10Hz 0.976541 -0.187871
+ 8.91e+10Hz 0.976498 -0.188078
+ 8.92e+10Hz 0.976455 -0.188284
+ 8.93e+10Hz 0.976412 -0.188491
+ 8.94e+10Hz 0.976368 -0.188697
+ 8.95e+10Hz 0.976325 -0.188904
+ 8.96e+10Hz 0.976282 -0.18911
+ 8.97e+10Hz 0.976239 -0.189317
+ 8.98e+10Hz 0.976195 -0.189523
+ 8.99e+10Hz 0.976152 -0.18973
+ 9e+10Hz 0.976108 -0.189936
+ 9.01e+10Hz 0.976065 -0.190143
+ 9.02e+10Hz 0.976021 -0.190349
+ 9.03e+10Hz 0.975978 -0.190556
+ 9.04e+10Hz 0.975934 -0.190762
+ 9.05e+10Hz 0.97589 -0.190969
+ 9.06e+10Hz 0.975847 -0.191175
+ 9.07e+10Hz 0.975803 -0.191382
+ 9.08e+10Hz 0.975759 -0.191588
+ 9.09e+10Hz 0.975715 -0.191794
+ 9.1e+10Hz 0.975672 -0.192001
+ 9.11e+10Hz 0.975627 -0.192207
+ 9.12e+10Hz 0.975584 -0.192414
+ 9.13e+10Hz 0.97554 -0.19262
+ 9.14e+10Hz 0.975495 -0.192826
+ 9.15e+10Hz 0.975451 -0.193033
+ 9.16e+10Hz 0.975407 -0.193239
+ 9.17e+10Hz 0.975363 -0.193445
+ 9.18e+10Hz 0.975319 -0.193652
+ 9.19e+10Hz 0.975275 -0.193858
+ 9.2e+10Hz 0.97523 -0.194065
+ 9.21e+10Hz 0.975186 -0.194271
+ 9.22e+10Hz 0.975141 -0.194477
+ 9.23e+10Hz 0.975097 -0.194684
+ 9.24e+10Hz 0.975052 -0.19489
+ 9.25e+10Hz 0.975008 -0.195096
+ 9.26e+10Hz 0.974963 -0.195302
+ 9.27e+10Hz 0.974919 -0.195509
+ 9.28e+10Hz 0.974874 -0.195715
+ 9.29e+10Hz 0.974829 -0.195921
+ 9.3e+10Hz 0.974785 -0.196128
+ 9.31e+10Hz 0.97474 -0.196334
+ 9.32e+10Hz 0.974695 -0.19654
+ 9.33e+10Hz 0.97465 -0.196746
+ 9.34e+10Hz 0.974605 -0.196953
+ 9.35e+10Hz 0.97456 -0.197159
+ 9.36e+10Hz 0.974515 -0.197365
+ 9.37e+10Hz 0.97447 -0.197572
+ 9.38e+10Hz 0.974425 -0.197778
+ 9.39e+10Hz 0.974379 -0.197984
+ 9.4e+10Hz 0.974334 -0.19819
+ 9.41e+10Hz 0.974289 -0.198397
+ 9.42e+10Hz 0.974244 -0.198603
+ 9.43e+10Hz 0.974198 -0.198809
+ 9.44e+10Hz 0.974153 -0.199015
+ 9.45e+10Hz 0.974107 -0.199221
+ 9.46e+10Hz 0.974062 -0.199428
+ 9.47e+10Hz 0.974016 -0.199634
+ 9.48e+10Hz 0.973971 -0.19984
+ 9.49e+10Hz 0.973925 -0.200046
+ 9.5e+10Hz 0.973879 -0.200252
+ 9.51e+10Hz 0.973834 -0.200458
+ 9.52e+10Hz 0.973788 -0.200665
+ 9.53e+10Hz 0.973742 -0.200871
+ 9.54e+10Hz 0.973696 -0.201077
+ 9.55e+10Hz 0.97365 -0.201283
+ 9.56e+10Hz 0.973604 -0.201489
+ 9.57e+10Hz 0.973558 -0.201695
+ 9.58e+10Hz 0.973512 -0.201901
+ 9.59e+10Hz 0.973466 -0.202107
+ 9.6e+10Hz 0.97342 -0.202314
+ 9.61e+10Hz 0.973374 -0.20252
+ 9.62e+10Hz 0.973327 -0.202726
+ 9.63e+10Hz 0.973281 -0.202932
+ 9.64e+10Hz 0.973235 -0.203138
+ 9.65e+10Hz 0.973188 -0.203344
+ 9.66e+10Hz 0.973142 -0.20355
+ 9.67e+10Hz 0.973095 -0.203756
+ 9.68e+10Hz 0.973048 -0.203962
+ 9.69e+10Hz 0.973002 -0.204168
+ 9.7e+10Hz 0.972955 -0.204374
+ 9.71e+10Hz 0.972908 -0.20458
+ 9.72e+10Hz 0.972862 -0.204786
+ 9.73e+10Hz 0.972815 -0.204992
+ 9.74e+10Hz 0.972768 -0.205198
+ 9.75e+10Hz 0.972721 -0.205404
+ 9.76e+10Hz 0.972674 -0.20561
+ 9.77e+10Hz 0.972627 -0.205816
+ 9.78e+10Hz 0.97258 -0.206022
+ 9.79e+10Hz 0.972533 -0.206228
+ 9.8e+10Hz 0.972486 -0.206434
+ 9.81e+10Hz 0.972438 -0.20664
+ 9.82e+10Hz 0.972391 -0.206846
+ 9.83e+10Hz 0.972344 -0.207052
+ 9.84e+10Hz 0.972296 -0.207258
+ 9.85e+10Hz 0.972249 -0.207464
+ 9.86e+10Hz 0.972202 -0.20767
+ 9.87e+10Hz 0.972154 -0.207876
+ 9.88e+10Hz 0.972106 -0.208082
+ 9.89e+10Hz 0.972059 -0.208287
+ 9.9e+10Hz 0.972011 -0.208493
+ 9.91e+10Hz 0.971963 -0.208699
+ 9.92e+10Hz 0.971916 -0.208905
+ 9.93e+10Hz 0.971868 -0.209111
+ 9.94e+10Hz 0.97182 -0.209317
+ 9.95e+10Hz 0.971772 -0.209523
+ 9.96e+10Hz 0.971724 -0.209728
+ 9.97e+10Hz 0.971676 -0.209934
+ 9.98e+10Hz 0.971628 -0.21014
+ 9.99e+10Hz 0.97158 -0.210346
+ 1e+11Hz 0.971531 -0.210551
+ 1.001e+11Hz 0.971483 -0.210757
+ 1.002e+11Hz 0.971435 -0.210963
+ 1.003e+11Hz 0.971387 -0.211169
+ 1.004e+11Hz 0.971338 -0.211374
+ 1.005e+11Hz 0.97129 -0.21158
+ 1.006e+11Hz 0.971241 -0.211786
+ 1.007e+11Hz 0.971193 -0.211991
+ 1.008e+11Hz 0.971144 -0.212197
+ 1.009e+11Hz 0.971096 -0.212403
+ 1.01e+11Hz 0.971047 -0.212608
+ 1.011e+11Hz 0.970998 -0.212814
+ 1.012e+11Hz 0.970949 -0.21302
+ 1.013e+11Hz 0.9709 -0.213225
+ 1.014e+11Hz 0.970851 -0.213431
+ 1.015e+11Hz 0.970803 -0.213636
+ 1.016e+11Hz 0.970754 -0.213842
+ 1.017e+11Hz 0.970704 -0.214047
+ 1.018e+11Hz 0.970655 -0.214253
+ 1.019e+11Hz 0.970606 -0.214458
+ 1.02e+11Hz 0.970557 -0.214664
+ 1.021e+11Hz 0.970508 -0.214869
+ 1.022e+11Hz 0.970459 -0.215075
+ 1.023e+11Hz 0.970409 -0.21528
+ 1.024e+11Hz 0.97036 -0.215486
+ 1.025e+11Hz 0.97031 -0.215691
+ 1.026e+11Hz 0.970261 -0.215897
+ 1.027e+11Hz 0.970211 -0.216102
+ 1.028e+11Hz 0.970162 -0.216307
+ 1.029e+11Hz 0.970112 -0.216513
+ 1.03e+11Hz 0.970062 -0.216718
+ 1.031e+11Hz 0.970013 -0.216923
+ 1.032e+11Hz 0.969963 -0.217129
+ 1.033e+11Hz 0.969913 -0.217334
+ 1.034e+11Hz 0.969863 -0.217539
+ 1.035e+11Hz 0.969813 -0.217745
+ 1.036e+11Hz 0.969763 -0.21795
+ 1.037e+11Hz 0.969713 -0.218155
+ 1.038e+11Hz 0.969663 -0.21836
+ 1.039e+11Hz 0.969613 -0.218565
+ 1.04e+11Hz 0.969563 -0.218771
+ 1.041e+11Hz 0.969513 -0.218976
+ 1.042e+11Hz 0.969462 -0.219181
+ 1.043e+11Hz 0.969412 -0.219386
+ 1.044e+11Hz 0.969362 -0.219591
+ 1.045e+11Hz 0.969311 -0.219796
+ 1.046e+11Hz 0.969261 -0.220001
+ 1.047e+11Hz 0.96921 -0.220206
+ 1.048e+11Hz 0.96916 -0.220411
+ 1.049e+11Hz 0.969109 -0.220616
+ 1.05e+11Hz 0.969059 -0.220821
+ 1.051e+11Hz 0.969008 -0.221026
+ 1.052e+11Hz 0.968957 -0.221231
+ 1.053e+11Hz 0.968906 -0.221436
+ 1.054e+11Hz 0.968856 -0.221641
+ 1.055e+11Hz 0.968805 -0.221846
+ 1.056e+11Hz 0.968754 -0.222051
+ 1.057e+11Hz 0.968703 -0.222256
+ 1.058e+11Hz 0.968652 -0.222461
+ 1.059e+11Hz 0.968601 -0.222666
+ 1.06e+11Hz 0.96855 -0.22287
+ 1.061e+11Hz 0.968499 -0.223075
+ 1.062e+11Hz 0.968448 -0.22328
+ 1.063e+11Hz 0.968396 -0.223485
+ 1.064e+11Hz 0.968345 -0.22369
+ 1.065e+11Hz 0.968294 -0.223894
+ 1.066e+11Hz 0.968242 -0.224099
+ 1.067e+11Hz 0.968191 -0.224304
+ 1.068e+11Hz 0.96814 -0.224508
+ 1.069e+11Hz 0.968088 -0.224713
+ 1.07e+11Hz 0.968036 -0.224918
+ 1.071e+11Hz 0.967985 -0.225122
+ 1.072e+11Hz 0.967933 -0.225327
+ 1.073e+11Hz 0.967882 -0.225531
+ 1.074e+11Hz 0.96783 -0.225736
+ 1.075e+11Hz 0.967778 -0.22594
+ 1.076e+11Hz 0.967727 -0.226145
+ 1.077e+11Hz 0.967675 -0.226349
+ 1.078e+11Hz 0.967623 -0.226554
+ 1.079e+11Hz 0.967571 -0.226758
+ 1.08e+11Hz 0.967519 -0.226963
+ 1.081e+11Hz 0.967467 -0.227167
+ 1.082e+11Hz 0.967415 -0.227372
+ 1.083e+11Hz 0.967363 -0.227576
+ 1.084e+11Hz 0.967311 -0.22778
+ 1.085e+11Hz 0.967259 -0.227985
+ 1.086e+11Hz 0.967207 -0.228189
+ 1.087e+11Hz 0.967155 -0.228393
+ 1.088e+11Hz 0.967102 -0.228598
+ 1.089e+11Hz 0.96705 -0.228802
+ 1.09e+11Hz 0.966998 -0.229006
+ 1.091e+11Hz 0.966945 -0.22921
+ 1.092e+11Hz 0.966893 -0.229415
+ 1.093e+11Hz 0.96684 -0.229619
+ 1.094e+11Hz 0.966788 -0.229823
+ 1.095e+11Hz 0.966735 -0.230027
+ 1.096e+11Hz 0.966683 -0.230231
+ 1.097e+11Hz 0.96663 -0.230435
+ 1.098e+11Hz 0.966578 -0.23064
+ 1.099e+11Hz 0.966525 -0.230844
+ 1.1e+11Hz 0.966472 -0.231048
+ 1.101e+11Hz 0.96642 -0.231252
+ 1.102e+11Hz 0.966367 -0.231456
+ 1.103e+11Hz 0.966314 -0.23166
+ 1.104e+11Hz 0.966261 -0.231864
+ 1.105e+11Hz 0.966208 -0.232068
+ 1.106e+11Hz 0.966155 -0.232272
+ 1.107e+11Hz 0.966102 -0.232476
+ 1.108e+11Hz 0.96605 -0.23268
+ 1.109e+11Hz 0.965997 -0.232884
+ 1.11e+11Hz 0.965943 -0.233088
+ 1.111e+11Hz 0.96589 -0.233292
+ 1.112e+11Hz 0.965837 -0.233495
+ 1.113e+11Hz 0.965784 -0.233699
+ 1.114e+11Hz 0.965731 -0.233903
+ 1.115e+11Hz 0.965678 -0.234107
+ 1.116e+11Hz 0.965624 -0.234311
+ 1.117e+11Hz 0.965571 -0.234515
+ 1.118e+11Hz 0.965518 -0.234718
+ 1.119e+11Hz 0.965464 -0.234922
+ 1.12e+11Hz 0.965411 -0.235126
+ 1.121e+11Hz 0.965357 -0.23533
+ 1.122e+11Hz 0.965304 -0.235533
+ 1.123e+11Hz 0.96525 -0.235737
+ 1.124e+11Hz 0.965197 -0.235941
+ 1.125e+11Hz 0.965143 -0.236145
+ 1.126e+11Hz 0.96509 -0.236348
+ 1.127e+11Hz 0.965036 -0.236552
+ 1.128e+11Hz 0.964982 -0.236756
+ 1.129e+11Hz 0.964928 -0.236959
+ 1.13e+11Hz 0.964875 -0.237163
+ 1.131e+11Hz 0.964821 -0.237366
+ 1.132e+11Hz 0.964767 -0.23757
+ 1.133e+11Hz 0.964713 -0.237774
+ 1.134e+11Hz 0.964659 -0.237977
+ 1.135e+11Hz 0.964605 -0.238181
+ 1.136e+11Hz 0.964551 -0.238384
+ 1.137e+11Hz 0.964497 -0.238588
+ 1.138e+11Hz 0.964443 -0.238791
+ 1.139e+11Hz 0.964389 -0.238995
+ 1.14e+11Hz 0.964335 -0.239198
+ 1.141e+11Hz 0.964281 -0.239402
+ 1.142e+11Hz 0.964227 -0.239605
+ 1.143e+11Hz 0.964173 -0.239809
+ 1.144e+11Hz 0.964118 -0.240012
+ 1.145e+11Hz 0.964064 -0.240216
+ 1.146e+11Hz 0.96401 -0.240419
+ 1.147e+11Hz 0.963955 -0.240623
+ 1.148e+11Hz 0.963901 -0.240826
+ 1.149e+11Hz 0.963847 -0.24103
+ 1.15e+11Hz 0.963792 -0.241233
+ 1.151e+11Hz 0.963738 -0.241436
+ 1.152e+11Hz 0.963683 -0.24164
+ 1.153e+11Hz 0.963628 -0.241843
+ 1.154e+11Hz 0.963574 -0.242046
+ 1.155e+11Hz 0.963519 -0.24225
+ 1.156e+11Hz 0.963464 -0.242453
+ 1.157e+11Hz 0.96341 -0.242657
+ 1.158e+11Hz 0.963355 -0.24286
+ 1.159e+11Hz 0.9633 -0.243063
+ 1.16e+11Hz 0.963245 -0.243267
+ 1.161e+11Hz 0.963191 -0.24347
+ 1.162e+11Hz 0.963136 -0.243673
+ 1.163e+11Hz 0.963081 -0.243876
+ 1.164e+11Hz 0.963026 -0.24408
+ 1.165e+11Hz 0.962971 -0.244283
+ 1.166e+11Hz 0.962916 -0.244486
+ 1.167e+11Hz 0.962861 -0.24469
+ 1.168e+11Hz 0.962805 -0.244893
+ 1.169e+11Hz 0.96275 -0.245096
+ 1.17e+11Hz 0.962695 -0.245299
+ 1.171e+11Hz 0.96264 -0.245503
+ 1.172e+11Hz 0.962584 -0.245706
+ 1.173e+11Hz 0.962529 -0.245909
+ 1.174e+11Hz 0.962474 -0.246112
+ 1.175e+11Hz 0.962418 -0.246316
+ 1.176e+11Hz 0.962363 -0.246519
+ 1.177e+11Hz 0.962307 -0.246722
+ 1.178e+11Hz 0.962252 -0.246925
+ 1.179e+11Hz 0.962196 -0.247128
+ 1.18e+11Hz 0.962141 -0.247332
+ 1.181e+11Hz 0.962085 -0.247535
+ 1.182e+11Hz 0.962029 -0.247738
+ 1.183e+11Hz 0.961974 -0.247941
+ 1.184e+11Hz 0.961918 -0.248144
+ 1.185e+11Hz 0.961862 -0.248347
+ 1.186e+11Hz 0.961806 -0.248551
+ 1.187e+11Hz 0.96175 -0.248754
+ 1.188e+11Hz 0.961694 -0.248957
+ 1.189e+11Hz 0.961638 -0.24916
+ 1.19e+11Hz 0.961582 -0.249363
+ 1.191e+11Hz 0.961526 -0.249566
+ 1.192e+11Hz 0.96147 -0.249769
+ 1.193e+11Hz 0.961414 -0.249972
+ 1.194e+11Hz 0.961358 -0.250175
+ 1.195e+11Hz 0.961302 -0.250379
+ 1.196e+11Hz 0.961245 -0.250582
+ 1.197e+11Hz 0.961189 -0.250785
+ 1.198e+11Hz 0.961132 -0.250988
+ 1.199e+11Hz 0.961076 -0.251191
+ 1.2e+11Hz 0.96102 -0.251394
+ 1.201e+11Hz 0.960963 -0.251597
+ 1.202e+11Hz 0.960906 -0.2518
+ 1.203e+11Hz 0.96085 -0.252003
+ 1.204e+11Hz 0.960793 -0.252206
+ 1.205e+11Hz 0.960737 -0.252409
+ 1.206e+11Hz 0.96068 -0.252612
+ 1.207e+11Hz 0.960623 -0.252815
+ 1.208e+11Hz 0.960566 -0.253018
+ 1.209e+11Hz 0.960509 -0.253221
+ 1.21e+11Hz 0.960452 -0.253424
+ 1.211e+11Hz 0.960395 -0.253627
+ 1.212e+11Hz 0.960338 -0.25383
+ 1.213e+11Hz 0.960281 -0.254033
+ 1.214e+11Hz 0.960224 -0.254236
+ 1.215e+11Hz 0.960167 -0.254439
+ 1.216e+11Hz 0.96011 -0.254642
+ 1.217e+11Hz 0.960052 -0.254845
+ 1.218e+11Hz 0.959995 -0.255048
+ 1.219e+11Hz 0.959938 -0.25525
+ 1.22e+11Hz 0.95988 -0.255453
+ 1.221e+11Hz 0.959823 -0.255656
+ 1.222e+11Hz 0.959765 -0.255859
+ 1.223e+11Hz 0.959708 -0.256062
+ 1.224e+11Hz 0.95965 -0.256265
+ 1.225e+11Hz 0.959592 -0.256468
+ 1.226e+11Hz 0.959534 -0.256671
+ 1.227e+11Hz 0.959477 -0.256873
+ 1.228e+11Hz 0.959419 -0.257076
+ 1.229e+11Hz 0.959361 -0.257279
+ 1.23e+11Hz 0.959303 -0.257482
+ 1.231e+11Hz 0.959245 -0.257684
+ 1.232e+11Hz 0.959187 -0.257887
+ 1.233e+11Hz 0.959129 -0.25809
+ 1.234e+11Hz 0.959071 -0.258293
+ 1.235e+11Hz 0.959012 -0.258495
+ 1.236e+11Hz 0.958954 -0.258698
+ 1.237e+11Hz 0.958896 -0.258901
+ 1.238e+11Hz 0.958837 -0.259103
+ 1.239e+11Hz 0.958779 -0.259306
+ 1.24e+11Hz 0.95872 -0.259509
+ 1.241e+11Hz 0.958662 -0.259711
+ 1.242e+11Hz 0.958603 -0.259914
+ 1.243e+11Hz 0.958545 -0.260117
+ 1.244e+11Hz 0.958486 -0.260319
+ 1.245e+11Hz 0.958427 -0.260522
+ 1.246e+11Hz 0.958368 -0.260724
+ 1.247e+11Hz 0.95831 -0.260927
+ 1.248e+11Hz 0.958251 -0.261129
+ 1.249e+11Hz 0.958192 -0.261332
+ 1.25e+11Hz 0.958133 -0.261534
+ 1.251e+11Hz 0.958073 -0.261737
+ 1.252e+11Hz 0.958014 -0.261939
+ 1.253e+11Hz 0.957955 -0.262142
+ 1.254e+11Hz 0.957896 -0.262344
+ 1.255e+11Hz 0.957836 -0.262546
+ 1.256e+11Hz 0.957777 -0.262749
+ 1.257e+11Hz 0.957718 -0.262951
+ 1.258e+11Hz 0.957658 -0.263153
+ 1.259e+11Hz 0.957599 -0.263356
+ 1.26e+11Hz 0.957539 -0.263558
+ 1.261e+11Hz 0.95748 -0.26376
+ 1.262e+11Hz 0.95742 -0.263962
+ 1.263e+11Hz 0.95736 -0.264165
+ 1.264e+11Hz 0.9573 -0.264367
+ 1.265e+11Hz 0.95724 -0.264569
+ 1.266e+11Hz 0.95718 -0.264771
+ 1.267e+11Hz 0.95712 -0.264973
+ 1.268e+11Hz 0.95706 -0.265175
+ 1.269e+11Hz 0.957 -0.265377
+ 1.27e+11Hz 0.95694 -0.265579
+ 1.271e+11Hz 0.95688 -0.265781
+ 1.272e+11Hz 0.95682 -0.265983
+ 1.273e+11Hz 0.956759 -0.266185
+ 1.274e+11Hz 0.956699 -0.266387
+ 1.275e+11Hz 0.956639 -0.266589
+ 1.276e+11Hz 0.956578 -0.266791
+ 1.277e+11Hz 0.956518 -0.266993
+ 1.278e+11Hz 0.956457 -0.267195
+ 1.279e+11Hz 0.956396 -0.267396
+ 1.28e+11Hz 0.956336 -0.267598
+ 1.281e+11Hz 0.956275 -0.2678
+ 1.282e+11Hz 0.956214 -0.268002
+ 1.283e+11Hz 0.956153 -0.268203
+ 1.284e+11Hz 0.956092 -0.268405
+ 1.285e+11Hz 0.956032 -0.268607
+ 1.286e+11Hz 0.95597 -0.268808
+ 1.287e+11Hz 0.955909 -0.26901
+ 1.288e+11Hz 0.955848 -0.269211
+ 1.289e+11Hz 0.955787 -0.269413
+ 1.29e+11Hz 0.955726 -0.269614
+ 1.291e+11Hz 0.955665 -0.269816
+ 1.292e+11Hz 0.955603 -0.270017
+ 1.293e+11Hz 0.955542 -0.270218
+ 1.294e+11Hz 0.955481 -0.27042
+ 1.295e+11Hz 0.955419 -0.270621
+ 1.296e+11Hz 0.955358 -0.270822
+ 1.297e+11Hz 0.955296 -0.271023
+ 1.298e+11Hz 0.955234 -0.271225
+ 1.299e+11Hz 0.955173 -0.271426
+ 1.3e+11Hz 0.955111 -0.271627
+ 1.301e+11Hz 0.955049 -0.271828
+ 1.302e+11Hz 0.954987 -0.272029
+ 1.303e+11Hz 0.954926 -0.27223
+ 1.304e+11Hz 0.954864 -0.272431
+ 1.305e+11Hz 0.954802 -0.272632
+ 1.306e+11Hz 0.95474 -0.272833
+ 1.307e+11Hz 0.954678 -0.273034
+ 1.308e+11Hz 0.954616 -0.273235
+ 1.309e+11Hz 0.954554 -0.273436
+ 1.31e+11Hz 0.954491 -0.273636
+ 1.311e+11Hz 0.954429 -0.273837
+ 1.312e+11Hz 0.954367 -0.274038
+ 1.313e+11Hz 0.954304 -0.274238
+ 1.314e+11Hz 0.954242 -0.274439
+ 1.315e+11Hz 0.95418 -0.27464
+ 1.316e+11Hz 0.954117 -0.27484
+ 1.317e+11Hz 0.954055 -0.275041
+ 1.318e+11Hz 0.953992 -0.275241
+ 1.319e+11Hz 0.95393 -0.275442
+ 1.32e+11Hz 0.953867 -0.275642
+ 1.321e+11Hz 0.953804 -0.275842
+ 1.322e+11Hz 0.953742 -0.276043
+ 1.323e+11Hz 0.953679 -0.276243
+ 1.324e+11Hz 0.953616 -0.276443
+ 1.325e+11Hz 0.953553 -0.276644
+ 1.326e+11Hz 0.953491 -0.276844
+ 1.327e+11Hz 0.953427 -0.277044
+ 1.328e+11Hz 0.953365 -0.277244
+ 1.329e+11Hz 0.953302 -0.277444
+ 1.33e+11Hz 0.953239 -0.277644
+ 1.331e+11Hz 0.953175 -0.277844
+ 1.332e+11Hz 0.953113 -0.278044
+ 1.333e+11Hz 0.953049 -0.278244
+ 1.334e+11Hz 0.952986 -0.278444
+ 1.335e+11Hz 0.952923 -0.278644
+ 1.336e+11Hz 0.95286 -0.278844
+ 1.337e+11Hz 0.952796 -0.279044
+ 1.338e+11Hz 0.952733 -0.279243
+ 1.339e+11Hz 0.95267 -0.279443
+ 1.34e+11Hz 0.952606 -0.279643
+ 1.341e+11Hz 0.952543 -0.279842
+ 1.342e+11Hz 0.95248 -0.280042
+ 1.343e+11Hz 0.952416 -0.280242
+ 1.344e+11Hz 0.952353 -0.280441
+ 1.345e+11Hz 0.952289 -0.280641
+ 1.346e+11Hz 0.952225 -0.28084
+ 1.347e+11Hz 0.952162 -0.28104
+ 1.348e+11Hz 0.952098 -0.281239
+ 1.349e+11Hz 0.952034 -0.281439
+ 1.35e+11Hz 0.951971 -0.281638
+ 1.351e+11Hz 0.951907 -0.281837
+ 1.352e+11Hz 0.951843 -0.282037
+ 1.353e+11Hz 0.951779 -0.282236
+ 1.354e+11Hz 0.951716 -0.282435
+ 1.355e+11Hz 0.951652 -0.282635
+ 1.356e+11Hz 0.951588 -0.282834
+ 1.357e+11Hz 0.951524 -0.283033
+ 1.358e+11Hz 0.95146 -0.283232
+ 1.359e+11Hz 0.951396 -0.283431
+ 1.36e+11Hz 0.951332 -0.28363
+ 1.361e+11Hz 0.951268 -0.283829
+ 1.362e+11Hz 0.951204 -0.284028
+ 1.363e+11Hz 0.95114 -0.284227
+ 1.364e+11Hz 0.951076 -0.284426
+ 1.365e+11Hz 0.951012 -0.284625
+ 1.366e+11Hz 0.950947 -0.284824
+ 1.367e+11Hz 0.950883 -0.285023
+ 1.368e+11Hz 0.950819 -0.285222
+ 1.369e+11Hz 0.950755 -0.285421
+ 1.37e+11Hz 0.95069 -0.28562
+ 1.371e+11Hz 0.950626 -0.285818
+ 1.372e+11Hz 0.950562 -0.286017
+ 1.373e+11Hz 0.950497 -0.286216
+ 1.374e+11Hz 0.950433 -0.286415
+ 1.375e+11Hz 0.950368 -0.286614
+ 1.376e+11Hz 0.950304 -0.286812
+ 1.377e+11Hz 0.95024 -0.287011
+ 1.378e+11Hz 0.950175 -0.28721
+ 1.379e+11Hz 0.950111 -0.287408
+ 1.38e+11Hz 0.950046 -0.287607
+ 1.381e+11Hz 0.949981 -0.287806
+ 1.382e+11Hz 0.949917 -0.288004
+ 1.383e+11Hz 0.949852 -0.288203
+ 1.384e+11Hz 0.949788 -0.288401
+ 1.385e+11Hz 0.949723 -0.2886
+ 1.386e+11Hz 0.949658 -0.288799
+ 1.387e+11Hz 0.949593 -0.288997
+ 1.388e+11Hz 0.949529 -0.289195
+ 1.389e+11Hz 0.949464 -0.289394
+ 1.39e+11Hz 0.949399 -0.289592
+ 1.391e+11Hz 0.949334 -0.289791
+ 1.392e+11Hz 0.949269 -0.28999
+ 1.393e+11Hz 0.949204 -0.290188
+ 1.394e+11Hz 0.949139 -0.290386
+ 1.395e+11Hz 0.949074 -0.290585
+ 1.396e+11Hz 0.949009 -0.290783
+ 1.397e+11Hz 0.948944 -0.290982
+ 1.398e+11Hz 0.948879 -0.29118
+ 1.399e+11Hz 0.948814 -0.291379
+ 1.4e+11Hz 0.948749 -0.291577
+ 1.401e+11Hz 0.948684 -0.291776
+ 1.402e+11Hz 0.948619 -0.291974
+ 1.403e+11Hz 0.948554 -0.292172
+ 1.404e+11Hz 0.948488 -0.292371
+ 1.405e+11Hz 0.948423 -0.292569
+ 1.406e+11Hz 0.948358 -0.292768
+ 1.407e+11Hz 0.948292 -0.292966
+ 1.408e+11Hz 0.948227 -0.293164
+ 1.409e+11Hz 0.948162 -0.293363
+ 1.41e+11Hz 0.948096 -0.293561
+ 1.411e+11Hz 0.948031 -0.29376
+ 1.412e+11Hz 0.947965 -0.293958
+ 1.413e+11Hz 0.9479 -0.294156
+ 1.414e+11Hz 0.947834 -0.294355
+ 1.415e+11Hz 0.947769 -0.294553
+ 1.416e+11Hz 0.947703 -0.294752
+ 1.417e+11Hz 0.947637 -0.29495
+ 1.418e+11Hz 0.947572 -0.295149
+ 1.419e+11Hz 0.947506 -0.295347
+ 1.42e+11Hz 0.94744 -0.295546
+ 1.421e+11Hz 0.947374 -0.295744
+ 1.422e+11Hz 0.947308 -0.295942
+ 1.423e+11Hz 0.947242 -0.296141
+ 1.424e+11Hz 0.947176 -0.296339
+ 1.425e+11Hz 0.94711 -0.296538
+ 1.426e+11Hz 0.947044 -0.296736
+ 1.427e+11Hz 0.946978 -0.296935
+ 1.428e+11Hz 0.946912 -0.297133
+ 1.429e+11Hz 0.946846 -0.297332
+ 1.43e+11Hz 0.94678 -0.29753
+ 1.431e+11Hz 0.946713 -0.297729
+ 1.432e+11Hz 0.946647 -0.297928
+ 1.433e+11Hz 0.946581 -0.298126
+ 1.434e+11Hz 0.946514 -0.298325
+ 1.435e+11Hz 0.946448 -0.298523
+ 1.436e+11Hz 0.946381 -0.298722
+ 1.437e+11Hz 0.946315 -0.298921
+ 1.438e+11Hz 0.946248 -0.299119
+ 1.439e+11Hz 0.946181 -0.299318
+ 1.44e+11Hz 0.946115 -0.299517
+ 1.441e+11Hz 0.946048 -0.299715
+ 1.442e+11Hz 0.945981 -0.299914
+ 1.443e+11Hz 0.945914 -0.300113
+ 1.444e+11Hz 0.945847 -0.300311
+ 1.445e+11Hz 0.94578 -0.30051
+ 1.446e+11Hz 0.945713 -0.300709
+ 1.447e+11Hz 0.945646 -0.300908
+ 1.448e+11Hz 0.945579 -0.301106
+ 1.449e+11Hz 0.945511 -0.301305
+ 1.45e+11Hz 0.945444 -0.301504
+ 1.451e+11Hz 0.945377 -0.301703
+ 1.452e+11Hz 0.945309 -0.301902
+ 1.453e+11Hz 0.945242 -0.3021
+ 1.454e+11Hz 0.945174 -0.302299
+ 1.455e+11Hz 0.945107 -0.302498
+ 1.456e+11Hz 0.945039 -0.302697
+ 1.457e+11Hz 0.944971 -0.302896
+ 1.458e+11Hz 0.944903 -0.303095
+ 1.459e+11Hz 0.944835 -0.303294
+ 1.46e+11Hz 0.944767 -0.303493
+ 1.461e+11Hz 0.944699 -0.303692
+ 1.462e+11Hz 0.944631 -0.303891
+ 1.463e+11Hz 0.944563 -0.30409
+ 1.464e+11Hz 0.944495 -0.304289
+ 1.465e+11Hz 0.944426 -0.304488
+ 1.466e+11Hz 0.944358 -0.304687
+ 1.467e+11Hz 0.944289 -0.304886
+ 1.468e+11Hz 0.944221 -0.305085
+ 1.469e+11Hz 0.944152 -0.305284
+ 1.47e+11Hz 0.944083 -0.305483
+ 1.471e+11Hz 0.944015 -0.305682
+ 1.472e+11Hz 0.943946 -0.305881
+ 1.473e+11Hz 0.943877 -0.30608
+ 1.474e+11Hz 0.943808 -0.306279
+ 1.475e+11Hz 0.943739 -0.306478
+ 1.476e+11Hz 0.943669 -0.306677
+ 1.477e+11Hz 0.9436 -0.306876
+ 1.478e+11Hz 0.943531 -0.307076
+ 1.479e+11Hz 0.943461 -0.307275
+ 1.48e+11Hz 0.943392 -0.307474
+ 1.481e+11Hz 0.943322 -0.307673
+ 1.482e+11Hz 0.943252 -0.307872
+ 1.483e+11Hz 0.943182 -0.308071
+ 1.484e+11Hz 0.943112 -0.308271
+ 1.485e+11Hz 0.943042 -0.30847
+ 1.486e+11Hz 0.942972 -0.308669
+ 1.487e+11Hz 0.942902 -0.308868
+ 1.488e+11Hz 0.942832 -0.309067
+ 1.489e+11Hz 0.942761 -0.309266
+ 1.49e+11Hz 0.942691 -0.309466
+ 1.491e+11Hz 0.94262 -0.309665
+ 1.492e+11Hz 0.94255 -0.309864
+ 1.493e+11Hz 0.942479 -0.310063
+ 1.494e+11Hz 0.942408 -0.310262
+ 1.495e+11Hz 0.942337 -0.310461
+ 1.496e+11Hz 0.942266 -0.31066
+ 1.497e+11Hz 0.942195 -0.310859
+ 1.498e+11Hz 0.942124 -0.311059
+ 1.499e+11Hz 0.942052 -0.311258
+ 1.5e+11Hz 0.941981 -0.311457
+ ]

A21 %vd(10 3) %vd(21, 22) xfer3
.model xfer3 xfer R_I=true table=[
+ 0Hz 0.99705 0
+ 1e+08Hz 0.99705 -0.000208397
+ 2e+08Hz 0.99705 -0.000416792
+ 3e+08Hz 0.99705 -0.000625183
+ 4e+08Hz 0.997049 -0.000833569
+ 5e+08Hz 0.997049 -0.00104195
+ 6e+08Hz 0.997048 -0.00125032
+ 7e+08Hz 0.997047 -0.00145868
+ 8e+08Hz 0.997046 -0.00166703
+ 9e+08Hz 0.997045 -0.00187536
+ 1e+09Hz 0.997044 -0.00208368
+ 1.1e+09Hz 0.997043 -0.00229198
+ 1.2e+09Hz 0.997041 -0.00250026
+ 1.3e+09Hz 0.997039 -0.00270852
+ 1.4e+09Hz 0.997038 -0.00291676
+ 1.5e+09Hz 0.997036 -0.00312497
+ 1.6e+09Hz 0.997034 -0.00333316
+ 1.7e+09Hz 0.997032 -0.00354133
+ 1.8e+09Hz 0.99703 -0.00374946
+ 1.9e+09Hz 0.997027 -0.00395756
+ 2e+09Hz 0.997025 -0.00416563
+ 2.1e+09Hz 0.997022 -0.00437366
+ 2.2e+09Hz 0.997019 -0.00458166
+ 2.3e+09Hz 0.997016 -0.00478963
+ 2.4e+09Hz 0.997014 -0.00499755
+ 2.5e+09Hz 0.997011 -0.00520544
+ 2.6e+09Hz 0.997007 -0.00541328
+ 2.7e+09Hz 0.997004 -0.00562108
+ 2.8e+09Hz 0.997 -0.00582884
+ 2.9e+09Hz 0.996997 -0.00603655
+ 3e+09Hz 0.996993 -0.00624421
+ 3.1e+09Hz 0.996989 -0.00645182
+ 3.2e+09Hz 0.996986 -0.00665939
+ 3.3e+09Hz 0.996981 -0.0068669
+ 3.4e+09Hz 0.996977 -0.00707436
+ 3.5e+09Hz 0.996973 -0.00728177
+ 3.6e+09Hz 0.996969 -0.00748912
+ 3.7e+09Hz 0.996964 -0.00769641
+ 3.8e+09Hz 0.99696 -0.00790365
+ 3.9e+09Hz 0.996955 -0.00811083
+ 4e+09Hz 0.99695 -0.00831795
+ 4.1e+09Hz 0.996945 -0.008525
+ 4.2e+09Hz 0.99694 -0.008732
+ 4.3e+09Hz 0.996935 -0.00893893
+ 4.4e+09Hz 0.99693 -0.0091458
+ 4.5e+09Hz 0.996925 -0.0093526
+ 4.6e+09Hz 0.996919 -0.00955934
+ 4.7e+09Hz 0.996914 -0.00976601
+ 4.8e+09Hz 0.996908 -0.00997261
+ 4.9e+09Hz 0.996903 -0.0101791
+ 5e+09Hz 0.996897 -0.0103856
+ 5.1e+09Hz 0.996891 -0.010592
+ 5.2e+09Hz 0.996885 -0.0107983
+ 5.3e+09Hz 0.996879 -0.0110046
+ 5.4e+09Hz 0.996873 -0.0112107
+ 5.5e+09Hz 0.996866 -0.0114168
+ 5.6e+09Hz 0.99686 -0.0116229
+ 5.7e+09Hz 0.996854 -0.0118288
+ 5.8e+09Hz 0.996847 -0.0120347
+ 5.9e+09Hz 0.996841 -0.0122405
+ 6e+09Hz 0.996834 -0.0124462
+ 6.1e+09Hz 0.996827 -0.0126519
+ 6.2e+09Hz 0.99682 -0.0128574
+ 6.3e+09Hz 0.996814 -0.0130629
+ 6.4e+09Hz 0.996807 -0.0132683
+ 6.5e+09Hz 0.9968 -0.0134737
+ 6.6e+09Hz 0.996792 -0.0136789
+ 6.7e+09Hz 0.996785 -0.0138841
+ 6.8e+09Hz 0.996778 -0.0140892
+ 6.9e+09Hz 0.996771 -0.0142942
+ 7e+09Hz 0.996763 -0.0144992
+ 7.1e+09Hz 0.996756 -0.014704
+ 7.2e+09Hz 0.996748 -0.0149088
+ 7.3e+09Hz 0.996741 -0.0151135
+ 7.4e+09Hz 0.996733 -0.0153181
+ 7.5e+09Hz 0.996725 -0.0155227
+ 7.6e+09Hz 0.996717 -0.0157271
+ 7.7e+09Hz 0.99671 -0.0159315
+ 7.8e+09Hz 0.996702 -0.0161358
+ 7.9e+09Hz 0.996694 -0.01634
+ 8e+09Hz 0.996686 -0.0165441
+ 8.1e+09Hz 0.996678 -0.0167482
+ 8.2e+09Hz 0.996669 -0.0169521
+ 8.3e+09Hz 0.996661 -0.017156
+ 8.4e+09Hz 0.996653 -0.0173598
+ 8.5e+09Hz 0.996645 -0.0175636
+ 8.6e+09Hz 0.996636 -0.0177672
+ 8.7e+09Hz 0.996628 -0.0179708
+ 8.8e+09Hz 0.99662 -0.0181743
+ 8.9e+09Hz 0.996611 -0.0183777
+ 9e+09Hz 0.996603 -0.0185811
+ 9.1e+09Hz 0.996594 -0.0187843
+ 9.2e+09Hz 0.996586 -0.0189875
+ 9.3e+09Hz 0.996577 -0.0191906
+ 9.4e+09Hz 0.996568 -0.0193936
+ 9.5e+09Hz 0.99656 -0.0195966
+ 9.6e+09Hz 0.996551 -0.0197995
+ 9.7e+09Hz 0.996542 -0.0200023
+ 9.8e+09Hz 0.996533 -0.020205
+ 9.9e+09Hz 0.996524 -0.0204077
+ 1e+10Hz 0.996515 -0.0206103
+ 1.01e+10Hz 0.996506 -0.0208128
+ 1.02e+10Hz 0.996498 -0.0210152
+ 1.03e+10Hz 0.996488 -0.0212176
+ 1.04e+10Hz 0.996479 -0.0214199
+ 1.05e+10Hz 0.99647 -0.0216221
+ 1.06e+10Hz 0.996461 -0.0218242
+ 1.07e+10Hz 0.996452 -0.0220263
+ 1.08e+10Hz 0.996443 -0.0222284
+ 1.09e+10Hz 0.996434 -0.0224303
+ 1.1e+10Hz 0.996425 -0.0226322
+ 1.11e+10Hz 0.996416 -0.022834
+ 1.12e+10Hz 0.996406 -0.0230358
+ 1.13e+10Hz 0.996397 -0.0232375
+ 1.14e+10Hz 0.996388 -0.0234391
+ 1.15e+10Hz 0.996379 -0.0236407
+ 1.16e+10Hz 0.996369 -0.0238422
+ 1.17e+10Hz 0.99636 -0.0240436
+ 1.18e+10Hz 0.996351 -0.024245
+ 1.19e+10Hz 0.996341 -0.0244463
+ 1.2e+10Hz 0.996332 -0.0246476
+ 1.21e+10Hz 0.996322 -0.0248488
+ 1.22e+10Hz 0.996313 -0.02505
+ 1.23e+10Hz 0.996304 -0.0252511
+ 1.24e+10Hz 0.996294 -0.0254521
+ 1.25e+10Hz 0.996285 -0.0256531
+ 1.26e+10Hz 0.996275 -0.025854
+ 1.27e+10Hz 0.996266 -0.0260549
+ 1.28e+10Hz 0.996256 -0.0262558
+ 1.29e+10Hz 0.996247 -0.0264565
+ 1.3e+10Hz 0.996237 -0.0266573
+ 1.31e+10Hz 0.996228 -0.026858
+ 1.32e+10Hz 0.996218 -0.0270586
+ 1.33e+10Hz 0.996209 -0.0272592
+ 1.34e+10Hz 0.996199 -0.0274597
+ 1.35e+10Hz 0.996189 -0.0276603
+ 1.36e+10Hz 0.99618 -0.0278607
+ 1.37e+10Hz 0.99617 -0.0280611
+ 1.38e+10Hz 0.996161 -0.0282615
+ 1.39e+10Hz 0.996151 -0.0284618
+ 1.4e+10Hz 0.996141 -0.0286621
+ 1.41e+10Hz 0.996132 -0.0288624
+ 1.42e+10Hz 0.996122 -0.0290626
+ 1.43e+10Hz 0.996112 -0.0292628
+ 1.44e+10Hz 0.996103 -0.0294629
+ 1.45e+10Hz 0.996093 -0.029663
+ 1.46e+10Hz 0.996083 -0.0298631
+ 1.47e+10Hz 0.996073 -0.0300632
+ 1.48e+10Hz 0.996064 -0.0302631
+ 1.49e+10Hz 0.996054 -0.0304631
+ 1.5e+10Hz 0.996044 -0.0306631
+ 1.51e+10Hz 0.996035 -0.030863
+ 1.52e+10Hz 0.996025 -0.0310629
+ 1.53e+10Hz 0.996015 -0.0312627
+ 1.54e+10Hz 0.996005 -0.0314626
+ 1.55e+10Hz 0.995995 -0.0316624
+ 1.56e+10Hz 0.995986 -0.0318622
+ 1.57e+10Hz 0.995976 -0.0320619
+ 1.58e+10Hz 0.995966 -0.0322617
+ 1.59e+10Hz 0.995956 -0.0324614
+ 1.6e+10Hz 0.995946 -0.032661
+ 1.61e+10Hz 0.995937 -0.0328607
+ 1.62e+10Hz 0.995927 -0.0330604
+ 1.63e+10Hz 0.995917 -0.03326
+ 1.64e+10Hz 0.995907 -0.0334596
+ 1.65e+10Hz 0.995897 -0.0336592
+ 1.66e+10Hz 0.995887 -0.0338587
+ 1.67e+10Hz 0.995877 -0.0340583
+ 1.68e+10Hz 0.995867 -0.0342578
+ 1.69e+10Hz 0.995857 -0.0344574
+ 1.7e+10Hz 0.995847 -0.0346569
+ 1.71e+10Hz 0.995837 -0.0348564
+ 1.72e+10Hz 0.995827 -0.0350558
+ 1.73e+10Hz 0.995817 -0.0352553
+ 1.74e+10Hz 0.995807 -0.0354548
+ 1.75e+10Hz 0.995797 -0.0356542
+ 1.76e+10Hz 0.995787 -0.0358537
+ 1.77e+10Hz 0.995777 -0.0360531
+ 1.78e+10Hz 0.995767 -0.0362525
+ 1.79e+10Hz 0.995757 -0.0364519
+ 1.8e+10Hz 0.995747 -0.0366513
+ 1.81e+10Hz 0.995737 -0.0368507
+ 1.82e+10Hz 0.995727 -0.0370501
+ 1.83e+10Hz 0.995717 -0.0372495
+ 1.84e+10Hz 0.995707 -0.0374489
+ 1.85e+10Hz 0.995696 -0.0376483
+ 1.86e+10Hz 0.995686 -0.0378476
+ 1.87e+10Hz 0.995676 -0.038047
+ 1.88e+10Hz 0.995666 -0.0382464
+ 1.89e+10Hz 0.995656 -0.0384457
+ 1.9e+10Hz 0.995645 -0.0386451
+ 1.91e+10Hz 0.995635 -0.0388445
+ 1.92e+10Hz 0.995625 -0.0390438
+ 1.93e+10Hz 0.995614 -0.0392432
+ 1.94e+10Hz 0.995604 -0.0394425
+ 1.95e+10Hz 0.995594 -0.0396419
+ 1.96e+10Hz 0.995583 -0.0398412
+ 1.97e+10Hz 0.995573 -0.0400406
+ 1.98e+10Hz 0.995563 -0.0402399
+ 1.99e+10Hz 0.995552 -0.0404393
+ 2e+10Hz 0.995542 -0.0406387
+ 2.01e+10Hz 0.995531 -0.040838
+ 2.02e+10Hz 0.995521 -0.0410374
+ 2.03e+10Hz 0.99551 -0.0412368
+ 2.04e+10Hz 0.995499 -0.0414361
+ 2.05e+10Hz 0.995489 -0.0416355
+ 2.06e+10Hz 0.995478 -0.0418349
+ 2.07e+10Hz 0.995467 -0.0420343
+ 2.08e+10Hz 0.995457 -0.0422337
+ 2.09e+10Hz 0.995446 -0.0424331
+ 2.1e+10Hz 0.995435 -0.0426325
+ 2.11e+10Hz 0.995425 -0.0428319
+ 2.12e+10Hz 0.995414 -0.0430313
+ 2.13e+10Hz 0.995403 -0.0432307
+ 2.14e+10Hz 0.995392 -0.0434302
+ 2.15e+10Hz 0.995381 -0.0436296
+ 2.16e+10Hz 0.99537 -0.043829
+ 2.17e+10Hz 0.995359 -0.0440285
+ 2.18e+10Hz 0.995348 -0.0442279
+ 2.19e+10Hz 0.995337 -0.0444274
+ 2.2e+10Hz 0.995326 -0.0446268
+ 2.21e+10Hz 0.995315 -0.0448263
+ 2.22e+10Hz 0.995304 -0.0450258
+ 2.23e+10Hz 0.995293 -0.0452253
+ 2.24e+10Hz 0.995282 -0.0454248
+ 2.25e+10Hz 0.995271 -0.0456243
+ 2.26e+10Hz 0.995259 -0.0458238
+ 2.27e+10Hz 0.995248 -0.0460233
+ 2.28e+10Hz 0.995237 -0.0462228
+ 2.29e+10Hz 0.995225 -0.0464223
+ 2.3e+10Hz 0.995214 -0.0466219
+ 2.31e+10Hz 0.995203 -0.0468214
+ 2.32e+10Hz 0.995191 -0.047021
+ 2.33e+10Hz 0.99518 -0.0472205
+ 2.34e+10Hz 0.995168 -0.0474201
+ 2.35e+10Hz 0.995156 -0.0476197
+ 2.36e+10Hz 0.995145 -0.0478193
+ 2.37e+10Hz 0.995133 -0.0480189
+ 2.38e+10Hz 0.995121 -0.0482185
+ 2.39e+10Hz 0.99511 -0.0484181
+ 2.4e+10Hz 0.995098 -0.0486177
+ 2.41e+10Hz 0.995086 -0.0488173
+ 2.42e+10Hz 0.995074 -0.0490169
+ 2.43e+10Hz 0.995062 -0.0492166
+ 2.44e+10Hz 0.99505 -0.0494162
+ 2.45e+10Hz 0.995038 -0.0496159
+ 2.46e+10Hz 0.995026 -0.0498155
+ 2.47e+10Hz 0.995014 -0.0500152
+ 2.48e+10Hz 0.995002 -0.0502149
+ 2.49e+10Hz 0.99499 -0.0504145
+ 2.5e+10Hz 0.994978 -0.0506142
+ 2.51e+10Hz 0.994966 -0.0508139
+ 2.52e+10Hz 0.994953 -0.0510136
+ 2.53e+10Hz 0.994941 -0.0512133
+ 2.54e+10Hz 0.994929 -0.051413
+ 2.55e+10Hz 0.994916 -0.0516127
+ 2.56e+10Hz 0.994904 -0.0518125
+ 2.57e+10Hz 0.994891 -0.0520122
+ 2.58e+10Hz 0.994879 -0.0522119
+ 2.59e+10Hz 0.994866 -0.0524117
+ 2.6e+10Hz 0.994853 -0.0526114
+ 2.61e+10Hz 0.994841 -0.0528112
+ 2.62e+10Hz 0.994828 -0.0530109
+ 2.63e+10Hz 0.994815 -0.0532107
+ 2.64e+10Hz 0.994802 -0.0534104
+ 2.65e+10Hz 0.994789 -0.0536102
+ 2.66e+10Hz 0.994776 -0.05381
+ 2.67e+10Hz 0.994764 -0.0540097
+ 2.68e+10Hz 0.99475 -0.0542095
+ 2.69e+10Hz 0.994737 -0.0544093
+ 2.7e+10Hz 0.994724 -0.0546091
+ 2.71e+10Hz 0.994711 -0.0548088
+ 2.72e+10Hz 0.994698 -0.0550086
+ 2.73e+10Hz 0.994685 -0.0552084
+ 2.74e+10Hz 0.994671 -0.0554082
+ 2.75e+10Hz 0.994658 -0.055608
+ 2.76e+10Hz 0.994645 -0.0558078
+ 2.77e+10Hz 0.994631 -0.0560076
+ 2.78e+10Hz 0.994618 -0.0562074
+ 2.79e+10Hz 0.994604 -0.0564072
+ 2.8e+10Hz 0.99459 -0.056607
+ 2.81e+10Hz 0.994577 -0.0568068
+ 2.82e+10Hz 0.994563 -0.0570066
+ 2.83e+10Hz 0.994549 -0.0572064
+ 2.84e+10Hz 0.994535 -0.0574062
+ 2.85e+10Hz 0.994521 -0.057606
+ 2.86e+10Hz 0.994508 -0.0578058
+ 2.87e+10Hz 0.994494 -0.0580056
+ 2.88e+10Hz 0.99448 -0.0582054
+ 2.89e+10Hz 0.994466 -0.0584052
+ 2.9e+10Hz 0.994452 -0.058605
+ 2.91e+10Hz 0.994437 -0.0588048
+ 2.92e+10Hz 0.994423 -0.0590046
+ 2.93e+10Hz 0.994409 -0.0592044
+ 2.94e+10Hz 0.994395 -0.0594042
+ 2.95e+10Hz 0.99438 -0.059604
+ 2.96e+10Hz 0.994366 -0.0598038
+ 2.97e+10Hz 0.994352 -0.0600036
+ 2.98e+10Hz 0.994337 -0.0602033
+ 2.99e+10Hz 0.994322 -0.0604031
+ 3e+10Hz 0.994308 -0.0606029
+ 3.01e+10Hz 0.994293 -0.0608027
+ 3.02e+10Hz 0.994278 -0.0610024
+ 3.03e+10Hz 0.994264 -0.0612022
+ 3.04e+10Hz 0.994249 -0.0614019
+ 3.05e+10Hz 0.994234 -0.0616017
+ 3.06e+10Hz 0.994219 -0.0618014
+ 3.07e+10Hz 0.994204 -0.0620012
+ 3.08e+10Hz 0.994189 -0.0622009
+ 3.09e+10Hz 0.994174 -0.0624007
+ 3.1e+10Hz 0.994159 -0.0626004
+ 3.11e+10Hz 0.994144 -0.0628001
+ 3.12e+10Hz 0.994129 -0.0629998
+ 3.13e+10Hz 0.994114 -0.0631995
+ 3.14e+10Hz 0.994098 -0.0633992
+ 3.15e+10Hz 0.994083 -0.0635989
+ 3.16e+10Hz 0.994068 -0.0637986
+ 3.17e+10Hz 0.994052 -0.0639983
+ 3.18e+10Hz 0.994037 -0.064198
+ 3.19e+10Hz 0.994021 -0.0643977
+ 3.2e+10Hz 0.994006 -0.0645973
+ 3.21e+10Hz 0.99399 -0.064797
+ 3.22e+10Hz 0.993975 -0.0649966
+ 3.23e+10Hz 0.993959 -0.0651963
+ 3.24e+10Hz 0.993943 -0.0653959
+ 3.25e+10Hz 0.993927 -0.0655955
+ 3.26e+10Hz 0.993912 -0.0657951
+ 3.27e+10Hz 0.993896 -0.0659948
+ 3.28e+10Hz 0.99388 -0.0661943
+ 3.29e+10Hz 0.993864 -0.0663939
+ 3.3e+10Hz 0.993848 -0.0665935
+ 3.31e+10Hz 0.993832 -0.0667931
+ 3.32e+10Hz 0.993816 -0.0669927
+ 3.33e+10Hz 0.993799 -0.0671922
+ 3.34e+10Hz 0.993783 -0.0673918
+ 3.35e+10Hz 0.993767 -0.0675913
+ 3.36e+10Hz 0.993751 -0.0677908
+ 3.37e+10Hz 0.993734 -0.0679904
+ 3.38e+10Hz 0.993718 -0.0681899
+ 3.39e+10Hz 0.993702 -0.0683894
+ 3.4e+10Hz 0.993685 -0.0685889
+ 3.41e+10Hz 0.993669 -0.0687884
+ 3.42e+10Hz 0.993652 -0.0689878
+ 3.43e+10Hz 0.993636 -0.0691873
+ 3.44e+10Hz 0.993619 -0.0693868
+ 3.45e+10Hz 0.993602 -0.0695862
+ 3.46e+10Hz 0.993586 -0.0697856
+ 3.47e+10Hz 0.993569 -0.0699851
+ 3.48e+10Hz 0.993552 -0.0701845
+ 3.49e+10Hz 0.993535 -0.0703839
+ 3.5e+10Hz 0.993518 -0.0705833
+ 3.51e+10Hz 0.993501 -0.0707827
+ 3.52e+10Hz 0.993484 -0.070982
+ 3.53e+10Hz 0.993467 -0.0711814
+ 3.54e+10Hz 0.99345 -0.0713808
+ 3.55e+10Hz 0.993433 -0.0715801
+ 3.56e+10Hz 0.993416 -0.0717794
+ 3.57e+10Hz 0.993399 -0.0719787
+ 3.58e+10Hz 0.993382 -0.0721781
+ 3.59e+10Hz 0.993364 -0.0723774
+ 3.6e+10Hz 0.993347 -0.0725767
+ 3.61e+10Hz 0.99333 -0.0727759
+ 3.62e+10Hz 0.993312 -0.0729752
+ 3.63e+10Hz 0.993295 -0.0731745
+ 3.64e+10Hz 0.993278 -0.0733737
+ 3.65e+10Hz 0.99326 -0.073573
+ 3.66e+10Hz 0.993243 -0.0737722
+ 3.67e+10Hz 0.993225 -0.0739714
+ 3.68e+10Hz 0.993207 -0.0741706
+ 3.69e+10Hz 0.99319 -0.0743698
+ 3.7e+10Hz 0.993172 -0.074569
+ 3.71e+10Hz 0.993154 -0.0747682
+ 3.72e+10Hz 0.993136 -0.0749674
+ 3.73e+10Hz 0.993119 -0.0751665
+ 3.74e+10Hz 0.993101 -0.0753657
+ 3.75e+10Hz 0.993083 -0.0755648
+ 3.76e+10Hz 0.993065 -0.0757639
+ 3.77e+10Hz 0.993047 -0.0759631
+ 3.78e+10Hz 0.993029 -0.0761622
+ 3.79e+10Hz 0.993011 -0.0763613
+ 3.8e+10Hz 0.992993 -0.0765604
+ 3.81e+10Hz 0.992975 -0.0767594
+ 3.82e+10Hz 0.992957 -0.0769585
+ 3.83e+10Hz 0.992939 -0.0771576
+ 3.84e+10Hz 0.99292 -0.0773566
+ 3.85e+10Hz 0.992902 -0.0775557
+ 3.86e+10Hz 0.992884 -0.0777547
+ 3.87e+10Hz 0.992866 -0.0779537
+ 3.88e+10Hz 0.992847 -0.0781527
+ 3.89e+10Hz 0.992829 -0.0783517
+ 3.9e+10Hz 0.99281 -0.0785507
+ 3.91e+10Hz 0.992792 -0.0787497
+ 3.92e+10Hz 0.992773 -0.0789487
+ 3.93e+10Hz 0.992755 -0.0791477
+ 3.94e+10Hz 0.992736 -0.0793466
+ 3.95e+10Hz 0.992718 -0.0795456
+ 3.96e+10Hz 0.992699 -0.0797445
+ 3.97e+10Hz 0.99268 -0.0799435
+ 3.98e+10Hz 0.992662 -0.0801424
+ 3.99e+10Hz 0.992643 -0.0803413
+ 4e+10Hz 0.992624 -0.0805402
+ 4.01e+10Hz 0.992605 -0.0807391
+ 4.02e+10Hz 0.992587 -0.080938
+ 4.03e+10Hz 0.992568 -0.0811369
+ 4.04e+10Hz 0.992549 -0.0813358
+ 4.05e+10Hz 0.99253 -0.0815347
+ 4.06e+10Hz 0.992511 -0.0817335
+ 4.07e+10Hz 0.992492 -0.0819324
+ 4.08e+10Hz 0.992473 -0.0821312
+ 4.09e+10Hz 0.992454 -0.0823301
+ 4.1e+10Hz 0.992435 -0.0825289
+ 4.11e+10Hz 0.992416 -0.0827277
+ 4.12e+10Hz 0.992396 -0.0829266
+ 4.13e+10Hz 0.992377 -0.0831254
+ 4.14e+10Hz 0.992358 -0.0833242
+ 4.15e+10Hz 0.992339 -0.083523
+ 4.16e+10Hz 0.992319 -0.0837218
+ 4.17e+10Hz 0.9923 -0.0839206
+ 4.18e+10Hz 0.992281 -0.0841194
+ 4.19e+10Hz 0.992261 -0.0843181
+ 4.2e+10Hz 0.992242 -0.0845169
+ 4.21e+10Hz 0.992222 -0.0847157
+ 4.22e+10Hz 0.992203 -0.0849144
+ 4.23e+10Hz 0.992183 -0.0851132
+ 4.24e+10Hz 0.992163 -0.0853119
+ 4.25e+10Hz 0.992144 -0.0855107
+ 4.26e+10Hz 0.992124 -0.0857094
+ 4.27e+10Hz 0.992105 -0.0859082
+ 4.28e+10Hz 0.992085 -0.0861069
+ 4.29e+10Hz 0.992065 -0.0863056
+ 4.3e+10Hz 0.992045 -0.0865043
+ 4.31e+10Hz 0.992026 -0.086703
+ 4.32e+10Hz 0.992006 -0.0869017
+ 4.33e+10Hz 0.991986 -0.0871004
+ 4.34e+10Hz 0.991966 -0.0872992
+ 4.35e+10Hz 0.991946 -0.0874979
+ 4.36e+10Hz 0.991926 -0.0876965
+ 4.37e+10Hz 0.991906 -0.0878952
+ 4.38e+10Hz 0.991886 -0.0880939
+ 4.39e+10Hz 0.991866 -0.0882926
+ 4.4e+10Hz 0.991846 -0.0884913
+ 4.41e+10Hz 0.991826 -0.0886899
+ 4.42e+10Hz 0.991805 -0.0888886
+ 4.43e+10Hz 0.991785 -0.0890873
+ 4.44e+10Hz 0.991765 -0.0892859
+ 4.45e+10Hz 0.991745 -0.0894846
+ 4.46e+10Hz 0.991724 -0.0896833
+ 4.47e+10Hz 0.991704 -0.0898819
+ 4.48e+10Hz 0.991684 -0.0900806
+ 4.49e+10Hz 0.991663 -0.0902792
+ 4.5e+10Hz 0.991643 -0.0904778
+ 4.51e+10Hz 0.991622 -0.0906765
+ 4.52e+10Hz 0.991602 -0.0908751
+ 4.53e+10Hz 0.991581 -0.0910738
+ 4.54e+10Hz 0.991561 -0.0912724
+ 4.55e+10Hz 0.99154 -0.091471
+ 4.56e+10Hz 0.991519 -0.0916697
+ 4.57e+10Hz 0.991499 -0.0918683
+ 4.58e+10Hz 0.991478 -0.0920669
+ 4.59e+10Hz 0.991457 -0.0922655
+ 4.6e+10Hz 0.991436 -0.0924642
+ 4.61e+10Hz 0.991416 -0.0926628
+ 4.62e+10Hz 0.991395 -0.0928614
+ 4.63e+10Hz 0.991374 -0.09306
+ 4.64e+10Hz 0.991353 -0.0932586
+ 4.65e+10Hz 0.991332 -0.0934572
+ 4.66e+10Hz 0.991311 -0.0936558
+ 4.67e+10Hz 0.99129 -0.0938545
+ 4.68e+10Hz 0.991269 -0.0940531
+ 4.69e+10Hz 0.991248 -0.0942517
+ 4.7e+10Hz 0.991227 -0.0944503
+ 4.71e+10Hz 0.991205 -0.0946489
+ 4.72e+10Hz 0.991184 -0.0948475
+ 4.73e+10Hz 0.991163 -0.0950461
+ 4.74e+10Hz 0.991142 -0.0952447
+ 4.75e+10Hz 0.99112 -0.0954433
+ 4.76e+10Hz 0.991099 -0.0956419
+ 4.77e+10Hz 0.991078 -0.0958405
+ 4.78e+10Hz 0.991056 -0.0960391
+ 4.79e+10Hz 0.991035 -0.0962376
+ 4.8e+10Hz 0.991013 -0.0964362
+ 4.81e+10Hz 0.990992 -0.0966348
+ 4.82e+10Hz 0.99097 -0.0968334
+ 4.83e+10Hz 0.990949 -0.097032
+ 4.84e+10Hz 0.990927 -0.0972306
+ 4.85e+10Hz 0.990905 -0.0974292
+ 4.86e+10Hz 0.990884 -0.0976278
+ 4.87e+10Hz 0.990862 -0.0978264
+ 4.88e+10Hz 0.99084 -0.0980249
+ 4.89e+10Hz 0.990818 -0.0982235
+ 4.9e+10Hz 0.990796 -0.0984221
+ 4.91e+10Hz 0.990774 -0.0986207
+ 4.92e+10Hz 0.990753 -0.0988193
+ 4.93e+10Hz 0.99073 -0.0990178
+ 4.94e+10Hz 0.990708 -0.0992164
+ 4.95e+10Hz 0.990686 -0.099415
+ 4.96e+10Hz 0.990664 -0.0996136
+ 4.97e+10Hz 0.990642 -0.0998121
+ 4.98e+10Hz 0.99062 -0.100011
+ 4.99e+10Hz 0.990598 -0.100209
+ 5e+10Hz 0.990576 -0.100408
+ 5.01e+10Hz 0.990553 -0.100606
+ 5.02e+10Hz 0.990531 -0.100805
+ 5.03e+10Hz 0.990509 -0.101004
+ 5.04e+10Hz 0.990486 -0.101202
+ 5.05e+10Hz 0.990464 -0.101401
+ 5.06e+10Hz 0.990441 -0.101599
+ 5.07e+10Hz 0.990419 -0.101798
+ 5.08e+10Hz 0.990396 -0.101996
+ 5.09e+10Hz 0.990374 -0.102195
+ 5.1e+10Hz 0.990351 -0.102393
+ 5.11e+10Hz 0.990328 -0.102592
+ 5.12e+10Hz 0.990306 -0.102791
+ 5.13e+10Hz 0.990283 -0.102989
+ 5.14e+10Hz 0.99026 -0.103188
+ 5.15e+10Hz 0.990237 -0.103386
+ 5.16e+10Hz 0.990214 -0.103585
+ 5.17e+10Hz 0.990192 -0.103783
+ 5.18e+10Hz 0.990169 -0.103982
+ 5.19e+10Hz 0.990146 -0.10418
+ 5.2e+10Hz 0.990123 -0.104379
+ 5.21e+10Hz 0.990099 -0.104578
+ 5.22e+10Hz 0.990076 -0.104776
+ 5.23e+10Hz 0.990053 -0.104975
+ 5.24e+10Hz 0.99003 -0.105173
+ 5.25e+10Hz 0.990007 -0.105372
+ 5.26e+10Hz 0.989984 -0.10557
+ 5.27e+10Hz 0.98996 -0.105769
+ 5.28e+10Hz 0.989937 -0.105967
+ 5.29e+10Hz 0.989913 -0.106166
+ 5.3e+10Hz 0.98989 -0.106364
+ 5.31e+10Hz 0.989866 -0.106563
+ 5.32e+10Hz 0.989843 -0.106761
+ 5.33e+10Hz 0.989819 -0.10696
+ 5.34e+10Hz 0.989796 -0.107158
+ 5.35e+10Hz 0.989772 -0.107357
+ 5.36e+10Hz 0.989748 -0.107555
+ 5.37e+10Hz 0.989725 -0.107754
+ 5.38e+10Hz 0.989701 -0.107952
+ 5.39e+10Hz 0.989677 -0.108151
+ 5.4e+10Hz 0.989653 -0.108349
+ 5.41e+10Hz 0.989629 -0.108548
+ 5.42e+10Hz 0.989605 -0.108746
+ 5.43e+10Hz 0.989581 -0.108945
+ 5.44e+10Hz 0.989557 -0.109143
+ 5.45e+10Hz 0.989533 -0.109342
+ 5.46e+10Hz 0.989509 -0.10954
+ 5.47e+10Hz 0.989485 -0.109739
+ 5.48e+10Hz 0.989461 -0.109937
+ 5.49e+10Hz 0.989437 -0.110135
+ 5.5e+10Hz 0.989412 -0.110334
+ 5.51e+10Hz 0.989388 -0.110532
+ 5.52e+10Hz 0.989363 -0.110731
+ 5.53e+10Hz 0.989339 -0.110929
+ 5.54e+10Hz 0.989315 -0.111128
+ 5.55e+10Hz 0.98929 -0.111326
+ 5.56e+10Hz 0.989266 -0.111525
+ 5.57e+10Hz 0.989241 -0.111723
+ 5.58e+10Hz 0.989216 -0.111921
+ 5.59e+10Hz 0.989192 -0.11212
+ 5.6e+10Hz 0.989167 -0.112318
+ 5.61e+10Hz 0.989142 -0.112517
+ 5.62e+10Hz 0.989117 -0.112715
+ 5.63e+10Hz 0.989093 -0.112913
+ 5.64e+10Hz 0.989068 -0.113112
+ 5.65e+10Hz 0.989043 -0.11331
+ 5.66e+10Hz 0.989018 -0.113508
+ 5.67e+10Hz 0.988993 -0.113707
+ 5.68e+10Hz 0.988968 -0.113905
+ 5.69e+10Hz 0.988942 -0.114103
+ 5.7e+10Hz 0.988917 -0.114302
+ 5.71e+10Hz 0.988892 -0.1145
+ 5.72e+10Hz 0.988867 -0.114698
+ 5.73e+10Hz 0.988842 -0.114897
+ 5.74e+10Hz 0.988816 -0.115095
+ 5.75e+10Hz 0.988791 -0.115293
+ 5.76e+10Hz 0.988765 -0.115492
+ 5.77e+10Hz 0.98874 -0.11569
+ 5.78e+10Hz 0.988715 -0.115888
+ 5.79e+10Hz 0.988689 -0.116086
+ 5.8e+10Hz 0.988663 -0.116285
+ 5.81e+10Hz 0.988638 -0.116483
+ 5.82e+10Hz 0.988612 -0.116681
+ 5.83e+10Hz 0.988586 -0.116879
+ 5.84e+10Hz 0.988561 -0.117078
+ 5.85e+10Hz 0.988535 -0.117276
+ 5.86e+10Hz 0.988509 -0.117474
+ 5.87e+10Hz 0.988483 -0.117672
+ 5.88e+10Hz 0.988457 -0.117871
+ 5.89e+10Hz 0.988431 -0.118069
+ 5.9e+10Hz 0.988405 -0.118267
+ 5.91e+10Hz 0.988379 -0.118465
+ 5.92e+10Hz 0.988353 -0.118663
+ 5.93e+10Hz 0.988327 -0.118861
+ 5.94e+10Hz 0.988301 -0.11906
+ 5.95e+10Hz 0.988274 -0.119258
+ 5.96e+10Hz 0.988248 -0.119456
+ 5.97e+10Hz 0.988222 -0.119654
+ 5.98e+10Hz 0.988195 -0.119852
+ 5.99e+10Hz 0.988169 -0.12005
+ 6e+10Hz 0.988143 -0.120248
+ 6.01e+10Hz 0.988116 -0.120446
+ 6.02e+10Hz 0.988089 -0.120644
+ 6.03e+10Hz 0.988063 -0.120843
+ 6.04e+10Hz 0.988036 -0.12104
+ 6.05e+10Hz 0.988009 -0.121239
+ 6.06e+10Hz 0.987983 -0.121437
+ 6.07e+10Hz 0.987956 -0.121635
+ 6.08e+10Hz 0.987929 -0.121833
+ 6.09e+10Hz 0.987902 -0.122031
+ 6.1e+10Hz 0.987876 -0.122229
+ 6.11e+10Hz 0.987849 -0.122427
+ 6.12e+10Hz 0.987822 -0.122625
+ 6.13e+10Hz 0.987795 -0.122823
+ 6.14e+10Hz 0.987768 -0.123021
+ 6.15e+10Hz 0.98774 -0.123218
+ 6.16e+10Hz 0.987713 -0.123416
+ 6.17e+10Hz 0.987686 -0.123614
+ 6.18e+10Hz 0.987659 -0.123812
+ 6.19e+10Hz 0.987632 -0.12401
+ 6.2e+10Hz 0.987604 -0.124208
+ 6.21e+10Hz 0.987577 -0.124406
+ 6.22e+10Hz 0.98755 -0.124604
+ 6.23e+10Hz 0.987522 -0.124801
+ 6.24e+10Hz 0.987495 -0.124999
+ 6.25e+10Hz 0.987467 -0.125197
+ 6.26e+10Hz 0.98744 -0.125395
+ 6.27e+10Hz 0.987412 -0.125593
+ 6.28e+10Hz 0.987384 -0.125791
+ 6.29e+10Hz 0.987357 -0.125988
+ 6.3e+10Hz 0.987329 -0.126186
+ 6.31e+10Hz 0.987301 -0.126384
+ 6.32e+10Hz 0.987273 -0.126582
+ 6.33e+10Hz 0.987245 -0.126779
+ 6.34e+10Hz 0.987217 -0.126977
+ 6.35e+10Hz 0.98719 -0.127175
+ 6.36e+10Hz 0.987162 -0.127373
+ 6.37e+10Hz 0.987134 -0.12757
+ 6.38e+10Hz 0.987105 -0.127768
+ 6.39e+10Hz 0.987077 -0.127966
+ 6.4e+10Hz 0.987049 -0.128163
+ 6.41e+10Hz 0.987021 -0.128361
+ 6.42e+10Hz 0.986993 -0.128559
+ 6.43e+10Hz 0.986965 -0.128756
+ 6.44e+10Hz 0.986936 -0.128954
+ 6.45e+10Hz 0.986908 -0.129151
+ 6.46e+10Hz 0.98688 -0.129349
+ 6.47e+10Hz 0.986851 -0.129547
+ 6.48e+10Hz 0.986823 -0.129744
+ 6.49e+10Hz 0.986794 -0.129942
+ 6.5e+10Hz 0.986766 -0.130139
+ 6.51e+10Hz 0.986737 -0.130337
+ 6.52e+10Hz 0.986708 -0.130534
+ 6.53e+10Hz 0.98668 -0.130732
+ 6.54e+10Hz 0.986651 -0.130929
+ 6.55e+10Hz 0.986622 -0.131127
+ 6.56e+10Hz 0.986594 -0.131324
+ 6.57e+10Hz 0.986565 -0.131522
+ 6.58e+10Hz 0.986536 -0.131719
+ 6.59e+10Hz 0.986507 -0.131916
+ 6.6e+10Hz 0.986478 -0.132114
+ 6.61e+10Hz 0.986449 -0.132311
+ 6.62e+10Hz 0.98642 -0.132509
+ 6.63e+10Hz 0.986391 -0.132706
+ 6.64e+10Hz 0.986362 -0.132904
+ 6.65e+10Hz 0.986333 -0.133101
+ 6.66e+10Hz 0.986303 -0.133298
+ 6.67e+10Hz 0.986274 -0.133496
+ 6.68e+10Hz 0.986245 -0.133693
+ 6.69e+10Hz 0.986216 -0.13389
+ 6.7e+10Hz 0.986186 -0.134088
+ 6.71e+10Hz 0.986157 -0.134285
+ 6.72e+10Hz 0.986128 -0.134482
+ 6.73e+10Hz 0.986098 -0.134679
+ 6.74e+10Hz 0.986069 -0.134877
+ 6.75e+10Hz 0.986039 -0.135074
+ 6.76e+10Hz 0.986009 -0.135271
+ 6.77e+10Hz 0.98598 -0.135468
+ 6.78e+10Hz 0.98595 -0.135666
+ 6.79e+10Hz 0.98592 -0.135863
+ 6.8e+10Hz 0.985891 -0.13606
+ 6.81e+10Hz 0.985861 -0.136257
+ 6.82e+10Hz 0.985831 -0.136454
+ 6.83e+10Hz 0.985801 -0.136652
+ 6.84e+10Hz 0.985771 -0.136849
+ 6.85e+10Hz 0.985742 -0.137046
+ 6.86e+10Hz 0.985711 -0.137243
+ 6.87e+10Hz 0.985681 -0.13744
+ 6.88e+10Hz 0.985652 -0.137637
+ 6.89e+10Hz 0.985621 -0.137834
+ 6.9e+10Hz 0.985591 -0.138031
+ 6.91e+10Hz 0.985561 -0.138229
+ 6.92e+10Hz 0.985531 -0.138426
+ 6.93e+10Hz 0.985501 -0.138623
+ 6.94e+10Hz 0.985471 -0.13882
+ 6.95e+10Hz 0.98544 -0.139017
+ 6.96e+10Hz 0.98541 -0.139214
+ 6.97e+10Hz 0.985379 -0.139411
+ 6.98e+10Hz 0.985349 -0.139608
+ 6.99e+10Hz 0.985318 -0.139805
+ 7e+10Hz 0.985288 -0.140002
+ 7.01e+10Hz 0.985258 -0.140199
+ 7.02e+10Hz 0.985227 -0.140396
+ 7.03e+10Hz 0.985196 -0.140593
+ 7.04e+10Hz 0.985166 -0.14079
+ 7.05e+10Hz 0.985135 -0.140986
+ 7.06e+10Hz 0.985104 -0.141183
+ 7.07e+10Hz 0.985074 -0.14138
+ 7.08e+10Hz 0.985043 -0.141577
+ 7.09e+10Hz 0.985012 -0.141774
+ 7.1e+10Hz 0.984981 -0.141971
+ 7.11e+10Hz 0.98495 -0.142168
+ 7.12e+10Hz 0.984919 -0.142365
+ 7.13e+10Hz 0.984888 -0.142562
+ 7.14e+10Hz 0.984857 -0.142759
+ 7.15e+10Hz 0.984826 -0.142955
+ 7.16e+10Hz 0.984795 -0.143152
+ 7.17e+10Hz 0.984764 -0.143349
+ 7.18e+10Hz 0.984733 -0.143546
+ 7.19e+10Hz 0.984701 -0.143743
+ 7.2e+10Hz 0.98467 -0.143939
+ 7.21e+10Hz 0.984639 -0.144136
+ 7.22e+10Hz 0.984607 -0.144333
+ 7.23e+10Hz 0.984576 -0.14453
+ 7.24e+10Hz 0.984545 -0.144727
+ 7.25e+10Hz 0.984513 -0.144923
+ 7.26e+10Hz 0.984482 -0.14512
+ 7.27e+10Hz 0.98445 -0.145317
+ 7.28e+10Hz 0.984419 -0.145514
+ 7.29e+10Hz 0.984387 -0.14571
+ 7.3e+10Hz 0.984355 -0.145907
+ 7.31e+10Hz 0.984324 -0.146104
+ 7.32e+10Hz 0.984292 -0.1463
+ 7.33e+10Hz 0.98426 -0.146497
+ 7.34e+10Hz 0.984228 -0.146694
+ 7.35e+10Hz 0.984197 -0.146891
+ 7.36e+10Hz 0.984165 -0.147087
+ 7.37e+10Hz 0.984133 -0.147284
+ 7.38e+10Hz 0.984101 -0.147481
+ 7.39e+10Hz 0.984069 -0.147677
+ 7.4e+10Hz 0.984037 -0.147874
+ 7.41e+10Hz 0.984005 -0.148071
+ 7.42e+10Hz 0.983973 -0.148267
+ 7.43e+10Hz 0.983941 -0.148464
+ 7.44e+10Hz 0.983908 -0.14866
+ 7.45e+10Hz 0.983876 -0.148857
+ 7.46e+10Hz 0.983844 -0.149054
+ 7.47e+10Hz 0.983812 -0.14925
+ 7.48e+10Hz 0.983779 -0.149447
+ 7.49e+10Hz 0.983747 -0.149643
+ 7.5e+10Hz 0.983715 -0.14984
+ 7.51e+10Hz 0.983682 -0.150037
+ 7.52e+10Hz 0.983649 -0.150233
+ 7.53e+10Hz 0.983617 -0.15043
+ 7.54e+10Hz 0.983584 -0.150626
+ 7.55e+10Hz 0.983552 -0.150823
+ 7.56e+10Hz 0.983519 -0.151019
+ 7.57e+10Hz 0.983487 -0.151216
+ 7.58e+10Hz 0.983454 -0.151412
+ 7.59e+10Hz 0.983421 -0.151609
+ 7.6e+10Hz 0.983388 -0.151805
+ 7.61e+10Hz 0.983355 -0.152002
+ 7.62e+10Hz 0.983322 -0.152198
+ 7.63e+10Hz 0.98329 -0.152395
+ 7.64e+10Hz 0.983256 -0.152591
+ 7.65e+10Hz 0.983224 -0.152788
+ 7.66e+10Hz 0.98319 -0.152984
+ 7.67e+10Hz 0.983157 -0.153181
+ 7.68e+10Hz 0.983124 -0.153377
+ 7.69e+10Hz 0.983091 -0.153574
+ 7.7e+10Hz 0.983058 -0.15377
+ 7.71e+10Hz 0.983025 -0.153967
+ 7.72e+10Hz 0.982991 -0.154163
+ 7.73e+10Hz 0.982958 -0.15436
+ 7.74e+10Hz 0.982925 -0.154556
+ 7.75e+10Hz 0.982891 -0.154752
+ 7.76e+10Hz 0.982858 -0.154949
+ 7.77e+10Hz 0.982824 -0.155145
+ 7.78e+10Hz 0.982791 -0.155342
+ 7.79e+10Hz 0.982757 -0.155538
+ 7.8e+10Hz 0.982723 -0.155734
+ 7.81e+10Hz 0.98269 -0.155931
+ 7.82e+10Hz 0.982656 -0.156127
+ 7.83e+10Hz 0.982622 -0.156324
+ 7.84e+10Hz 0.982588 -0.15652
+ 7.85e+10Hz 0.982555 -0.156716
+ 7.86e+10Hz 0.982521 -0.156913
+ 7.87e+10Hz 0.982487 -0.157109
+ 7.88e+10Hz 0.982453 -0.157305
+ 7.89e+10Hz 0.982419 -0.157502
+ 7.9e+10Hz 0.982385 -0.157698
+ 7.91e+10Hz 0.982351 -0.157894
+ 7.92e+10Hz 0.982317 -0.158091
+ 7.93e+10Hz 0.982282 -0.158287
+ 7.94e+10Hz 0.982248 -0.158483
+ 7.95e+10Hz 0.982214 -0.15868
+ 7.96e+10Hz 0.98218 -0.158876
+ 7.97e+10Hz 0.982145 -0.159072
+ 7.98e+10Hz 0.982111 -0.159269
+ 7.99e+10Hz 0.982077 -0.159465
+ 8e+10Hz 0.982042 -0.159661
+ 8.01e+10Hz 0.982008 -0.159857
+ 8.02e+10Hz 0.981973 -0.160054
+ 8.03e+10Hz 0.981939 -0.16025
+ 8.04e+10Hz 0.981904 -0.160446
+ 8.05e+10Hz 0.981869 -0.160642
+ 8.06e+10Hz 0.981835 -0.160839
+ 8.07e+10Hz 0.9818 -0.161035
+ 8.08e+10Hz 0.981765 -0.161231
+ 8.09e+10Hz 0.98173 -0.161427
+ 8.1e+10Hz 0.981695 -0.161624
+ 8.11e+10Hz 0.98166 -0.16182
+ 8.12e+10Hz 0.981625 -0.162016
+ 8.13e+10Hz 0.98159 -0.162212
+ 8.14e+10Hz 0.981555 -0.162408
+ 8.15e+10Hz 0.98152 -0.162605
+ 8.16e+10Hz 0.981485 -0.162801
+ 8.17e+10Hz 0.98145 -0.162997
+ 8.18e+10Hz 0.981414 -0.163193
+ 8.19e+10Hz 0.981379 -0.163389
+ 8.2e+10Hz 0.981344 -0.163585
+ 8.21e+10Hz 0.981308 -0.163781
+ 8.22e+10Hz 0.981273 -0.163978
+ 8.23e+10Hz 0.981237 -0.164174
+ 8.24e+10Hz 0.981202 -0.16437
+ 8.25e+10Hz 0.981167 -0.164566
+ 8.26e+10Hz 0.981131 -0.164762
+ 8.27e+10Hz 0.981095 -0.164958
+ 8.28e+10Hz 0.98106 -0.165154
+ 8.29e+10Hz 0.981024 -0.16535
+ 8.3e+10Hz 0.980988 -0.165546
+ 8.31e+10Hz 0.980952 -0.165742
+ 8.32e+10Hz 0.980916 -0.165939
+ 8.33e+10Hz 0.980881 -0.166135
+ 8.34e+10Hz 0.980845 -0.166331
+ 8.35e+10Hz 0.980808 -0.166527
+ 8.36e+10Hz 0.980773 -0.166723
+ 8.37e+10Hz 0.980736 -0.166919
+ 8.38e+10Hz 0.9807 -0.167115
+ 8.39e+10Hz 0.980664 -0.167311
+ 8.4e+10Hz 0.980628 -0.167507
+ 8.41e+10Hz 0.980592 -0.167703
+ 8.42e+10Hz 0.980555 -0.167899
+ 8.43e+10Hz 0.980519 -0.168095
+ 8.44e+10Hz 0.980483 -0.168291
+ 8.45e+10Hz 0.980446 -0.168487
+ 8.46e+10Hz 0.98041 -0.168683
+ 8.47e+10Hz 0.980373 -0.168879
+ 8.48e+10Hz 0.980336 -0.169075
+ 8.49e+10Hz 0.9803 -0.169271
+ 8.5e+10Hz 0.980263 -0.169466
+ 8.51e+10Hz 0.980226 -0.169662
+ 8.52e+10Hz 0.98019 -0.169858
+ 8.53e+10Hz 0.980153 -0.170054
+ 8.54e+10Hz 0.980116 -0.17025
+ 8.55e+10Hz 0.980079 -0.170446
+ 8.56e+10Hz 0.980042 -0.170642
+ 8.57e+10Hz 0.980005 -0.170838
+ 8.58e+10Hz 0.979968 -0.171034
+ 8.59e+10Hz 0.979931 -0.17123
+ 8.6e+10Hz 0.979894 -0.171425
+ 8.61e+10Hz 0.979857 -0.171621
+ 8.62e+10Hz 0.979819 -0.171817
+ 8.63e+10Hz 0.979782 -0.172013
+ 8.64e+10Hz 0.979745 -0.172209
+ 8.65e+10Hz 0.979708 -0.172404
+ 8.66e+10Hz 0.97967 -0.1726
+ 8.67e+10Hz 0.979633 -0.172796
+ 8.68e+10Hz 0.979595 -0.172992
+ 8.69e+10Hz 0.979558 -0.173187
+ 8.7e+10Hz 0.97952 -0.173383
+ 8.71e+10Hz 0.979483 -0.173579
+ 8.72e+10Hz 0.979445 -0.173775
+ 8.73e+10Hz 0.979407 -0.17397
+ 8.74e+10Hz 0.97937 -0.174166
+ 8.75e+10Hz 0.979332 -0.174362
+ 8.76e+10Hz 0.979294 -0.174558
+ 8.77e+10Hz 0.979256 -0.174753
+ 8.78e+10Hz 0.979218 -0.174949
+ 8.79e+10Hz 0.97918 -0.175145
+ 8.8e+10Hz 0.979142 -0.17534
+ 8.81e+10Hz 0.979104 -0.175536
+ 8.82e+10Hz 0.979066 -0.175731
+ 8.83e+10Hz 0.979028 -0.175927
+ 8.84e+10Hz 0.978989 -0.176123
+ 8.85e+10Hz 0.978951 -0.176318
+ 8.86e+10Hz 0.978913 -0.176514
+ 8.87e+10Hz 0.978875 -0.176709
+ 8.88e+10Hz 0.978836 -0.176905
+ 8.89e+10Hz 0.978798 -0.1771
+ 8.9e+10Hz 0.978759 -0.177296
+ 8.91e+10Hz 0.978721 -0.177491
+ 8.92e+10Hz 0.978682 -0.177687
+ 8.93e+10Hz 0.978644 -0.177882
+ 8.94e+10Hz 0.978605 -0.178078
+ 8.95e+10Hz 0.978566 -0.178274
+ 8.96e+10Hz 0.978528 -0.178469
+ 8.97e+10Hz 0.978489 -0.178664
+ 8.98e+10Hz 0.97845 -0.17886
+ 8.99e+10Hz 0.978411 -0.179055
+ 9e+10Hz 0.978372 -0.179251
+ 9.01e+10Hz 0.978333 -0.179446
+ 9.02e+10Hz 0.978294 -0.179642
+ 9.03e+10Hz 0.978255 -0.179837
+ 9.04e+10Hz 0.978216 -0.180032
+ 9.05e+10Hz 0.978177 -0.180228
+ 9.06e+10Hz 0.978138 -0.180423
+ 9.07e+10Hz 0.978099 -0.180618
+ 9.08e+10Hz 0.978059 -0.180814
+ 9.09e+10Hz 0.97802 -0.181009
+ 9.1e+10Hz 0.977981 -0.181204
+ 9.11e+10Hz 0.977941 -0.181399
+ 9.12e+10Hz 0.977902 -0.181595
+ 9.13e+10Hz 0.977862 -0.18179
+ 9.14e+10Hz 0.977823 -0.181985
+ 9.15e+10Hz 0.977784 -0.18218
+ 9.16e+10Hz 0.977744 -0.182376
+ 9.17e+10Hz 0.977704 -0.182571
+ 9.18e+10Hz 0.977665 -0.182766
+ 9.19e+10Hz 0.977625 -0.182961
+ 9.2e+10Hz 0.977585 -0.183156
+ 9.21e+10Hz 0.977545 -0.183352
+ 9.22e+10Hz 0.977506 -0.183547
+ 9.23e+10Hz 0.977466 -0.183742
+ 9.24e+10Hz 0.977426 -0.183937
+ 9.25e+10Hz 0.977386 -0.184132
+ 9.26e+10Hz 0.977346 -0.184327
+ 9.27e+10Hz 0.977306 -0.184522
+ 9.28e+10Hz 0.977266 -0.184718
+ 9.29e+10Hz 0.977225 -0.184913
+ 9.3e+10Hz 0.977185 -0.185108
+ 9.31e+10Hz 0.977145 -0.185303
+ 9.32e+10Hz 0.977105 -0.185498
+ 9.33e+10Hz 0.977064 -0.185693
+ 9.34e+10Hz 0.977024 -0.185888
+ 9.35e+10Hz 0.976984 -0.186083
+ 9.36e+10Hz 0.976943 -0.186278
+ 9.37e+10Hz 0.976903 -0.186473
+ 9.38e+10Hz 0.976862 -0.186667
+ 9.39e+10Hz 0.976822 -0.186862
+ 9.4e+10Hz 0.976781 -0.187057
+ 9.41e+10Hz 0.976741 -0.187252
+ 9.42e+10Hz 0.9767 -0.187447
+ 9.43e+10Hz 0.976659 -0.187642
+ 9.44e+10Hz 0.976618 -0.187837
+ 9.45e+10Hz 0.976578 -0.188032
+ 9.46e+10Hz 0.976537 -0.188227
+ 9.47e+10Hz 0.976496 -0.188421
+ 9.48e+10Hz 0.976455 -0.188616
+ 9.49e+10Hz 0.976414 -0.188811
+ 9.5e+10Hz 0.976373 -0.189006
+ 9.51e+10Hz 0.976332 -0.189201
+ 9.52e+10Hz 0.976291 -0.189395
+ 9.53e+10Hz 0.97625 -0.18959
+ 9.54e+10Hz 0.976209 -0.189785
+ 9.55e+10Hz 0.976168 -0.18998
+ 9.56e+10Hz 0.976127 -0.190174
+ 9.57e+10Hz 0.976085 -0.190369
+ 9.58e+10Hz 0.976044 -0.190564
+ 9.59e+10Hz 0.976003 -0.190758
+ 9.6e+10Hz 0.975961 -0.190953
+ 9.61e+10Hz 0.97592 -0.191148
+ 9.62e+10Hz 0.975878 -0.191342
+ 9.63e+10Hz 0.975837 -0.191537
+ 9.64e+10Hz 0.975796 -0.191732
+ 9.65e+10Hz 0.975754 -0.191926
+ 9.66e+10Hz 0.975712 -0.192121
+ 9.67e+10Hz 0.975671 -0.192315
+ 9.68e+10Hz 0.975629 -0.19251
+ 9.69e+10Hz 0.975587 -0.192705
+ 9.7e+10Hz 0.975546 -0.192899
+ 9.71e+10Hz 0.975504 -0.193094
+ 9.72e+10Hz 0.975462 -0.193288
+ 9.73e+10Hz 0.97542 -0.193483
+ 9.74e+10Hz 0.975378 -0.193677
+ 9.75e+10Hz 0.975336 -0.193872
+ 9.76e+10Hz 0.975294 -0.194066
+ 9.77e+10Hz 0.975252 -0.194261
+ 9.78e+10Hz 0.97521 -0.194455
+ 9.79e+10Hz 0.975168 -0.19465
+ 9.8e+10Hz 0.975126 -0.194844
+ 9.81e+10Hz 0.975084 -0.195038
+ 9.82e+10Hz 0.975042 -0.195233
+ 9.83e+10Hz 0.975 -0.195427
+ 9.84e+10Hz 0.974957 -0.195622
+ 9.85e+10Hz 0.974915 -0.195816
+ 9.86e+10Hz 0.974873 -0.19601
+ 9.87e+10Hz 0.97483 -0.196205
+ 9.88e+10Hz 0.974788 -0.196399
+ 9.89e+10Hz 0.974745 -0.196593
+ 9.9e+10Hz 0.974703 -0.196788
+ 9.91e+10Hz 0.97466 -0.196982
+ 9.92e+10Hz 0.974618 -0.197176
+ 9.93e+10Hz 0.974575 -0.197371
+ 9.94e+10Hz 0.974533 -0.197565
+ 9.95e+10Hz 0.97449 -0.197759
+ 9.96e+10Hz 0.974447 -0.197954
+ 9.97e+10Hz 0.974405 -0.198148
+ 9.98e+10Hz 0.974362 -0.198342
+ 9.99e+10Hz 0.974319 -0.198536
+ 1e+11Hz 0.974276 -0.198731
+ 1.001e+11Hz 0.974233 -0.198925
+ 1.002e+11Hz 0.97419 -0.199119
+ 1.003e+11Hz 0.974147 -0.199313
+ 1.004e+11Hz 0.974104 -0.199507
+ 1.005e+11Hz 0.974061 -0.199702
+ 1.006e+11Hz 0.974018 -0.199896
+ 1.007e+11Hz 0.973975 -0.20009
+ 1.008e+11Hz 0.973932 -0.200284
+ 1.009e+11Hz 0.973889 -0.200478
+ 1.01e+11Hz 0.973846 -0.200672
+ 1.011e+11Hz 0.973803 -0.200866
+ 1.012e+11Hz 0.973759 -0.201061
+ 1.013e+11Hz 0.973716 -0.201255
+ 1.014e+11Hz 0.973673 -0.201449
+ 1.015e+11Hz 0.973629 -0.201643
+ 1.016e+11Hz 0.973586 -0.201837
+ 1.017e+11Hz 0.973542 -0.202031
+ 1.018e+11Hz 0.973499 -0.202225
+ 1.019e+11Hz 0.973455 -0.202419
+ 1.02e+11Hz 0.973412 -0.202613
+ 1.021e+11Hz 0.973368 -0.202807
+ 1.022e+11Hz 0.973325 -0.203001
+ 1.023e+11Hz 0.973281 -0.203195
+ 1.024e+11Hz 0.973237 -0.203389
+ 1.025e+11Hz 0.973194 -0.203583
+ 1.026e+11Hz 0.97315 -0.203777
+ 1.027e+11Hz 0.973106 -0.203971
+ 1.028e+11Hz 0.973062 -0.204165
+ 1.029e+11Hz 0.973018 -0.204359
+ 1.03e+11Hz 0.972974 -0.204553
+ 1.031e+11Hz 0.97293 -0.204747
+ 1.032e+11Hz 0.972886 -0.204941
+ 1.033e+11Hz 0.972842 -0.205135
+ 1.034e+11Hz 0.972798 -0.205329
+ 1.035e+11Hz 0.972754 -0.205523
+ 1.036e+11Hz 0.97271 -0.205717
+ 1.037e+11Hz 0.972666 -0.205911
+ 1.038e+11Hz 0.972622 -0.206105
+ 1.039e+11Hz 0.972577 -0.206299
+ 1.04e+11Hz 0.972533 -0.206493
+ 1.041e+11Hz 0.972489 -0.206687
+ 1.042e+11Hz 0.972445 -0.20688
+ 1.043e+11Hz 0.9724 -0.207074
+ 1.044e+11Hz 0.972356 -0.207268
+ 1.045e+11Hz 0.972311 -0.207462
+ 1.046e+11Hz 0.972267 -0.207656
+ 1.047e+11Hz 0.972222 -0.20785
+ 1.048e+11Hz 0.972178 -0.208044
+ 1.049e+11Hz 0.972133 -0.208237
+ 1.05e+11Hz 0.972089 -0.208431
+ 1.051e+11Hz 0.972044 -0.208625
+ 1.052e+11Hz 0.971999 -0.208819
+ 1.053e+11Hz 0.971954 -0.209013
+ 1.054e+11Hz 0.97191 -0.209207
+ 1.055e+11Hz 0.971865 -0.2094
+ 1.056e+11Hz 0.97182 -0.209594
+ 1.057e+11Hz 0.971775 -0.209788
+ 1.058e+11Hz 0.97173 -0.209982
+ 1.059e+11Hz 0.971685 -0.210176
+ 1.06e+11Hz 0.97164 -0.210369
+ 1.061e+11Hz 0.971595 -0.210563
+ 1.062e+11Hz 0.97155 -0.210757
+ 1.063e+11Hz 0.971505 -0.210951
+ 1.064e+11Hz 0.97146 -0.211145
+ 1.065e+11Hz 0.971414 -0.211338
+ 1.066e+11Hz 0.971369 -0.211532
+ 1.067e+11Hz 0.971324 -0.211726
+ 1.068e+11Hz 0.971279 -0.21192
+ 1.069e+11Hz 0.971233 -0.212113
+ 1.07e+11Hz 0.971188 -0.212307
+ 1.071e+11Hz 0.971143 -0.212501
+ 1.072e+11Hz 0.971097 -0.212695
+ 1.073e+11Hz 0.971051 -0.212888
+ 1.074e+11Hz 0.971006 -0.213082
+ 1.075e+11Hz 0.97096 -0.213276
+ 1.076e+11Hz 0.970915 -0.213469
+ 1.077e+11Hz 0.970869 -0.213663
+ 1.078e+11Hz 0.970823 -0.213857
+ 1.079e+11Hz 0.970778 -0.21405
+ 1.08e+11Hz 0.970732 -0.214244
+ 1.081e+11Hz 0.970686 -0.214438
+ 1.082e+11Hz 0.97064 -0.214631
+ 1.083e+11Hz 0.970594 -0.214825
+ 1.084e+11Hz 0.970548 -0.215019
+ 1.085e+11Hz 0.970502 -0.215212
+ 1.086e+11Hz 0.970456 -0.215406
+ 1.087e+11Hz 0.97041 -0.2156
+ 1.088e+11Hz 0.970364 -0.215793
+ 1.089e+11Hz 0.970318 -0.215987
+ 1.09e+11Hz 0.970272 -0.21618
+ 1.091e+11Hz 0.970226 -0.216374
+ 1.092e+11Hz 0.970179 -0.216568
+ 1.093e+11Hz 0.970133 -0.216761
+ 1.094e+11Hz 0.970087 -0.216955
+ 1.095e+11Hz 0.97004 -0.217148
+ 1.096e+11Hz 0.969994 -0.217342
+ 1.097e+11Hz 0.969948 -0.217536
+ 1.098e+11Hz 0.969901 -0.217729
+ 1.099e+11Hz 0.969854 -0.217923
+ 1.1e+11Hz 0.969808 -0.218116
+ 1.101e+11Hz 0.969761 -0.21831
+ 1.102e+11Hz 0.969715 -0.218503
+ 1.103e+11Hz 0.969668 -0.218697
+ 1.104e+11Hz 0.969621 -0.21889
+ 1.105e+11Hz 0.969574 -0.219084
+ 1.106e+11Hz 0.969528 -0.219277
+ 1.107e+11Hz 0.969481 -0.219471
+ 1.108e+11Hz 0.969434 -0.219664
+ 1.109e+11Hz 0.969387 -0.219858
+ 1.11e+11Hz 0.96934 -0.220051
+ 1.111e+11Hz 0.969293 -0.220245
+ 1.112e+11Hz 0.969246 -0.220438
+ 1.113e+11Hz 0.969199 -0.220632
+ 1.114e+11Hz 0.969151 -0.220825
+ 1.115e+11Hz 0.969104 -0.221019
+ 1.116e+11Hz 0.969057 -0.221212
+ 1.117e+11Hz 0.96901 -0.221406
+ 1.118e+11Hz 0.968962 -0.221599
+ 1.119e+11Hz 0.968915 -0.221792
+ 1.12e+11Hz 0.968867 -0.221986
+ 1.121e+11Hz 0.96882 -0.222179
+ 1.122e+11Hz 0.968773 -0.222373
+ 1.123e+11Hz 0.968725 -0.222566
+ 1.124e+11Hz 0.968677 -0.222759
+ 1.125e+11Hz 0.96863 -0.222953
+ 1.126e+11Hz 0.968582 -0.223146
+ 1.127e+11Hz 0.968534 -0.223339
+ 1.128e+11Hz 0.968487 -0.223533
+ 1.129e+11Hz 0.968439 -0.223726
+ 1.13e+11Hz 0.968391 -0.223919
+ 1.131e+11Hz 0.968343 -0.224112
+ 1.132e+11Hz 0.968295 -0.224306
+ 1.133e+11Hz 0.968247 -0.224499
+ 1.134e+11Hz 0.968199 -0.224692
+ 1.135e+11Hz 0.968151 -0.224886
+ 1.136e+11Hz 0.968103 -0.225079
+ 1.137e+11Hz 0.968055 -0.225272
+ 1.138e+11Hz 0.968007 -0.225465
+ 1.139e+11Hz 0.967958 -0.225659
+ 1.14e+11Hz 0.96791 -0.225852
+ 1.141e+11Hz 0.967862 -0.226045
+ 1.142e+11Hz 0.967813 -0.226238
+ 1.143e+11Hz 0.967765 -0.226431
+ 1.144e+11Hz 0.967716 -0.226624
+ 1.145e+11Hz 0.967668 -0.226818
+ 1.146e+11Hz 0.967619 -0.227011
+ 1.147e+11Hz 0.967571 -0.227204
+ 1.148e+11Hz 0.967522 -0.227397
+ 1.149e+11Hz 0.967473 -0.22759
+ 1.15e+11Hz 0.967425 -0.227783
+ 1.151e+11Hz 0.967376 -0.227976
+ 1.152e+11Hz 0.967327 -0.228169
+ 1.153e+11Hz 0.967278 -0.228362
+ 1.154e+11Hz 0.967229 -0.228555
+ 1.155e+11Hz 0.96718 -0.228748
+ 1.156e+11Hz 0.967132 -0.228941
+ 1.157e+11Hz 0.967082 -0.229134
+ 1.158e+11Hz 0.967033 -0.229327
+ 1.159e+11Hz 0.966984 -0.22952
+ 1.16e+11Hz 0.966935 -0.229713
+ 1.161e+11Hz 0.966886 -0.229906
+ 1.162e+11Hz 0.966837 -0.230099
+ 1.163e+11Hz 0.966787 -0.230292
+ 1.164e+11Hz 0.966738 -0.230485
+ 1.165e+11Hz 0.966689 -0.230677
+ 1.166e+11Hz 0.966639 -0.23087
+ 1.167e+11Hz 0.96659 -0.231063
+ 1.168e+11Hz 0.96654 -0.231256
+ 1.169e+11Hz 0.966491 -0.231449
+ 1.17e+11Hz 0.966441 -0.231642
+ 1.171e+11Hz 0.966391 -0.231834
+ 1.172e+11Hz 0.966342 -0.232027
+ 1.173e+11Hz 0.966292 -0.23222
+ 1.174e+11Hz 0.966242 -0.232412
+ 1.175e+11Hz 0.966192 -0.232605
+ 1.176e+11Hz 0.966143 -0.232798
+ 1.177e+11Hz 0.966093 -0.23299
+ 1.178e+11Hz 0.966043 -0.233183
+ 1.179e+11Hz 0.965993 -0.233376
+ 1.18e+11Hz 0.965943 -0.233568
+ 1.181e+11Hz 0.965893 -0.233761
+ 1.182e+11Hz 0.965843 -0.233954
+ 1.183e+11Hz 0.965792 -0.234146
+ 1.184e+11Hz 0.965742 -0.234339
+ 1.185e+11Hz 0.965692 -0.234531
+ 1.186e+11Hz 0.965642 -0.234724
+ 1.187e+11Hz 0.965591 -0.234916
+ 1.188e+11Hz 0.965541 -0.235108
+ 1.189e+11Hz 0.965491 -0.235301
+ 1.19e+11Hz 0.96544 -0.235493
+ 1.191e+11Hz 0.96539 -0.235686
+ 1.192e+11Hz 0.965339 -0.235878
+ 1.193e+11Hz 0.965289 -0.23607
+ 1.194e+11Hz 0.965238 -0.236263
+ 1.195e+11Hz 0.965187 -0.236455
+ 1.196e+11Hz 0.965137 -0.236648
+ 1.197e+11Hz 0.965086 -0.23684
+ 1.198e+11Hz 0.965035 -0.237032
+ 1.199e+11Hz 0.964984 -0.237224
+ 1.2e+11Hz 0.964933 -0.237416
+ 1.201e+11Hz 0.964883 -0.237609
+ 1.202e+11Hz 0.964832 -0.237801
+ 1.203e+11Hz 0.964781 -0.237993
+ 1.204e+11Hz 0.96473 -0.238185
+ 1.205e+11Hz 0.964679 -0.238377
+ 1.206e+11Hz 0.964627 -0.238569
+ 1.207e+11Hz 0.964576 -0.238761
+ 1.208e+11Hz 0.964525 -0.238953
+ 1.209e+11Hz 0.964474 -0.239145
+ 1.21e+11Hz 0.964423 -0.239337
+ 1.211e+11Hz 0.964372 -0.239529
+ 1.212e+11Hz 0.96432 -0.239721
+ 1.213e+11Hz 0.964269 -0.239913
+ 1.214e+11Hz 0.964217 -0.240105
+ 1.215e+11Hz 0.964166 -0.240297
+ 1.216e+11Hz 0.964114 -0.240489
+ 1.217e+11Hz 0.964063 -0.240681
+ 1.218e+11Hz 0.964011 -0.240873
+ 1.219e+11Hz 0.96396 -0.241064
+ 1.22e+11Hz 0.963908 -0.241256
+ 1.221e+11Hz 0.963857 -0.241448
+ 1.222e+11Hz 0.963805 -0.24164
+ 1.223e+11Hz 0.963753 -0.241831
+ 1.224e+11Hz 0.963701 -0.242023
+ 1.225e+11Hz 0.96365 -0.242215
+ 1.226e+11Hz 0.963598 -0.242406
+ 1.227e+11Hz 0.963546 -0.242598
+ 1.228e+11Hz 0.963494 -0.24279
+ 1.229e+11Hz 0.963442 -0.242981
+ 1.23e+11Hz 0.96339 -0.243173
+ 1.231e+11Hz 0.963338 -0.243364
+ 1.232e+11Hz 0.963286 -0.243556
+ 1.233e+11Hz 0.963234 -0.243747
+ 1.234e+11Hz 0.963182 -0.243939
+ 1.235e+11Hz 0.963129 -0.24413
+ 1.236e+11Hz 0.963077 -0.244322
+ 1.237e+11Hz 0.963025 -0.244513
+ 1.238e+11Hz 0.962973 -0.244704
+ 1.239e+11Hz 0.96292 -0.244896
+ 1.24e+11Hz 0.962868 -0.245087
+ 1.241e+11Hz 0.962816 -0.245278
+ 1.242e+11Hz 0.962763 -0.24547
+ 1.243e+11Hz 0.962711 -0.245661
+ 1.244e+11Hz 0.962658 -0.245852
+ 1.245e+11Hz 0.962606 -0.246043
+ 1.246e+11Hz 0.962553 -0.246234
+ 1.247e+11Hz 0.962501 -0.246426
+ 1.248e+11Hz 0.962448 -0.246617
+ 1.249e+11Hz 0.962395 -0.246808
+ 1.25e+11Hz 0.962343 -0.246999
+ 1.251e+11Hz 0.96229 -0.24719
+ 1.252e+11Hz 0.962237 -0.247381
+ 1.253e+11Hz 0.962185 -0.247572
+ 1.254e+11Hz 0.962132 -0.247763
+ 1.255e+11Hz 0.962079 -0.247954
+ 1.256e+11Hz 0.962026 -0.248145
+ 1.257e+11Hz 0.961973 -0.248336
+ 1.258e+11Hz 0.96192 -0.248527
+ 1.259e+11Hz 0.961867 -0.248718
+ 1.26e+11Hz 0.961814 -0.248909
+ 1.261e+11Hz 0.961761 -0.2491
+ 1.262e+11Hz 0.961708 -0.24929
+ 1.263e+11Hz 0.961655 -0.249481
+ 1.264e+11Hz 0.961602 -0.249672
+ 1.265e+11Hz 0.961549 -0.249863
+ 1.266e+11Hz 0.961496 -0.250054
+ 1.267e+11Hz 0.961442 -0.250244
+ 1.268e+11Hz 0.961389 -0.250435
+ 1.269e+11Hz 0.961336 -0.250626
+ 1.27e+11Hz 0.961283 -0.250816
+ 1.271e+11Hz 0.961229 -0.251007
+ 1.272e+11Hz 0.961176 -0.251198
+ 1.273e+11Hz 0.961123 -0.251388
+ 1.274e+11Hz 0.961069 -0.251579
+ 1.275e+11Hz 0.961016 -0.251769
+ 1.276e+11Hz 0.960962 -0.25196
+ 1.277e+11Hz 0.960909 -0.252151
+ 1.278e+11Hz 0.960855 -0.252341
+ 1.279e+11Hz 0.960802 -0.252532
+ 1.28e+11Hz 0.960748 -0.252722
+ 1.281e+11Hz 0.960694 -0.252912
+ 1.282e+11Hz 0.960641 -0.253103
+ 1.283e+11Hz 0.960587 -0.253293
+ 1.284e+11Hz 0.960533 -0.253484
+ 1.285e+11Hz 0.96048 -0.253674
+ 1.286e+11Hz 0.960426 -0.253865
+ 1.287e+11Hz 0.960372 -0.254055
+ 1.288e+11Hz 0.960318 -0.254245
+ 1.289e+11Hz 0.960264 -0.254436
+ 1.29e+11Hz 0.96021 -0.254626
+ 1.291e+11Hz 0.960157 -0.254816
+ 1.292e+11Hz 0.960103 -0.255006
+ 1.293e+11Hz 0.960049 -0.255197
+ 1.294e+11Hz 0.959995 -0.255387
+ 1.295e+11Hz 0.959941 -0.255577
+ 1.296e+11Hz 0.959887 -0.255767
+ 1.297e+11Hz 0.959832 -0.255958
+ 1.298e+11Hz 0.959778 -0.256148
+ 1.299e+11Hz 0.959724 -0.256338
+ 1.3e+11Hz 0.95967 -0.256528
+ 1.301e+11Hz 0.959616 -0.256718
+ 1.302e+11Hz 0.959562 -0.256908
+ 1.303e+11Hz 0.959507 -0.257098
+ 1.304e+11Hz 0.959453 -0.257288
+ 1.305e+11Hz 0.959399 -0.257479
+ 1.306e+11Hz 0.959344 -0.257669
+ 1.307e+11Hz 0.95929 -0.257859
+ 1.308e+11Hz 0.959236 -0.258049
+ 1.309e+11Hz 0.959181 -0.258239
+ 1.31e+11Hz 0.959127 -0.258429
+ 1.311e+11Hz 0.959072 -0.258619
+ 1.312e+11Hz 0.959018 -0.258809
+ 1.313e+11Hz 0.958963 -0.258999
+ 1.314e+11Hz 0.958909 -0.259189
+ 1.315e+11Hz 0.958854 -0.259379
+ 1.316e+11Hz 0.958799 -0.259569
+ 1.317e+11Hz 0.958744 -0.259759
+ 1.318e+11Hz 0.95869 -0.259949
+ 1.319e+11Hz 0.958635 -0.260138
+ 1.32e+11Hz 0.95858 -0.260328
+ 1.321e+11Hz 0.958525 -0.260518
+ 1.322e+11Hz 0.958471 -0.260708
+ 1.323e+11Hz 0.958416 -0.260898
+ 1.324e+11Hz 0.958361 -0.261088
+ 1.325e+11Hz 0.958306 -0.261278
+ 1.326e+11Hz 0.958251 -0.261468
+ 1.327e+11Hz 0.958196 -0.261657
+ 1.328e+11Hz 0.958141 -0.261847
+ 1.329e+11Hz 0.958086 -0.262037
+ 1.33e+11Hz 0.958031 -0.262227
+ 1.331e+11Hz 0.957975 -0.262417
+ 1.332e+11Hz 0.95792 -0.262607
+ 1.333e+11Hz 0.957865 -0.262796
+ 1.334e+11Hz 0.95781 -0.262986
+ 1.335e+11Hz 0.957755 -0.263176
+ 1.336e+11Hz 0.957699 -0.263366
+ 1.337e+11Hz 0.957644 -0.263555
+ 1.338e+11Hz 0.957589 -0.263745
+ 1.339e+11Hz 0.957533 -0.263935
+ 1.34e+11Hz 0.957478 -0.264125
+ 1.341e+11Hz 0.957422 -0.264314
+ 1.342e+11Hz 0.957367 -0.264504
+ 1.343e+11Hz 0.957311 -0.264694
+ 1.344e+11Hz 0.957256 -0.264884
+ 1.345e+11Hz 0.9572 -0.265073
+ 1.346e+11Hz 0.957144 -0.265263
+ 1.347e+11Hz 0.957089 -0.265453
+ 1.348e+11Hz 0.957033 -0.265643
+ 1.349e+11Hz 0.956977 -0.265832
+ 1.35e+11Hz 0.956921 -0.266022
+ 1.351e+11Hz 0.956865 -0.266212
+ 1.352e+11Hz 0.956809 -0.266401
+ 1.353e+11Hz 0.956753 -0.266591
+ 1.354e+11Hz 0.956697 -0.266781
+ 1.355e+11Hz 0.956641 -0.26697
+ 1.356e+11Hz 0.956585 -0.26716
+ 1.357e+11Hz 0.956529 -0.26735
+ 1.358e+11Hz 0.956473 -0.267539
+ 1.359e+11Hz 0.956417 -0.267729
+ 1.36e+11Hz 0.956361 -0.267919
+ 1.361e+11Hz 0.956304 -0.268108
+ 1.362e+11Hz 0.956248 -0.268298
+ 1.363e+11Hz 0.956192 -0.268488
+ 1.364e+11Hz 0.956135 -0.268677
+ 1.365e+11Hz 0.956079 -0.268867
+ 1.366e+11Hz 0.956022 -0.269057
+ 1.367e+11Hz 0.955966 -0.269246
+ 1.368e+11Hz 0.955909 -0.269436
+ 1.369e+11Hz 0.955852 -0.269626
+ 1.37e+11Hz 0.955796 -0.269815
+ 1.371e+11Hz 0.955739 -0.270005
+ 1.372e+11Hz 0.955682 -0.270195
+ 1.373e+11Hz 0.955626 -0.270384
+ 1.374e+11Hz 0.955569 -0.270574
+ 1.375e+11Hz 0.955512 -0.270763
+ 1.376e+11Hz 0.955455 -0.270953
+ 1.377e+11Hz 0.955398 -0.271143
+ 1.378e+11Hz 0.955341 -0.271332
+ 1.379e+11Hz 0.955283 -0.271522
+ 1.38e+11Hz 0.955226 -0.271712
+ 1.381e+11Hz 0.955169 -0.271901
+ 1.382e+11Hz 0.955112 -0.272091
+ 1.383e+11Hz 0.955055 -0.27228
+ 1.384e+11Hz 0.954997 -0.27247
+ 1.385e+11Hz 0.95494 -0.27266
+ 1.386e+11Hz 0.954882 -0.272849
+ 1.387e+11Hz 0.954825 -0.273039
+ 1.388e+11Hz 0.954767 -0.273228
+ 1.389e+11Hz 0.954709 -0.273418
+ 1.39e+11Hz 0.954652 -0.273608
+ 1.391e+11Hz 0.954594 -0.273797
+ 1.392e+11Hz 0.954536 -0.273987
+ 1.393e+11Hz 0.954478 -0.274176
+ 1.394e+11Hz 0.95442 -0.274366
+ 1.395e+11Hz 0.954363 -0.274556
+ 1.396e+11Hz 0.954304 -0.274745
+ 1.397e+11Hz 0.954246 -0.274935
+ 1.398e+11Hz 0.954188 -0.275124
+ 1.399e+11Hz 0.95413 -0.275314
+ 1.4e+11Hz 0.954072 -0.275503
+ 1.401e+11Hz 0.954013 -0.275693
+ 1.402e+11Hz 0.953955 -0.275882
+ 1.403e+11Hz 0.953897 -0.276072
+ 1.404e+11Hz 0.953838 -0.276261
+ 1.405e+11Hz 0.95378 -0.276451
+ 1.406e+11Hz 0.953721 -0.27664
+ 1.407e+11Hz 0.953662 -0.27683
+ 1.408e+11Hz 0.953604 -0.277019
+ 1.409e+11Hz 0.953545 -0.277209
+ 1.41e+11Hz 0.953486 -0.277398
+ 1.411e+11Hz 0.953427 -0.277588
+ 1.412e+11Hz 0.953368 -0.277777
+ 1.413e+11Hz 0.953309 -0.277967
+ 1.414e+11Hz 0.95325 -0.278156
+ 1.415e+11Hz 0.953191 -0.278346
+ 1.416e+11Hz 0.953131 -0.278535
+ 1.417e+11Hz 0.953072 -0.278725
+ 1.418e+11Hz 0.953013 -0.278914
+ 1.419e+11Hz 0.952953 -0.279103
+ 1.42e+11Hz 0.952894 -0.279293
+ 1.421e+11Hz 0.952834 -0.279482
+ 1.422e+11Hz 0.952774 -0.279672
+ 1.423e+11Hz 0.952715 -0.279861
+ 1.424e+11Hz 0.952655 -0.28005
+ 1.425e+11Hz 0.952595 -0.28024
+ 1.426e+11Hz 0.952535 -0.280429
+ 1.427e+11Hz 0.952475 -0.280618
+ 1.428e+11Hz 0.952415 -0.280808
+ 1.429e+11Hz 0.952355 -0.280997
+ 1.43e+11Hz 0.952295 -0.281186
+ 1.431e+11Hz 0.952235 -0.281375
+ 1.432e+11Hz 0.952175 -0.281565
+ 1.433e+11Hz 0.952114 -0.281754
+ 1.434e+11Hz 0.952054 -0.281943
+ 1.435e+11Hz 0.951993 -0.282132
+ 1.436e+11Hz 0.951933 -0.282322
+ 1.437e+11Hz 0.951872 -0.282511
+ 1.438e+11Hz 0.951811 -0.2827
+ 1.439e+11Hz 0.95175 -0.282889
+ 1.44e+11Hz 0.95169 -0.283078
+ 1.441e+11Hz 0.951629 -0.283267
+ 1.442e+11Hz 0.951568 -0.283456
+ 1.443e+11Hz 0.951507 -0.283645
+ 1.444e+11Hz 0.951446 -0.283834
+ 1.445e+11Hz 0.951384 -0.284023
+ 1.446e+11Hz 0.951323 -0.284212
+ 1.447e+11Hz 0.951262 -0.284401
+ 1.448e+11Hz 0.9512 -0.28459
+ 1.449e+11Hz 0.951139 -0.284779
+ 1.45e+11Hz 0.951077 -0.284968
+ 1.451e+11Hz 0.951016 -0.285157
+ 1.452e+11Hz 0.950954 -0.285346
+ 1.453e+11Hz 0.950892 -0.285535
+ 1.454e+11Hz 0.950831 -0.285724
+ 1.455e+11Hz 0.950769 -0.285912
+ 1.456e+11Hz 0.950707 -0.286101
+ 1.457e+11Hz 0.950645 -0.28629
+ 1.458e+11Hz 0.950582 -0.286479
+ 1.459e+11Hz 0.95052 -0.286667
+ 1.46e+11Hz 0.950458 -0.286856
+ 1.461e+11Hz 0.950396 -0.287045
+ 1.462e+11Hz 0.950334 -0.287233
+ 1.463e+11Hz 0.950271 -0.287422
+ 1.464e+11Hz 0.950209 -0.28761
+ 1.465e+11Hz 0.950146 -0.287799
+ 1.466e+11Hz 0.950083 -0.287988
+ 1.467e+11Hz 0.950021 -0.288176
+ 1.468e+11Hz 0.949958 -0.288364
+ 1.469e+11Hz 0.949895 -0.288553
+ 1.47e+11Hz 0.949832 -0.288741
+ 1.471e+11Hz 0.949769 -0.28893
+ 1.472e+11Hz 0.949706 -0.289118
+ 1.473e+11Hz 0.949643 -0.289306
+ 1.474e+11Hz 0.94958 -0.289494
+ 1.475e+11Hz 0.949517 -0.289683
+ 1.476e+11Hz 0.949453 -0.289871
+ 1.477e+11Hz 0.94939 -0.290059
+ 1.478e+11Hz 0.949327 -0.290247
+ 1.479e+11Hz 0.949263 -0.290435
+ 1.48e+11Hz 0.9492 -0.290623
+ 1.481e+11Hz 0.949136 -0.290811
+ 1.482e+11Hz 0.949072 -0.290999
+ 1.483e+11Hz 0.949009 -0.291187
+ 1.484e+11Hz 0.948945 -0.291375
+ 1.485e+11Hz 0.948881 -0.291563
+ 1.486e+11Hz 0.948817 -0.291751
+ 1.487e+11Hz 0.948753 -0.291939
+ 1.488e+11Hz 0.948689 -0.292126
+ 1.489e+11Hz 0.948625 -0.292314
+ 1.49e+11Hz 0.948561 -0.292502
+ 1.491e+11Hz 0.948497 -0.292689
+ 1.492e+11Hz 0.948433 -0.292877
+ 1.493e+11Hz 0.948368 -0.293065
+ 1.494e+11Hz 0.948304 -0.293252
+ 1.495e+11Hz 0.94824 -0.29344
+ 1.496e+11Hz 0.948175 -0.293627
+ 1.497e+11Hz 0.948111 -0.293815
+ 1.498e+11Hz 0.948046 -0.294002
+ 1.499e+11Hz 0.947982 -0.294189
+ 1.5e+11Hz 0.947917 -0.294377
+ ]

A22 %vd(20 3) %vd(22, 3) xfer4
.model xfer4 xfer R_I=true table=[
+ 0Hz 0.00293424 0
+ 1e+08Hz 0.00293429 5.75275e-05
+ 2e+08Hz 0.00293444 0.000115054
+ 3e+08Hz 0.00293469 0.000172577
+ 4e+08Hz 0.00293504 0.000230096
+ 5e+08Hz 0.00293549 0.00028761
+ 6e+08Hz 0.00293604 0.000345117
+ 7e+08Hz 0.00293669 0.000402615
+ 8e+08Hz 0.00293744 0.000460104
+ 9e+08Hz 0.00293828 0.000517582
+ 1e+09Hz 0.00293923 0.000575048
+ 1.1e+09Hz 0.00294027 0.0006325
+ 1.2e+09Hz 0.00294142 0.000689936
+ 1.3e+09Hz 0.00294266 0.000747357
+ 1.4e+09Hz 0.002944 0.00080476
+ 1.5e+09Hz 0.00294543 0.000862143
+ 1.6e+09Hz 0.00294697 0.000919506
+ 1.7e+09Hz 0.0029486 0.000976848
+ 1.8e+09Hz 0.00295032 0.00103417
+ 1.9e+09Hz 0.00295214 0.00109146
+ 2e+09Hz 0.00295406 0.00114873
+ 2.1e+09Hz 0.00295607 0.00120597
+ 2.2e+09Hz 0.00295817 0.00126319
+ 2.3e+09Hz 0.00296037 0.00132037
+ 2.4e+09Hz 0.00296267 0.00137753
+ 2.5e+09Hz 0.00296505 0.00143465
+ 2.6e+09Hz 0.00296752 0.00149174
+ 2.7e+09Hz 0.00297009 0.00154879
+ 2.8e+09Hz 0.00297275 0.00160581
+ 2.9e+09Hz 0.00297549 0.0016628
+ 3e+09Hz 0.00297833 0.00171975
+ 3.1e+09Hz 0.00298125 0.00177665
+ 3.2e+09Hz 0.00298427 0.00183352
+ 3.3e+09Hz 0.00298737 0.00189035
+ 3.4e+09Hz 0.00299055 0.00194714
+ 3.5e+09Hz 0.00299382 0.00200388
+ 3.6e+09Hz 0.00299717 0.00206058
+ 3.7e+09Hz 0.00300061 0.00211723
+ 3.8e+09Hz 0.00300413 0.00217384
+ 3.9e+09Hz 0.00300773 0.0022304
+ 4e+09Hz 0.00301141 0.00228692
+ 4.1e+09Hz 0.00301517 0.00234338
+ 4.2e+09Hz 0.00301901 0.0023998
+ 4.3e+09Hz 0.00302293 0.00245616
+ 4.4e+09Hz 0.00302693 0.00251248
+ 4.5e+09Hz 0.003031 0.00256874
+ 4.6e+09Hz 0.00303514 0.00262495
+ 4.7e+09Hz 0.00303937 0.00268111
+ 4.8e+09Hz 0.00304366 0.00273721
+ 4.9e+09Hz 0.00304803 0.00279325
+ 5e+09Hz 0.00305246 0.00284924
+ 5.1e+09Hz 0.00305697 0.00290517
+ 5.2e+09Hz 0.00306154 0.00296105
+ 5.3e+09Hz 0.00306619 0.00301687
+ 5.4e+09Hz 0.0030709 0.00307263
+ 5.5e+09Hz 0.00307567 0.00312833
+ 5.6e+09Hz 0.00308051 0.00318397
+ 5.7e+09Hz 0.00308542 0.00323955
+ 5.8e+09Hz 0.00309038 0.00329507
+ 5.9e+09Hz 0.00309541 0.00335053
+ 6e+09Hz 0.0031005 0.00340593
+ 6.1e+09Hz 0.00310564 0.00346126
+ 6.2e+09Hz 0.00311085 0.00351653
+ 6.3e+09Hz 0.00311611 0.00357174
+ 6.4e+09Hz 0.00312143 0.00362689
+ 6.5e+09Hz 0.0031268 0.00368197
+ 6.6e+09Hz 0.00313222 0.00373699
+ 6.7e+09Hz 0.0031377 0.00379194
+ 6.8e+09Hz 0.00314323 0.00384683
+ 6.9e+09Hz 0.00314881 0.00390166
+ 7e+09Hz 0.00315444 0.00395641
+ 7.1e+09Hz 0.00316011 0.00401111
+ 7.2e+09Hz 0.00316583 0.00406574
+ 7.3e+09Hz 0.0031716 0.0041203
+ 7.4e+09Hz 0.00317741 0.0041748
+ 7.5e+09Hz 0.00318327 0.00422923
+ 7.6e+09Hz 0.00318916 0.00428359
+ 7.7e+09Hz 0.0031951 0.00433789
+ 7.8e+09Hz 0.00320108 0.00439212
+ 7.9e+09Hz 0.0032071 0.00444629
+ 8e+09Hz 0.00321315 0.00450039
+ 8.1e+09Hz 0.00321924 0.00455442
+ 8.2e+09Hz 0.00322537 0.00460839
+ 8.3e+09Hz 0.00323153 0.00466229
+ 8.4e+09Hz 0.00323772 0.00471613
+ 8.5e+09Hz 0.00324395 0.0047699
+ 8.6e+09Hz 0.00325021 0.0048236
+ 8.7e+09Hz 0.0032565 0.00487724
+ 8.8e+09Hz 0.00326282 0.00493081
+ 8.9e+09Hz 0.00326916 0.00498432
+ 9e+09Hz 0.00327553 0.00503776
+ 9.1e+09Hz 0.00328193 0.00509114
+ 9.2e+09Hz 0.00328836 0.00514445
+ 9.3e+09Hz 0.0032948 0.0051977
+ 9.4e+09Hz 0.00330128 0.00525089
+ 9.5e+09Hz 0.00330777 0.00530401
+ 9.6e+09Hz 0.00331428 0.00535707
+ 9.7e+09Hz 0.00332082 0.00541006
+ 9.8e+09Hz 0.00332737 0.00546299
+ 9.9e+09Hz 0.00333394 0.00551586
+ 1e+10Hz 0.00334053 0.00556867
+ 1.01e+10Hz 0.00334714 0.00562141
+ 1.02e+10Hz 0.00335376 0.0056741
+ 1.03e+10Hz 0.0033604 0.00572672
+ 1.04e+10Hz 0.00336705 0.00577929
+ 1.05e+10Hz 0.00337371 0.00583179
+ 1.06e+10Hz 0.00338039 0.00588423
+ 1.07e+10Hz 0.00338707 0.00593662
+ 1.08e+10Hz 0.00339377 0.00598894
+ 1.09e+10Hz 0.00340048 0.00604121
+ 1.1e+10Hz 0.0034072 0.00609342
+ 1.11e+10Hz 0.00341392 0.00614558
+ 1.12e+10Hz 0.00342065 0.00619768
+ 1.13e+10Hz 0.00342739 0.00624972
+ 1.14e+10Hz 0.00343414 0.00630171
+ 1.15e+10Hz 0.00344089 0.00635364
+ 1.16e+10Hz 0.00344765 0.00640552
+ 1.17e+10Hz 0.0034544 0.00645734
+ 1.18e+10Hz 0.00346117 0.00650911
+ 1.19e+10Hz 0.00346793 0.00656083
+ 1.2e+10Hz 0.0034747 0.0066125
+ 1.21e+10Hz 0.00348147 0.00666412
+ 1.22e+10Hz 0.00348824 0.00671568
+ 1.23e+10Hz 0.00349501 0.0067672
+ 1.24e+10Hz 0.00350178 0.00681867
+ 1.25e+10Hz 0.00350855 0.00687008
+ 1.26e+10Hz 0.00351532 0.00692146
+ 1.27e+10Hz 0.00352209 0.00697278
+ 1.28e+10Hz 0.00352885 0.00702406
+ 1.29e+10Hz 0.00353562 0.00707529
+ 1.3e+10Hz 0.00354237 0.00712648
+ 1.31e+10Hz 0.00354913 0.00717762
+ 1.32e+10Hz 0.00355588 0.00722872
+ 1.33e+10Hz 0.00356263 0.00727977
+ 1.34e+10Hz 0.00356937 0.00733078
+ 1.35e+10Hz 0.0035761 0.00738175
+ 1.36e+10Hz 0.00358283 0.00743268
+ 1.37e+10Hz 0.00358956 0.00748357
+ 1.38e+10Hz 0.00359628 0.00753442
+ 1.39e+10Hz 0.00360299 0.00758523
+ 1.4e+10Hz 0.00360969 0.00763601
+ 1.41e+10Hz 0.00361639 0.00768674
+ 1.42e+10Hz 0.00362308 0.00773744
+ 1.43e+10Hz 0.00362976 0.0077881
+ 1.44e+10Hz 0.00363644 0.00783873
+ 1.45e+10Hz 0.0036431 0.00788932
+ 1.46e+10Hz 0.00364976 0.00793988
+ 1.47e+10Hz 0.00365641 0.0079904
+ 1.48e+10Hz 0.00366305 0.00804089
+ 1.49e+10Hz 0.00366968 0.00809135
+ 1.5e+10Hz 0.0036763 0.00814178
+ 1.51e+10Hz 0.00368291 0.00819218
+ 1.52e+10Hz 0.00368951 0.00824255
+ 1.53e+10Hz 0.0036961 0.00829289
+ 1.54e+10Hz 0.00370269 0.0083432
+ 1.55e+10Hz 0.00370926 0.00839348
+ 1.56e+10Hz 0.00371582 0.00844374
+ 1.57e+10Hz 0.00372237 0.00849397
+ 1.58e+10Hz 0.00372892 0.00854417
+ 1.59e+10Hz 0.00373545 0.00859435
+ 1.6e+10Hz 0.00374197 0.0086445
+ 1.61e+10Hz 0.00374849 0.00869463
+ 1.62e+10Hz 0.00375499 0.00874474
+ 1.63e+10Hz 0.00376148 0.00879482
+ 1.64e+10Hz 0.00376796 0.00884489
+ 1.65e+10Hz 0.00377443 0.00889493
+ 1.66e+10Hz 0.00378089 0.00894495
+ 1.67e+10Hz 0.00378735 0.00899495
+ 1.68e+10Hz 0.00379379 0.00904493
+ 1.69e+10Hz 0.00380022 0.00909489
+ 1.7e+10Hz 0.00380664 0.00914483
+ 1.71e+10Hz 0.00381305 0.00919476
+ 1.72e+10Hz 0.00381945 0.00924467
+ 1.73e+10Hz 0.00382585 0.00929456
+ 1.74e+10Hz 0.00383223 0.00934444
+ 1.75e+10Hz 0.0038386 0.0093943
+ 1.76e+10Hz 0.00384497 0.00944414
+ 1.77e+10Hz 0.00385132 0.00949398
+ 1.78e+10Hz 0.00385767 0.0095438
+ 1.79e+10Hz 0.00386401 0.0095936
+ 1.8e+10Hz 0.00387034 0.00964339
+ 1.81e+10Hz 0.00387666 0.00969317
+ 1.82e+10Hz 0.00388297 0.00974294
+ 1.83e+10Hz 0.00388928 0.0097927
+ 1.84e+10Hz 0.00389557 0.00984245
+ 1.85e+10Hz 0.00390186 0.00989219
+ 1.86e+10Hz 0.00390814 0.00994192
+ 1.87e+10Hz 0.00391442 0.00999163
+ 1.88e+10Hz 0.00392069 0.0100413
+ 1.89e+10Hz 0.00392695 0.0100911
+ 1.9e+10Hz 0.0039332 0.0101407
+ 1.91e+10Hz 0.00393945 0.0101904
+ 1.92e+10Hz 0.00394569 0.0102401
+ 1.93e+10Hz 0.00395193 0.0102898
+ 1.94e+10Hz 0.00395816 0.0103395
+ 1.95e+10Hz 0.00396439 0.0103891
+ 1.96e+10Hz 0.00397061 0.0104388
+ 1.97e+10Hz 0.00397683 0.0104884
+ 1.98e+10Hz 0.00398304 0.0105381
+ 1.99e+10Hz 0.00398925 0.0105877
+ 2e+10Hz 0.00399545 0.0106374
+ 2.01e+10Hz 0.00400165 0.010687
+ 2.02e+10Hz 0.00400785 0.0107366
+ 2.03e+10Hz 0.00401404 0.0107862
+ 2.04e+10Hz 0.00402023 0.0108359
+ 2.05e+10Hz 0.00402643 0.0108855
+ 2.06e+10Hz 0.00403261 0.0109351
+ 2.07e+10Hz 0.0040388 0.0109847
+ 2.08e+10Hz 0.00404498 0.0110344
+ 2.09e+10Hz 0.00405117 0.011084
+ 2.1e+10Hz 0.00405735 0.0111336
+ 2.11e+10Hz 0.00406353 0.0111832
+ 2.12e+10Hz 0.00406971 0.0112328
+ 2.13e+10Hz 0.00407589 0.0112825
+ 2.14e+10Hz 0.00408208 0.0113321
+ 2.15e+10Hz 0.00408826 0.0113817
+ 2.16e+10Hz 0.00409444 0.0114313
+ 2.17e+10Hz 0.00410063 0.0114809
+ 2.18e+10Hz 0.00410682 0.0115306
+ 2.19e+10Hz 0.00411301 0.0115802
+ 2.2e+10Hz 0.0041192 0.0116298
+ 2.21e+10Hz 0.00412539 0.0116794
+ 2.22e+10Hz 0.00413159 0.0117291
+ 2.23e+10Hz 0.00413779 0.0117787
+ 2.24e+10Hz 0.004144 0.0118283
+ 2.25e+10Hz 0.0041502 0.011878
+ 2.26e+10Hz 0.00415642 0.0119276
+ 2.27e+10Hz 0.00416263 0.0119773
+ 2.28e+10Hz 0.00416886 0.0120269
+ 2.29e+10Hz 0.00417508 0.0120766
+ 2.3e+10Hz 0.00418132 0.0121262
+ 2.31e+10Hz 0.00418756 0.0121759
+ 2.32e+10Hz 0.0041938 0.0122255
+ 2.33e+10Hz 0.00420005 0.0122752
+ 2.34e+10Hz 0.00420631 0.0123248
+ 2.35e+10Hz 0.00421258 0.0123745
+ 2.36e+10Hz 0.00421885 0.0124242
+ 2.37e+10Hz 0.00422513 0.0124738
+ 2.38e+10Hz 0.00423142 0.0125235
+ 2.39e+10Hz 0.00423772 0.0125732
+ 2.4e+10Hz 0.00424402 0.0126229
+ 2.41e+10Hz 0.00425034 0.0126726
+ 2.42e+10Hz 0.00425666 0.0127223
+ 2.43e+10Hz 0.004263 0.012772
+ 2.44e+10Hz 0.00426934 0.0128217
+ 2.45e+10Hz 0.00427569 0.0128714
+ 2.46e+10Hz 0.00428206 0.0129211
+ 2.47e+10Hz 0.00428843 0.0129708
+ 2.48e+10Hz 0.00429482 0.0130205
+ 2.49e+10Hz 0.00430121 0.0130703
+ 2.5e+10Hz 0.00430762 0.01312
+ 2.51e+10Hz 0.00431404 0.0131697
+ 2.52e+10Hz 0.00432047 0.0132194
+ 2.53e+10Hz 0.00432692 0.0132692
+ 2.54e+10Hz 0.00433337 0.0133189
+ 2.55e+10Hz 0.00433984 0.0133687
+ 2.56e+10Hz 0.00434632 0.0134184
+ 2.57e+10Hz 0.00435282 0.0134682
+ 2.58e+10Hz 0.00435933 0.0135179
+ 2.59e+10Hz 0.00436585 0.0135677
+ 2.6e+10Hz 0.00437239 0.0136174
+ 2.61e+10Hz 0.00437894 0.0136672
+ 2.62e+10Hz 0.0043855 0.013717
+ 2.63e+10Hz 0.00439208 0.0137668
+ 2.64e+10Hz 0.00439867 0.0138165
+ 2.65e+10Hz 0.00440528 0.0138663
+ 2.66e+10Hz 0.00441191 0.0139161
+ 2.67e+10Hz 0.00441855 0.0139659
+ 2.68e+10Hz 0.0044252 0.0140157
+ 2.69e+10Hz 0.00443187 0.0140655
+ 2.7e+10Hz 0.00443856 0.0141153
+ 2.71e+10Hz 0.00444526 0.0141651
+ 2.72e+10Hz 0.00445198 0.0142149
+ 2.73e+10Hz 0.00445872 0.0142647
+ 2.74e+10Hz 0.00446547 0.0143145
+ 2.75e+10Hz 0.00447224 0.0143643
+ 2.76e+10Hz 0.00447903 0.0144141
+ 2.77e+10Hz 0.00448583 0.0144639
+ 2.78e+10Hz 0.00449265 0.0145137
+ 2.79e+10Hz 0.00449949 0.0145635
+ 2.8e+10Hz 0.00450635 0.0146133
+ 2.81e+10Hz 0.00451322 0.0146632
+ 2.82e+10Hz 0.00452011 0.014713
+ 2.83e+10Hz 0.00452702 0.0147628
+ 2.84e+10Hz 0.00453395 0.0148126
+ 2.85e+10Hz 0.0045409 0.0148624
+ 2.86e+10Hz 0.00454786 0.0149123
+ 2.87e+10Hz 0.00455485 0.0149621
+ 2.88e+10Hz 0.00456185 0.0150119
+ 2.89e+10Hz 0.00456887 0.0150617
+ 2.9e+10Hz 0.00457591 0.0151116
+ 2.91e+10Hz 0.00458297 0.0151614
+ 2.92e+10Hz 0.00459004 0.0152112
+ 2.93e+10Hz 0.00459714 0.015261
+ 2.94e+10Hz 0.00460426 0.0153109
+ 2.95e+10Hz 0.00461139 0.0153607
+ 2.96e+10Hz 0.00461855 0.0154105
+ 2.97e+10Hz 0.00462572 0.0154603
+ 2.98e+10Hz 0.00463291 0.0155102
+ 2.99e+10Hz 0.00464013 0.01556
+ 3e+10Hz 0.00464736 0.0156098
+ 3.01e+10Hz 0.00465461 0.0156596
+ 3.02e+10Hz 0.00466189 0.0157094
+ 3.03e+10Hz 0.00466918 0.0157593
+ 3.04e+10Hz 0.00467649 0.0158091
+ 3.05e+10Hz 0.00468382 0.0158589
+ 3.06e+10Hz 0.00469118 0.0159087
+ 3.07e+10Hz 0.00469855 0.0159585
+ 3.08e+10Hz 0.00470594 0.0160083
+ 3.09e+10Hz 0.00471335 0.0160581
+ 3.1e+10Hz 0.00472078 0.0161079
+ 3.11e+10Hz 0.00472824 0.0161577
+ 3.12e+10Hz 0.00473571 0.0162075
+ 3.13e+10Hz 0.0047432 0.0162573
+ 3.14e+10Hz 0.00475071 0.0163071
+ 3.15e+10Hz 0.00475825 0.0163569
+ 3.16e+10Hz 0.0047658 0.0164067
+ 3.17e+10Hz 0.00477337 0.0164565
+ 3.18e+10Hz 0.00478097 0.0165062
+ 3.19e+10Hz 0.00478858 0.016556
+ 3.2e+10Hz 0.00479622 0.0166058
+ 3.21e+10Hz 0.00480387 0.0166555
+ 3.22e+10Hz 0.00481154 0.0167053
+ 3.23e+10Hz 0.00481924 0.0167551
+ 3.24e+10Hz 0.00482695 0.0168048
+ 3.25e+10Hz 0.00483469 0.0168546
+ 3.26e+10Hz 0.00484244 0.0169043
+ 3.27e+10Hz 0.00485021 0.016954
+ 3.28e+10Hz 0.00485801 0.0170038
+ 3.29e+10Hz 0.00486582 0.0170535
+ 3.3e+10Hz 0.00487366 0.0171032
+ 3.31e+10Hz 0.00488151 0.017153
+ 3.32e+10Hz 0.00488938 0.0172027
+ 3.33e+10Hz 0.00489728 0.0172524
+ 3.34e+10Hz 0.00490519 0.0173021
+ 3.35e+10Hz 0.00491312 0.0173518
+ 3.36e+10Hz 0.00492108 0.0174015
+ 3.37e+10Hz 0.00492905 0.0174512
+ 3.38e+10Hz 0.00493704 0.0175008
+ 3.39e+10Hz 0.00494505 0.0175505
+ 3.4e+10Hz 0.00495308 0.0176002
+ 3.41e+10Hz 0.00496113 0.0176499
+ 3.42e+10Hz 0.0049692 0.0176995
+ 3.43e+10Hz 0.00497729 0.0177492
+ 3.44e+10Hz 0.0049854 0.0177988
+ 3.45e+10Hz 0.00499353 0.0178484
+ 3.46e+10Hz 0.00500167 0.0178981
+ 3.47e+10Hz 0.00500984 0.0179477
+ 3.48e+10Hz 0.00501802 0.0179973
+ 3.49e+10Hz 0.00502622 0.0180469
+ 3.5e+10Hz 0.00503445 0.0180965
+ 3.51e+10Hz 0.00504268 0.0181461
+ 3.52e+10Hz 0.00505094 0.0181957
+ 3.53e+10Hz 0.00505922 0.0182453
+ 3.54e+10Hz 0.00506752 0.0182949
+ 3.55e+10Hz 0.00507583 0.0183445
+ 3.56e+10Hz 0.00508416 0.018394
+ 3.57e+10Hz 0.00509252 0.0184436
+ 3.58e+10Hz 0.00510089 0.0184931
+ 3.59e+10Hz 0.00510927 0.0185427
+ 3.6e+10Hz 0.00511768 0.0185922
+ 3.61e+10Hz 0.0051261 0.0186417
+ 3.62e+10Hz 0.00513454 0.0186912
+ 3.63e+10Hz 0.005143 0.0187408
+ 3.64e+10Hz 0.00515148 0.0187903
+ 3.65e+10Hz 0.00515997 0.0188397
+ 3.66e+10Hz 0.00516848 0.0188892
+ 3.67e+10Hz 0.00517701 0.0189387
+ 3.68e+10Hz 0.00518556 0.0189882
+ 3.69e+10Hz 0.00519412 0.0190376
+ 3.7e+10Hz 0.0052027 0.0190871
+ 3.71e+10Hz 0.0052113 0.0191366
+ 3.72e+10Hz 0.00521991 0.019186
+ 3.73e+10Hz 0.00522855 0.0192354
+ 3.74e+10Hz 0.00523719 0.0192848
+ 3.75e+10Hz 0.00524586 0.0193343
+ 3.76e+10Hz 0.00525454 0.0193837
+ 3.77e+10Hz 0.00526324 0.0194331
+ 3.78e+10Hz 0.00527195 0.0194825
+ 3.79e+10Hz 0.00528069 0.0195319
+ 3.8e+10Hz 0.00528943 0.0195812
+ 3.81e+10Hz 0.0052982 0.0196306
+ 3.82e+10Hz 0.00530698 0.01968
+ 3.83e+10Hz 0.00531577 0.0197293
+ 3.84e+10Hz 0.00532458 0.0197787
+ 3.85e+10Hz 0.00533341 0.019828
+ 3.86e+10Hz 0.00534226 0.0198773
+ 3.87e+10Hz 0.00535112 0.0199267
+ 3.88e+10Hz 0.00535999 0.019976
+ 3.89e+10Hz 0.00536888 0.0200253
+ 3.9e+10Hz 0.00537779 0.0200746
+ 3.91e+10Hz 0.00538671 0.0201239
+ 3.92e+10Hz 0.00539565 0.0201731
+ 3.93e+10Hz 0.0054046 0.0202224
+ 3.94e+10Hz 0.00541357 0.0202717
+ 3.95e+10Hz 0.00542255 0.0203209
+ 3.96e+10Hz 0.00543155 0.0203702
+ 3.97e+10Hz 0.00544056 0.0204194
+ 3.98e+10Hz 0.00544959 0.0204687
+ 3.99e+10Hz 0.00545863 0.0205179
+ 4e+10Hz 0.00546769 0.0205671
+ 4.01e+10Hz 0.00547676 0.0206163
+ 4.02e+10Hz 0.00548585 0.0206655
+ 4.03e+10Hz 0.00549495 0.0207147
+ 4.04e+10Hz 0.00550407 0.0207639
+ 4.05e+10Hz 0.0055132 0.0208131
+ 4.06e+10Hz 0.00552234 0.0208623
+ 4.07e+10Hz 0.0055315 0.0209114
+ 4.08e+10Hz 0.00554068 0.0209606
+ 4.09e+10Hz 0.00554986 0.0210097
+ 4.1e+10Hz 0.00555906 0.0210589
+ 4.11e+10Hz 0.00556828 0.021108
+ 4.12e+10Hz 0.00557751 0.0211571
+ 4.13e+10Hz 0.00558675 0.0212063
+ 4.14e+10Hz 0.00559601 0.0212554
+ 4.15e+10Hz 0.00560528 0.0213045
+ 4.16e+10Hz 0.00561457 0.0213536
+ 4.17e+10Hz 0.00562387 0.0214027
+ 4.18e+10Hz 0.00563318 0.0214518
+ 4.19e+10Hz 0.00564251 0.0215009
+ 4.2e+10Hz 0.00565185 0.0215499
+ 4.21e+10Hz 0.0056612 0.021599
+ 4.22e+10Hz 0.00567057 0.021648
+ 4.23e+10Hz 0.00567995 0.0216971
+ 4.24e+10Hz 0.00568935 0.0217461
+ 4.25e+10Hz 0.00569876 0.0217952
+ 4.26e+10Hz 0.00570818 0.0218442
+ 4.27e+10Hz 0.00571761 0.0218932
+ 4.28e+10Hz 0.00572706 0.0219423
+ 4.29e+10Hz 0.00573653 0.0219913
+ 4.3e+10Hz 0.005746 0.0220403
+ 4.31e+10Hz 0.00575549 0.0220893
+ 4.32e+10Hz 0.00576499 0.0221383
+ 4.33e+10Hz 0.00577451 0.0221873
+ 4.34e+10Hz 0.00578403 0.0222363
+ 4.35e+10Hz 0.00579358 0.0222852
+ 4.36e+10Hz 0.00580313 0.0223342
+ 4.37e+10Hz 0.0058127 0.0223832
+ 4.38e+10Hz 0.00582228 0.0224321
+ 4.39e+10Hz 0.00583188 0.0224811
+ 4.4e+10Hz 0.00584148 0.02253
+ 4.41e+10Hz 0.0058511 0.022579
+ 4.42e+10Hz 0.00586074 0.0226279
+ 4.43e+10Hz 0.00587038 0.0226768
+ 4.44e+10Hz 0.00588004 0.0227258
+ 4.45e+10Hz 0.00588972 0.0227747
+ 4.46e+10Hz 0.0058994 0.0228236
+ 4.47e+10Hz 0.0059091 0.0228725
+ 4.48e+10Hz 0.00591882 0.0229214
+ 4.49e+10Hz 0.00592854 0.0229703
+ 4.5e+10Hz 0.00593828 0.0230192
+ 4.51e+10Hz 0.00594803 0.0230681
+ 4.52e+10Hz 0.0059578 0.023117
+ 4.53e+10Hz 0.00596757 0.0231659
+ 4.54e+10Hz 0.00597737 0.0232147
+ 4.55e+10Hz 0.00598717 0.0232636
+ 4.56e+10Hz 0.00599699 0.0233125
+ 4.57e+10Hz 0.00600682 0.0233613
+ 4.58e+10Hz 0.00601666 0.0234102
+ 4.59e+10Hz 0.00602652 0.023459
+ 4.6e+10Hz 0.00603639 0.0235079
+ 4.61e+10Hz 0.00604627 0.0235567
+ 4.62e+10Hz 0.00605617 0.0236055
+ 4.63e+10Hz 0.00606608 0.0236544
+ 4.64e+10Hz 0.006076 0.0237032
+ 4.65e+10Hz 0.00608594 0.023752
+ 4.66e+10Hz 0.00609589 0.0238008
+ 4.67e+10Hz 0.00610585 0.0238497
+ 4.68e+10Hz 0.00611583 0.0238985
+ 4.69e+10Hz 0.00612582 0.0239473
+ 4.7e+10Hz 0.00613582 0.0239961
+ 4.71e+10Hz 0.00614584 0.0240449
+ 4.72e+10Hz 0.00615587 0.0240937
+ 4.73e+10Hz 0.00616591 0.0241425
+ 4.74e+10Hz 0.00617597 0.0241913
+ 4.75e+10Hz 0.00618604 0.02424
+ 4.76e+10Hz 0.00619612 0.0242888
+ 4.77e+10Hz 0.00620622 0.0243376
+ 4.78e+10Hz 0.00621633 0.0243864
+ 4.79e+10Hz 0.00622646 0.0244351
+ 4.8e+10Hz 0.0062366 0.0244839
+ 4.81e+10Hz 0.00624675 0.0245327
+ 4.82e+10Hz 0.00625692 0.0245814
+ 4.83e+10Hz 0.0062671 0.0246302
+ 4.84e+10Hz 0.00627729 0.0246789
+ 4.85e+10Hz 0.0062875 0.0247277
+ 4.86e+10Hz 0.00629773 0.0247764
+ 4.87e+10Hz 0.00630796 0.0248252
+ 4.88e+10Hz 0.00631822 0.0248739
+ 4.89e+10Hz 0.00632848 0.0249226
+ 4.9e+10Hz 0.00633876 0.0249714
+ 4.91e+10Hz 0.00634905 0.0250201
+ 4.92e+10Hz 0.00635936 0.0250688
+ 4.93e+10Hz 0.00636968 0.0251175
+ 4.94e+10Hz 0.00638002 0.0251663
+ 4.95e+10Hz 0.00639037 0.025215
+ 4.96e+10Hz 0.00640074 0.0252637
+ 4.97e+10Hz 0.00641112 0.0253124
+ 4.98e+10Hz 0.00642151 0.0253611
+ 4.99e+10Hz 0.00643192 0.0254098
+ 5e+10Hz 0.00644235 0.0254585
+ 5.01e+10Hz 0.00645279 0.0255072
+ 5.02e+10Hz 0.00646324 0.0255559
+ 5.03e+10Hz 0.00647371 0.0256046
+ 5.04e+10Hz 0.00648419 0.0256533
+ 5.05e+10Hz 0.00649469 0.025702
+ 5.06e+10Hz 0.00650521 0.0257506
+ 5.07e+10Hz 0.00651573 0.0257993
+ 5.08e+10Hz 0.00652628 0.025848
+ 5.09e+10Hz 0.00653684 0.0258967
+ 5.1e+10Hz 0.00654741 0.0259453
+ 5.11e+10Hz 0.006558 0.025994
+ 5.12e+10Hz 0.00656861 0.0260427
+ 5.13e+10Hz 0.00657923 0.0260913
+ 5.14e+10Hz 0.00658986 0.02614
+ 5.15e+10Hz 0.00660051 0.0261886
+ 5.16e+10Hz 0.00661118 0.0262373
+ 5.17e+10Hz 0.00662186 0.0262859
+ 5.18e+10Hz 0.00663256 0.0263346
+ 5.19e+10Hz 0.00664328 0.0263832
+ 5.2e+10Hz 0.00665401 0.0264319
+ 5.21e+10Hz 0.00666475 0.0264805
+ 5.22e+10Hz 0.00667551 0.0265292
+ 5.23e+10Hz 0.00668629 0.0265778
+ 5.24e+10Hz 0.00669708 0.0266264
+ 5.25e+10Hz 0.00670789 0.026675
+ 5.26e+10Hz 0.00671872 0.0267237
+ 5.27e+10Hz 0.00672956 0.0267723
+ 5.28e+10Hz 0.00674042 0.0268209
+ 5.29e+10Hz 0.00675129 0.0268695
+ 5.3e+10Hz 0.00676219 0.0269181
+ 5.31e+10Hz 0.00677309 0.0269668
+ 5.32e+10Hz 0.00678402 0.0270154
+ 5.33e+10Hz 0.00679496 0.027064
+ 5.34e+10Hz 0.00680591 0.0271126
+ 5.35e+10Hz 0.00681689 0.0271612
+ 5.36e+10Hz 0.00682788 0.0272098
+ 5.37e+10Hz 0.00683888 0.0272583
+ 5.38e+10Hz 0.00684991 0.0273069
+ 5.39e+10Hz 0.00686095 0.0273555
+ 5.4e+10Hz 0.006872 0.0274041
+ 5.41e+10Hz 0.00688308 0.0274527
+ 5.42e+10Hz 0.00689417 0.0275013
+ 5.43e+10Hz 0.00690527 0.0275498
+ 5.44e+10Hz 0.0069164 0.0275984
+ 5.45e+10Hz 0.00692754 0.027647
+ 5.46e+10Hz 0.0069387 0.0276955
+ 5.47e+10Hz 0.00694988 0.0277441
+ 5.48e+10Hz 0.00696107 0.0277926
+ 5.49e+10Hz 0.00697228 0.0278412
+ 5.5e+10Hz 0.00698351 0.0278898
+ 5.51e+10Hz 0.00699476 0.0279383
+ 5.52e+10Hz 0.00700602 0.0279868
+ 5.53e+10Hz 0.0070173 0.0280354
+ 5.54e+10Hz 0.0070286 0.0280839
+ 5.55e+10Hz 0.00703991 0.0281324
+ 5.56e+10Hz 0.00705124 0.028181
+ 5.57e+10Hz 0.00706259 0.0282295
+ 5.58e+10Hz 0.00707396 0.028278
+ 5.59e+10Hz 0.00708535 0.0283265
+ 5.6e+10Hz 0.00709675 0.028375
+ 5.61e+10Hz 0.00710817 0.0284236
+ 5.62e+10Hz 0.00711961 0.0284721
+ 5.63e+10Hz 0.00713107 0.0285206
+ 5.64e+10Hz 0.00714254 0.0285691
+ 5.65e+10Hz 0.00715404 0.0286176
+ 5.66e+10Hz 0.00716554 0.028666
+ 5.67e+10Hz 0.00717707 0.0287145
+ 5.68e+10Hz 0.00718862 0.028763
+ 5.69e+10Hz 0.00720018 0.0288115
+ 5.7e+10Hz 0.00721177 0.02886
+ 5.71e+10Hz 0.00722337 0.0289084
+ 5.72e+10Hz 0.00723498 0.0289569
+ 5.73e+10Hz 0.00724662 0.0290054
+ 5.74e+10Hz 0.00725827 0.0290538
+ 5.75e+10Hz 0.00726995 0.0291023
+ 5.76e+10Hz 0.00728164 0.0291507
+ 5.77e+10Hz 0.00729335 0.0291992
+ 5.78e+10Hz 0.00730508 0.0292476
+ 5.79e+10Hz 0.00731682 0.029296
+ 5.8e+10Hz 0.00732858 0.0293445
+ 5.81e+10Hz 0.00734037 0.0293929
+ 5.82e+10Hz 0.00735217 0.0294413
+ 5.83e+10Hz 0.00736398 0.0294897
+ 5.84e+10Hz 0.00737582 0.0295381
+ 5.85e+10Hz 0.00738768 0.0295865
+ 5.86e+10Hz 0.00739955 0.0296349
+ 5.87e+10Hz 0.00741144 0.0296833
+ 5.88e+10Hz 0.00742335 0.0297317
+ 5.89e+10Hz 0.00743528 0.0297801
+ 5.9e+10Hz 0.00744723 0.0298285
+ 5.91e+10Hz 0.00745919 0.0298768
+ 5.92e+10Hz 0.00747118 0.0299252
+ 5.93e+10Hz 0.00748318 0.0299736
+ 5.94e+10Hz 0.0074952 0.0300219
+ 5.95e+10Hz 0.00750724 0.0300703
+ 5.96e+10Hz 0.0075193 0.0301186
+ 5.97e+10Hz 0.00753137 0.030167
+ 5.98e+10Hz 0.00754347 0.0302153
+ 5.99e+10Hz 0.00755558 0.0302636
+ 6e+10Hz 0.00756771 0.030312
+ 6.01e+10Hz 0.00757986 0.0303603
+ 6.02e+10Hz 0.00759203 0.0304086
+ 6.03e+10Hz 0.00760422 0.0304569
+ 6.04e+10Hz 0.00761642 0.0305052
+ 6.05e+10Hz 0.00762865 0.0305535
+ 6.06e+10Hz 0.00764089 0.0306018
+ 6.07e+10Hz 0.00765315 0.0306501
+ 6.08e+10Hz 0.00766543 0.0306984
+ 6.09e+10Hz 0.00767772 0.0307466
+ 6.1e+10Hz 0.00769004 0.0307949
+ 6.11e+10Hz 0.00770237 0.0308432
+ 6.12e+10Hz 0.00771473 0.0308914
+ 6.13e+10Hz 0.0077271 0.0309397
+ 6.14e+10Hz 0.00773949 0.0309879
+ 6.15e+10Hz 0.00775189 0.0310361
+ 6.16e+10Hz 0.00776432 0.0310844
+ 6.17e+10Hz 0.00777676 0.0311326
+ 6.18e+10Hz 0.00778923 0.0311808
+ 6.19e+10Hz 0.00780171 0.031229
+ 6.2e+10Hz 0.00781421 0.0312772
+ 6.21e+10Hz 0.00782672 0.0313254
+ 6.22e+10Hz 0.00783926 0.0313736
+ 6.23e+10Hz 0.00785181 0.0314218
+ 6.24e+10Hz 0.00786439 0.03147
+ 6.25e+10Hz 0.00787698 0.0315181
+ 6.26e+10Hz 0.00788958 0.0315663
+ 6.27e+10Hz 0.00790221 0.0316145
+ 6.28e+10Hz 0.00791486 0.0316626
+ 6.29e+10Hz 0.00792752 0.0317108
+ 6.3e+10Hz 0.0079402 0.0317589
+ 6.31e+10Hz 0.0079529 0.031807
+ 6.32e+10Hz 0.00796562 0.0318551
+ 6.33e+10Hz 0.00797835 0.0319033
+ 6.34e+10Hz 0.00799111 0.0319514
+ 6.35e+10Hz 0.00800388 0.0319995
+ 6.36e+10Hz 0.00801667 0.0320476
+ 6.37e+10Hz 0.00802947 0.0320956
+ 6.38e+10Hz 0.0080423 0.0321437
+ 6.39e+10Hz 0.00805514 0.0321918
+ 6.4e+10Hz 0.008068 0.0322399
+ 6.41e+10Hz 0.00808088 0.0322879
+ 6.42e+10Hz 0.00809378 0.032336
+ 6.43e+10Hz 0.00810669 0.032384
+ 6.44e+10Hz 0.00811963 0.032432
+ 6.45e+10Hz 0.00813258 0.0324801
+ 6.46e+10Hz 0.00814554 0.0325281
+ 6.47e+10Hz 0.00815853 0.0325761
+ 6.48e+10Hz 0.00817153 0.0326241
+ 6.49e+10Hz 0.00818455 0.0326721
+ 6.5e+10Hz 0.00819759 0.0327201
+ 6.51e+10Hz 0.00821065 0.0327681
+ 6.52e+10Hz 0.00822372 0.0328161
+ 6.53e+10Hz 0.00823681 0.032864
+ 6.54e+10Hz 0.00824992 0.032912
+ 6.55e+10Hz 0.00826305 0.03296
+ 6.56e+10Hz 0.00827619 0.0330079
+ 6.57e+10Hz 0.00828935 0.0330558
+ 6.58e+10Hz 0.00830253 0.0331038
+ 6.59e+10Hz 0.00831572 0.0331517
+ 6.6e+10Hz 0.00832894 0.0331996
+ 6.61e+10Hz 0.00834217 0.0332475
+ 6.62e+10Hz 0.00835541 0.0332954
+ 6.63e+10Hz 0.00836868 0.0333433
+ 6.64e+10Hz 0.00838196 0.0333912
+ 6.65e+10Hz 0.00839526 0.0334391
+ 6.66e+10Hz 0.00840857 0.0334869
+ 6.67e+10Hz 0.00842191 0.0335348
+ 6.68e+10Hz 0.00843526 0.0335827
+ 6.69e+10Hz 0.00844862 0.0336305
+ 6.7e+10Hz 0.00846201 0.0336784
+ 6.71e+10Hz 0.00847541 0.0337262
+ 6.72e+10Hz 0.00848883 0.033774
+ 6.73e+10Hz 0.00850226 0.0338218
+ 6.74e+10Hz 0.00851572 0.0338696
+ 6.75e+10Hz 0.00852918 0.0339174
+ 6.76e+10Hz 0.00854267 0.0339652
+ 6.77e+10Hz 0.00855617 0.034013
+ 6.78e+10Hz 0.00856969 0.0340608
+ 6.79e+10Hz 0.00858323 0.0341086
+ 6.8e+10Hz 0.00859678 0.0341563
+ 6.81e+10Hz 0.00861035 0.0342041
+ 6.82e+10Hz 0.00862393 0.0342518
+ 6.83e+10Hz 0.00863754 0.0342995
+ 6.84e+10Hz 0.00865115 0.0343473
+ 6.85e+10Hz 0.00866479 0.034395
+ 6.86e+10Hz 0.00867844 0.0344427
+ 6.87e+10Hz 0.00869211 0.0344904
+ 6.88e+10Hz 0.0087058 0.0345381
+ 6.89e+10Hz 0.0087195 0.0345858
+ 6.9e+10Hz 0.00873321 0.0346335
+ 6.91e+10Hz 0.00874695 0.0346812
+ 6.92e+10Hz 0.0087607 0.0347288
+ 6.93e+10Hz 0.00877447 0.0347765
+ 6.94e+10Hz 0.00878825 0.0348242
+ 6.95e+10Hz 0.00880205 0.0348718
+ 6.96e+10Hz 0.00881586 0.0349194
+ 6.97e+10Hz 0.0088297 0.0349671
+ 6.98e+10Hz 0.00884354 0.0350147
+ 6.99e+10Hz 0.00885741 0.0350623
+ 7e+10Hz 0.00887129 0.0351099
+ 7.01e+10Hz 0.00888519 0.0351575
+ 7.02e+10Hz 0.0088991 0.0352051
+ 7.03e+10Hz 0.00891303 0.0352527
+ 7.04e+10Hz 0.00892697 0.0353003
+ 7.05e+10Hz 0.00894093 0.0353479
+ 7.06e+10Hz 0.00895491 0.0353954
+ 7.07e+10Hz 0.0089689 0.035443
+ 7.08e+10Hz 0.00898291 0.0354905
+ 7.09e+10Hz 0.00899694 0.0355381
+ 7.1e+10Hz 0.00901098 0.0355856
+ 7.11e+10Hz 0.00902503 0.0356331
+ 7.12e+10Hz 0.00903911 0.0356806
+ 7.13e+10Hz 0.0090532 0.0357281
+ 7.14e+10Hz 0.0090673 0.0357756
+ 7.15e+10Hz 0.00908142 0.0358231
+ 7.16e+10Hz 0.00909556 0.0358706
+ 7.17e+10Hz 0.00910971 0.0359181
+ 7.18e+10Hz 0.00912388 0.0359656
+ 7.19e+10Hz 0.00913806 0.036013
+ 7.2e+10Hz 0.00915226 0.0360605
+ 7.21e+10Hz 0.00916648 0.036108
+ 7.22e+10Hz 0.00918071 0.0361554
+ 7.23e+10Hz 0.00919496 0.0362028
+ 7.24e+10Hz 0.00920922 0.0362503
+ 7.25e+10Hz 0.0092235 0.0362977
+ 7.26e+10Hz 0.00923779 0.0363451
+ 7.27e+10Hz 0.0092521 0.0363925
+ 7.28e+10Hz 0.00926643 0.0364399
+ 7.29e+10Hz 0.00928077 0.0364873
+ 7.3e+10Hz 0.00929513 0.0365347
+ 7.31e+10Hz 0.0093095 0.0365821
+ 7.32e+10Hz 0.00932389 0.0366295
+ 7.33e+10Hz 0.00933829 0.0366768
+ 7.34e+10Hz 0.00935271 0.0367242
+ 7.35e+10Hz 0.00936715 0.0367716
+ 7.36e+10Hz 0.0093816 0.0368189
+ 7.37e+10Hz 0.00939607 0.0368662
+ 7.38e+10Hz 0.00941055 0.0369136
+ 7.39e+10Hz 0.00942505 0.0369609
+ 7.4e+10Hz 0.00943957 0.0370082
+ 7.41e+10Hz 0.0094541 0.0370555
+ 7.42e+10Hz 0.00946864 0.0371028
+ 7.43e+10Hz 0.0094832 0.0371501
+ 7.44e+10Hz 0.00949778 0.0371974
+ 7.45e+10Hz 0.00951237 0.0372447
+ 7.46e+10Hz 0.00952698 0.037292
+ 7.47e+10Hz 0.00954161 0.0373393
+ 7.48e+10Hz 0.00955625 0.0373865
+ 7.49e+10Hz 0.0095709 0.0374338
+ 7.5e+10Hz 0.00958558 0.037481
+ 7.51e+10Hz 0.00960026 0.0375283
+ 7.52e+10Hz 0.00961497 0.0375755
+ 7.53e+10Hz 0.00962969 0.0376228
+ 7.54e+10Hz 0.00964442 0.03767
+ 7.55e+10Hz 0.00965917 0.0377172
+ 7.56e+10Hz 0.00967394 0.0377644
+ 7.57e+10Hz 0.00968872 0.0378116
+ 7.58e+10Hz 0.00970352 0.0378588
+ 7.59e+10Hz 0.00971833 0.037906
+ 7.6e+10Hz 0.00973316 0.0379532
+ 7.61e+10Hz 0.00974801 0.0380004
+ 7.62e+10Hz 0.00976287 0.0380476
+ 7.63e+10Hz 0.00977774 0.0380947
+ 7.64e+10Hz 0.00979264 0.0381419
+ 7.65e+10Hz 0.00980755 0.0381891
+ 7.66e+10Hz 0.00982247 0.0382362
+ 7.67e+10Hz 0.00983741 0.0382834
+ 7.68e+10Hz 0.00985237 0.0383305
+ 7.69e+10Hz 0.00986734 0.0383776
+ 7.7e+10Hz 0.00988233 0.0384248
+ 7.71e+10Hz 0.00989734 0.0384719
+ 7.72e+10Hz 0.00991236 0.038519
+ 7.73e+10Hz 0.0099274 0.0385661
+ 7.74e+10Hz 0.00994245 0.0386132
+ 7.75e+10Hz 0.00995752 0.0386603
+ 7.76e+10Hz 0.0099726 0.0387074
+ 7.77e+10Hz 0.0099877 0.0387545
+ 7.78e+10Hz 0.0100028 0.0388015
+ 7.79e+10Hz 0.010018 0.0388486
+ 7.8e+10Hz 0.0100331 0.0388957
+ 7.81e+10Hz 0.0100483 0.0389427
+ 7.82e+10Hz 0.0100635 0.0389898
+ 7.83e+10Hz 0.0100786 0.0390368
+ 7.84e+10Hz 0.0100939 0.0390839
+ 7.85e+10Hz 0.0101091 0.0391309
+ 7.86e+10Hz 0.0101244 0.039178
+ 7.87e+10Hz 0.0101396 0.039225
+ 7.88e+10Hz 0.0101549 0.039272
+ 7.89e+10Hz 0.0101702 0.039319
+ 7.9e+10Hz 0.0101855 0.039366
+ 7.91e+10Hz 0.0102008 0.039413
+ 7.92e+10Hz 0.0102162 0.03946
+ 7.93e+10Hz 0.0102315 0.039507
+ 7.94e+10Hz 0.0102469 0.039554
+ 7.95e+10Hz 0.0102623 0.039601
+ 7.96e+10Hz 0.0102777 0.0396479
+ 7.97e+10Hz 0.0102932 0.0396949
+ 7.98e+10Hz 0.0103086 0.0397419
+ 7.99e+10Hz 0.0103241 0.0397888
+ 8e+10Hz 0.0103395 0.0398358
+ 8.01e+10Hz 0.010355 0.0398827
+ 8.02e+10Hz 0.0103706 0.0399296
+ 8.03e+10Hz 0.0103861 0.0399766
+ 8.04e+10Hz 0.0104016 0.0400235
+ 8.05e+10Hz 0.0104172 0.0400704
+ 8.06e+10Hz 0.0104328 0.0401173
+ 8.07e+10Hz 0.0104484 0.0401642
+ 8.08e+10Hz 0.010464 0.0402112
+ 8.09e+10Hz 0.0104796 0.040258
+ 8.1e+10Hz 0.0104953 0.0403049
+ 8.11e+10Hz 0.0105109 0.0403518
+ 8.12e+10Hz 0.0105266 0.0403987
+ 8.13e+10Hz 0.0105423 0.0404456
+ 8.14e+10Hz 0.010558 0.0404924
+ 8.15e+10Hz 0.0105738 0.0405393
+ 8.16e+10Hz 0.0105895 0.0405862
+ 8.17e+10Hz 0.0106053 0.040633
+ 8.18e+10Hz 0.0106211 0.0406798
+ 8.19e+10Hz 0.0106369 0.0407267
+ 8.2e+10Hz 0.0106527 0.0407735
+ 8.21e+10Hz 0.0106685 0.0408203
+ 8.22e+10Hz 0.0106844 0.0408672
+ 8.23e+10Hz 0.0107002 0.040914
+ 8.24e+10Hz 0.0107161 0.0409608
+ 8.25e+10Hz 0.010732 0.0410076
+ 8.26e+10Hz 0.010748 0.0410544
+ 8.27e+10Hz 0.0107639 0.0411012
+ 8.28e+10Hz 0.0107799 0.041148
+ 8.29e+10Hz 0.0107958 0.0411948
+ 8.3e+10Hz 0.0108118 0.0412415
+ 8.31e+10Hz 0.0108278 0.0412883
+ 8.32e+10Hz 0.0108439 0.041335
+ 8.33e+10Hz 0.0108599 0.0413818
+ 8.34e+10Hz 0.010876 0.0414286
+ 8.35e+10Hz 0.0108921 0.0414753
+ 8.36e+10Hz 0.0109082 0.041522
+ 8.37e+10Hz 0.0109243 0.0415688
+ 8.38e+10Hz 0.0109404 0.0416155
+ 8.39e+10Hz 0.0109566 0.0416622
+ 8.4e+10Hz 0.0109727 0.0417089
+ 8.41e+10Hz 0.0109889 0.0417556
+ 8.42e+10Hz 0.0110051 0.0418023
+ 8.43e+10Hz 0.0110213 0.041849
+ 8.44e+10Hz 0.0110376 0.0418957
+ 8.45e+10Hz 0.0110539 0.0419424
+ 8.46e+10Hz 0.0110701 0.0419891
+ 8.47e+10Hz 0.0110864 0.0420357
+ 8.48e+10Hz 0.0111027 0.0420824
+ 8.49e+10Hz 0.0111191 0.042129
+ 8.5e+10Hz 0.0111354 0.0421757
+ 8.51e+10Hz 0.0111518 0.0422223
+ 8.52e+10Hz 0.0111682 0.042269
+ 8.53e+10Hz 0.0111846 0.0423156
+ 8.54e+10Hz 0.011201 0.0423622
+ 8.55e+10Hz 0.0112174 0.0424088
+ 8.56e+10Hz 0.0112339 0.0424554
+ 8.57e+10Hz 0.0112504 0.042502
+ 8.58e+10Hz 0.0112669 0.0425486
+ 8.59e+10Hz 0.0112834 0.0425952
+ 8.6e+10Hz 0.0112999 0.0426418
+ 8.61e+10Hz 0.0113165 0.0426884
+ 8.62e+10Hz 0.011333 0.042735
+ 8.63e+10Hz 0.0113496 0.0427815
+ 8.64e+10Hz 0.0113662 0.0428281
+ 8.65e+10Hz 0.0113828 0.0428746
+ 8.66e+10Hz 0.0113995 0.0429212
+ 8.67e+10Hz 0.0114161 0.0429677
+ 8.68e+10Hz 0.0114328 0.0430142
+ 8.69e+10Hz 0.0114495 0.0430608
+ 8.7e+10Hz 0.0114662 0.0431073
+ 8.71e+10Hz 0.0114829 0.0431538
+ 8.72e+10Hz 0.0114997 0.0432003
+ 8.73e+10Hz 0.0115164 0.0432468
+ 8.74e+10Hz 0.0115332 0.0432932
+ 8.75e+10Hz 0.01155 0.0433397
+ 8.76e+10Hz 0.0115668 0.0433862
+ 8.77e+10Hz 0.0115837 0.0434327
+ 8.78e+10Hz 0.0116005 0.0434791
+ 8.79e+10Hz 0.0116174 0.0435256
+ 8.8e+10Hz 0.0116343 0.043572
+ 8.81e+10Hz 0.0116512 0.0436185
+ 8.82e+10Hz 0.0116682 0.0436649
+ 8.83e+10Hz 0.0116851 0.0437113
+ 8.84e+10Hz 0.0117021 0.0437577
+ 8.85e+10Hz 0.011719 0.0438041
+ 8.86e+10Hz 0.011736 0.0438505
+ 8.87e+10Hz 0.0117531 0.0438969
+ 8.88e+10Hz 0.0117701 0.0439433
+ 8.89e+10Hz 0.0117872 0.0439896
+ 8.9e+10Hz 0.0118043 0.044036
+ 8.91e+10Hz 0.0118213 0.0440824
+ 8.92e+10Hz 0.0118385 0.0441287
+ 8.93e+10Hz 0.0118556 0.0441751
+ 8.94e+10Hz 0.0118727 0.0442214
+ 8.95e+10Hz 0.0118899 0.0442677
+ 8.96e+10Hz 0.0119071 0.0443141
+ 8.97e+10Hz 0.0119243 0.0443604
+ 8.98e+10Hz 0.0119415 0.0444067
+ 8.99e+10Hz 0.0119588 0.044453
+ 9e+10Hz 0.011976 0.0444992
+ 9.01e+10Hz 0.0119933 0.0445455
+ 9.02e+10Hz 0.0120106 0.0445918
+ 9.03e+10Hz 0.0120279 0.0446381
+ 9.04e+10Hz 0.0120452 0.0446843
+ 9.05e+10Hz 0.0120626 0.0447306
+ 9.06e+10Hz 0.0120799 0.0447768
+ 9.07e+10Hz 0.0120973 0.044823
+ 9.08e+10Hz 0.0121147 0.0448692
+ 9.09e+10Hz 0.0121321 0.0449155
+ 9.1e+10Hz 0.0121496 0.0449617
+ 9.11e+10Hz 0.0121671 0.0450079
+ 9.12e+10Hz 0.0121845 0.0450541
+ 9.13e+10Hz 0.012202 0.0451002
+ 9.14e+10Hz 0.0122195 0.0451464
+ 9.15e+10Hz 0.012237 0.0451926
+ 9.16e+10Hz 0.0122546 0.0452387
+ 9.17e+10Hz 0.0122722 0.0452849
+ 9.18e+10Hz 0.0122897 0.045331
+ 9.19e+10Hz 0.0123073 0.0453771
+ 9.2e+10Hz 0.012325 0.0454233
+ 9.21e+10Hz 0.0123426 0.0454694
+ 9.22e+10Hz 0.0123602 0.0455155
+ 9.23e+10Hz 0.0123779 0.0455616
+ 9.24e+10Hz 0.0123956 0.0456076
+ 9.25e+10Hz 0.0124133 0.0456537
+ 9.26e+10Hz 0.012431 0.0456998
+ 9.27e+10Hz 0.0124488 0.0457459
+ 9.28e+10Hz 0.0124665 0.0457919
+ 9.29e+10Hz 0.0124843 0.045838
+ 9.3e+10Hz 0.0125021 0.045884
+ 9.31e+10Hz 0.0125199 0.04593
+ 9.32e+10Hz 0.0125378 0.045976
+ 9.33e+10Hz 0.0125556 0.046022
+ 9.34e+10Hz 0.0125735 0.046068
+ 9.35e+10Hz 0.0125913 0.046114
+ 9.36e+10Hz 0.0126092 0.04616
+ 9.37e+10Hz 0.0126272 0.046206
+ 9.38e+10Hz 0.0126451 0.0462519
+ 9.39e+10Hz 0.012663 0.0462979
+ 9.4e+10Hz 0.012681 0.0463438
+ 9.41e+10Hz 0.012699 0.0463897
+ 9.42e+10Hz 0.012717 0.0464357
+ 9.43e+10Hz 0.012735 0.0464816
+ 9.44e+10Hz 0.012753 0.0465275
+ 9.45e+10Hz 0.0127711 0.0465734
+ 9.46e+10Hz 0.0127892 0.0466193
+ 9.47e+10Hz 0.0128072 0.0466651
+ 9.48e+10Hz 0.0128253 0.046711
+ 9.49e+10Hz 0.0128435 0.0467569
+ 9.5e+10Hz 0.0128616 0.0468027
+ 9.51e+10Hz 0.0128798 0.0468486
+ 9.52e+10Hz 0.0128979 0.0468944
+ 9.53e+10Hz 0.0129161 0.0469402
+ 9.54e+10Hz 0.0129343 0.046986
+ 9.55e+10Hz 0.0129525 0.0470318
+ 9.56e+10Hz 0.0129708 0.0470776
+ 9.57e+10Hz 0.012989 0.0471234
+ 9.58e+10Hz 0.0130073 0.0471692
+ 9.59e+10Hz 0.0130256 0.047215
+ 9.6e+10Hz 0.0130439 0.0472607
+ 9.61e+10Hz 0.0130622 0.0473065
+ 9.62e+10Hz 0.0130805 0.0473522
+ 9.63e+10Hz 0.0130989 0.0473979
+ 9.64e+10Hz 0.0131173 0.0474436
+ 9.65e+10Hz 0.0131357 0.0474894
+ 9.66e+10Hz 0.0131541 0.0475351
+ 9.67e+10Hz 0.0131725 0.0475808
+ 9.68e+10Hz 0.0131909 0.0476264
+ 9.69e+10Hz 0.0132094 0.0476721
+ 9.7e+10Hz 0.0132278 0.0477178
+ 9.71e+10Hz 0.0132463 0.0477634
+ 9.72e+10Hz 0.0132648 0.0478091
+ 9.73e+10Hz 0.0132833 0.0478547
+ 9.74e+10Hz 0.0133019 0.0479003
+ 9.75e+10Hz 0.0133204 0.047946
+ 9.76e+10Hz 0.013339 0.0479916
+ 9.77e+10Hz 0.0133575 0.0480372
+ 9.78e+10Hz 0.0133761 0.0480828
+ 9.79e+10Hz 0.0133948 0.0481283
+ 9.8e+10Hz 0.0134134 0.0481739
+ 9.81e+10Hz 0.013432 0.0482195
+ 9.82e+10Hz 0.0134507 0.048265
+ 9.83e+10Hz 0.0134693 0.0483106
+ 9.84e+10Hz 0.013488 0.0483561
+ 9.85e+10Hz 0.0135067 0.0484016
+ 9.86e+10Hz 0.0135255 0.0484471
+ 9.87e+10Hz 0.0135442 0.0484926
+ 9.88e+10Hz 0.013563 0.0485381
+ 9.89e+10Hz 0.0135817 0.0485836
+ 9.9e+10Hz 0.0136005 0.0486291
+ 9.91e+10Hz 0.0136193 0.0486746
+ 9.92e+10Hz 0.0136381 0.04872
+ 9.93e+10Hz 0.0136569 0.0487655
+ 9.94e+10Hz 0.0136758 0.0488109
+ 9.95e+10Hz 0.0136946 0.0488564
+ 9.96e+10Hz 0.0137135 0.0489018
+ 9.97e+10Hz 0.0137324 0.0489472
+ 9.98e+10Hz 0.0137513 0.0489926
+ 9.99e+10Hz 0.0137702 0.049038
+ 1e+11Hz 0.0137892 0.0490834
+ 1.001e+11Hz 0.0138081 0.0491288
+ 1.002e+11Hz 0.0138271 0.0491741
+ 1.003e+11Hz 0.0138461 0.0492195
+ 1.004e+11Hz 0.0138651 0.0492649
+ 1.005e+11Hz 0.0138841 0.0493102
+ 1.006e+11Hz 0.0139031 0.0493555
+ 1.007e+11Hz 0.0139221 0.0494009
+ 1.008e+11Hz 0.0139412 0.0494462
+ 1.009e+11Hz 0.0139603 0.0494915
+ 1.01e+11Hz 0.0139794 0.0495368
+ 1.011e+11Hz 0.0139985 0.0495821
+ 1.012e+11Hz 0.0140176 0.0496274
+ 1.013e+11Hz 0.0140367 0.0496726
+ 1.014e+11Hz 0.0140558 0.0497179
+ 1.015e+11Hz 0.014075 0.0497632
+ 1.016e+11Hz 0.0140942 0.0498084
+ 1.017e+11Hz 0.0141134 0.0498536
+ 1.018e+11Hz 0.0141326 0.0498989
+ 1.019e+11Hz 0.0141518 0.0499441
+ 1.02e+11Hz 0.014171 0.0499893
+ 1.021e+11Hz 0.0141903 0.0500345
+ 1.022e+11Hz 0.0142095 0.0500797
+ 1.023e+11Hz 0.0142288 0.0501249
+ 1.024e+11Hz 0.0142481 0.0501701
+ 1.025e+11Hz 0.0142674 0.0502152
+ 1.026e+11Hz 0.0142868 0.0502604
+ 1.027e+11Hz 0.0143061 0.0503056
+ 1.028e+11Hz 0.0143254 0.0503507
+ 1.029e+11Hz 0.0143448 0.0503958
+ 1.03e+11Hz 0.0143642 0.050441
+ 1.031e+11Hz 0.0143836 0.0504861
+ 1.032e+11Hz 0.014403 0.0505312
+ 1.033e+11Hz 0.0144224 0.0505763
+ 1.034e+11Hz 0.0144419 0.0506214
+ 1.035e+11Hz 0.0144613 0.0506665
+ 1.036e+11Hz 0.0144808 0.0507116
+ 1.037e+11Hz 0.0145003 0.0507566
+ 1.038e+11Hz 0.0145198 0.0508017
+ 1.039e+11Hz 0.0145393 0.0508468
+ 1.04e+11Hz 0.0145588 0.0508918
+ 1.041e+11Hz 0.0145784 0.0509368
+ 1.042e+11Hz 0.0145979 0.0509819
+ 1.043e+11Hz 0.0146175 0.0510269
+ 1.044e+11Hz 0.0146371 0.0510719
+ 1.045e+11Hz 0.0146567 0.0511169
+ 1.046e+11Hz 0.0146763 0.0511619
+ 1.047e+11Hz 0.0146959 0.0512069
+ 1.048e+11Hz 0.0147156 0.0512519
+ 1.049e+11Hz 0.0147352 0.0512969
+ 1.05e+11Hz 0.0147549 0.0513418
+ 1.051e+11Hz 0.0147746 0.0513868
+ 1.052e+11Hz 0.0147943 0.0514317
+ 1.053e+11Hz 0.014814 0.0514767
+ 1.054e+11Hz 0.0148337 0.0515216
+ 1.055e+11Hz 0.0148535 0.0515666
+ 1.056e+11Hz 0.0148733 0.0516115
+ 1.057e+11Hz 0.014893 0.0516564
+ 1.058e+11Hz 0.0149128 0.0517013
+ 1.059e+11Hz 0.0149326 0.0517462
+ 1.06e+11Hz 0.0149525 0.0517911
+ 1.061e+11Hz 0.0149723 0.051836
+ 1.062e+11Hz 0.0149921 0.0518808
+ 1.063e+11Hz 0.015012 0.0519257
+ 1.064e+11Hz 0.0150319 0.0519706
+ 1.065e+11Hz 0.0150518 0.0520154
+ 1.066e+11Hz 0.0150717 0.0520603
+ 1.067e+11Hz 0.0150916 0.0521051
+ 1.068e+11Hz 0.0151116 0.05215
+ 1.069e+11Hz 0.0151315 0.0521948
+ 1.07e+11Hz 0.0151515 0.0522396
+ 1.071e+11Hz 0.0151715 0.0522844
+ 1.072e+11Hz 0.0151915 0.0523292
+ 1.073e+11Hz 0.0152115 0.052374
+ 1.074e+11Hz 0.0152315 0.0524188
+ 1.075e+11Hz 0.0152516 0.0524636
+ 1.076e+11Hz 0.0152716 0.0525083
+ 1.077e+11Hz 0.0152917 0.0525531
+ 1.078e+11Hz 0.0153118 0.0525979
+ 1.079e+11Hz 0.0153319 0.0526426
+ 1.08e+11Hz 0.015352 0.0526874
+ 1.081e+11Hz 0.0153722 0.0527321
+ 1.082e+11Hz 0.0153923 0.0527768
+ 1.083e+11Hz 0.0154125 0.0528215
+ 1.084e+11Hz 0.0154327 0.0528663
+ 1.085e+11Hz 0.0154529 0.052911
+ 1.086e+11Hz 0.0154731 0.0529557
+ 1.087e+11Hz 0.0154933 0.0530004
+ 1.088e+11Hz 0.0155135 0.0530451
+ 1.089e+11Hz 0.0155338 0.0530897
+ 1.09e+11Hz 0.0155541 0.0531344
+ 1.091e+11Hz 0.0155744 0.0531791
+ 1.092e+11Hz 0.0155947 0.0532237
+ 1.093e+11Hz 0.015615 0.0532684
+ 1.094e+11Hz 0.0156353 0.053313
+ 1.095e+11Hz 0.0156557 0.0533576
+ 1.096e+11Hz 0.015676 0.0534023
+ 1.097e+11Hz 0.0156964 0.0534469
+ 1.098e+11Hz 0.0157168 0.0534915
+ 1.099e+11Hz 0.0157372 0.0535361
+ 1.1e+11Hz 0.0157577 0.0535807
+ 1.101e+11Hz 0.0157781 0.0536253
+ 1.102e+11Hz 0.0157986 0.0536699
+ 1.103e+11Hz 0.015819 0.0537145
+ 1.104e+11Hz 0.0158395 0.053759
+ 1.105e+11Hz 0.01586 0.0538036
+ 1.106e+11Hz 0.0158806 0.0538482
+ 1.107e+11Hz 0.0159011 0.0538927
+ 1.108e+11Hz 0.0159217 0.0539372
+ 1.109e+11Hz 0.0159422 0.0539818
+ 1.11e+11Hz 0.0159628 0.0540263
+ 1.111e+11Hz 0.0159834 0.0540708
+ 1.112e+11Hz 0.016004 0.0541153
+ 1.113e+11Hz 0.0160247 0.0541598
+ 1.114e+11Hz 0.0160453 0.0542043
+ 1.115e+11Hz 0.016066 0.0542488
+ 1.116e+11Hz 0.0160867 0.0542933
+ 1.117e+11Hz 0.0161074 0.0543378
+ 1.118e+11Hz 0.0161281 0.0543823
+ 1.119e+11Hz 0.0161488 0.0544267
+ 1.12e+11Hz 0.0161696 0.0544712
+ 1.121e+11Hz 0.0161903 0.0545156
+ 1.122e+11Hz 0.0162111 0.05456
+ 1.123e+11Hz 0.0162319 0.0546045
+ 1.124e+11Hz 0.0162527 0.0546489
+ 1.125e+11Hz 0.0162736 0.0546933
+ 1.126e+11Hz 0.0162944 0.0547377
+ 1.127e+11Hz 0.0163153 0.0547821
+ 1.128e+11Hz 0.0163362 0.0548265
+ 1.129e+11Hz 0.0163571 0.0548709
+ 1.13e+11Hz 0.016378 0.0549153
+ 1.131e+11Hz 0.0163989 0.0549596
+ 1.132e+11Hz 0.0164199 0.055004
+ 1.133e+11Hz 0.0164408 0.0550483
+ 1.134e+11Hz 0.0164618 0.0550927
+ 1.135e+11Hz 0.0164828 0.055137
+ 1.136e+11Hz 0.0165038 0.0551813
+ 1.137e+11Hz 0.0165249 0.0552257
+ 1.138e+11Hz 0.0165459 0.05527
+ 1.139e+11Hz 0.016567 0.0553143
+ 1.14e+11Hz 0.016588 0.0553586
+ 1.141e+11Hz 0.0166091 0.0554029
+ 1.142e+11Hz 0.0166303 0.0554471
+ 1.143e+11Hz 0.0166514 0.0554914
+ 1.144e+11Hz 0.0166725 0.0555357
+ 1.145e+11Hz 0.0166937 0.0555799
+ 1.146e+11Hz 0.0167149 0.0556242
+ 1.147e+11Hz 0.0167361 0.0556684
+ 1.148e+11Hz 0.0167573 0.0557126
+ 1.149e+11Hz 0.0167785 0.0557569
+ 1.15e+11Hz 0.0167998 0.0558011
+ 1.151e+11Hz 0.0168211 0.0558453
+ 1.152e+11Hz 0.0168423 0.0558895
+ 1.153e+11Hz 0.0168637 0.0559337
+ 1.154e+11Hz 0.016885 0.0559778
+ 1.155e+11Hz 0.0169063 0.056022
+ 1.156e+11Hz 0.0169277 0.0560661
+ 1.157e+11Hz 0.016949 0.0561103
+ 1.158e+11Hz 0.0169704 0.0561544
+ 1.159e+11Hz 0.0169918 0.0561986
+ 1.16e+11Hz 0.0170132 0.0562427
+ 1.161e+11Hz 0.0170347 0.0562868
+ 1.162e+11Hz 0.0170561 0.0563309
+ 1.163e+11Hz 0.0170776 0.056375
+ 1.164e+11Hz 0.0170991 0.0564191
+ 1.165e+11Hz 0.0171206 0.0564631
+ 1.166e+11Hz 0.0171421 0.0565072
+ 1.167e+11Hz 0.0171637 0.0565513
+ 1.168e+11Hz 0.0171852 0.0565953
+ 1.169e+11Hz 0.0172068 0.0566394
+ 1.17e+11Hz 0.0172284 0.0566834
+ 1.171e+11Hz 0.01725 0.0567274
+ 1.172e+11Hz 0.0172716 0.0567714
+ 1.173e+11Hz 0.0172933 0.0568154
+ 1.174e+11Hz 0.017315 0.0568594
+ 1.175e+11Hz 0.0173366 0.0569034
+ 1.176e+11Hz 0.0173583 0.0569473
+ 1.177e+11Hz 0.0173801 0.0569913
+ 1.178e+11Hz 0.0174018 0.0570352
+ 1.179e+11Hz 0.0174235 0.0570792
+ 1.18e+11Hz 0.0174453 0.0571231
+ 1.181e+11Hz 0.0174671 0.057167
+ 1.182e+11Hz 0.0174889 0.0572109
+ 1.183e+11Hz 0.0175107 0.0572548
+ 1.184e+11Hz 0.0175325 0.0572987
+ 1.185e+11Hz 0.0175544 0.0573426
+ 1.186e+11Hz 0.0175763 0.0573864
+ 1.187e+11Hz 0.0175981 0.0574303
+ 1.188e+11Hz 0.01762 0.0574741
+ 1.189e+11Hz 0.0176419 0.057518
+ 1.19e+11Hz 0.0176639 0.0575618
+ 1.191e+11Hz 0.0176858 0.0576056
+ 1.192e+11Hz 0.0177078 0.0576494
+ 1.193e+11Hz 0.0177298 0.0576932
+ 1.194e+11Hz 0.0177518 0.057737
+ 1.195e+11Hz 0.0177738 0.0577807
+ 1.196e+11Hz 0.0177959 0.0578245
+ 1.197e+11Hz 0.0178179 0.0578682
+ 1.198e+11Hz 0.01784 0.0579119
+ 1.199e+11Hz 0.0178621 0.0579557
+ 1.2e+11Hz 0.0178842 0.0579994
+ 1.201e+11Hz 0.0179063 0.0580431
+ 1.202e+11Hz 0.0179284 0.0580867
+ 1.203e+11Hz 0.0179506 0.0581304
+ 1.204e+11Hz 0.0179727 0.0581741
+ 1.205e+11Hz 0.0179949 0.0582177
+ 1.206e+11Hz 0.0180171 0.0582614
+ 1.207e+11Hz 0.0180394 0.058305
+ 1.208e+11Hz 0.0180616 0.0583486
+ 1.209e+11Hz 0.0180838 0.0583922
+ 1.21e+11Hz 0.0181061 0.0584358
+ 1.211e+11Hz 0.0181284 0.0584794
+ 1.212e+11Hz 0.0181507 0.0585229
+ 1.213e+11Hz 0.018173 0.0585665
+ 1.214e+11Hz 0.0181954 0.05861
+ 1.215e+11Hz 0.0182177 0.0586536
+ 1.216e+11Hz 0.0182401 0.0586971
+ 1.217e+11Hz 0.0182625 0.0587406
+ 1.218e+11Hz 0.0182848 0.0587841
+ 1.219e+11Hz 0.0183073 0.0588276
+ 1.22e+11Hz 0.0183297 0.058871
+ 1.221e+11Hz 0.0183521 0.0589145
+ 1.222e+11Hz 0.0183746 0.0589579
+ 1.223e+11Hz 0.0183971 0.0590014
+ 1.224e+11Hz 0.0184196 0.0590448
+ 1.225e+11Hz 0.0184421 0.0590882
+ 1.226e+11Hz 0.0184646 0.0591316
+ 1.227e+11Hz 0.0184871 0.0591749
+ 1.228e+11Hz 0.0185097 0.0592183
+ 1.229e+11Hz 0.0185323 0.0592617
+ 1.23e+11Hz 0.0185549 0.059305
+ 1.231e+11Hz 0.0185774 0.0593483
+ 1.232e+11Hz 0.0186001 0.0593916
+ 1.233e+11Hz 0.0186227 0.0594349
+ 1.234e+11Hz 0.0186454 0.0594782
+ 1.235e+11Hz 0.018668 0.0595215
+ 1.236e+11Hz 0.0186907 0.0595648
+ 1.237e+11Hz 0.0187134 0.059608
+ 1.238e+11Hz 0.0187361 0.0596512
+ 1.239e+11Hz 0.0187588 0.0596945
+ 1.24e+11Hz 0.0187815 0.0597377
+ 1.241e+11Hz 0.0188043 0.0597809
+ 1.242e+11Hz 0.0188271 0.059824
+ 1.243e+11Hz 0.0188498 0.0598672
+ 1.244e+11Hz 0.0188726 0.0599104
+ 1.245e+11Hz 0.0188954 0.0599535
+ 1.246e+11Hz 0.0189183 0.0599966
+ 1.247e+11Hz 0.0189411 0.0600398
+ 1.248e+11Hz 0.0189639 0.0600829
+ 1.249e+11Hz 0.0189868 0.0601259
+ 1.25e+11Hz 0.0190097 0.060169
+ 1.251e+11Hz 0.0190326 0.0602121
+ 1.252e+11Hz 0.0190555 0.0602551
+ 1.253e+11Hz 0.0190784 0.0602982
+ 1.254e+11Hz 0.0191013 0.0603412
+ 1.255e+11Hz 0.0191243 0.0603842
+ 1.256e+11Hz 0.0191473 0.0604272
+ 1.257e+11Hz 0.0191702 0.0604702
+ 1.258e+11Hz 0.0191932 0.0605131
+ 1.259e+11Hz 0.0192162 0.0605561
+ 1.26e+11Hz 0.0192392 0.060599
+ 1.261e+11Hz 0.0192623 0.060642
+ 1.262e+11Hz 0.0192853 0.0606849
+ 1.263e+11Hz 0.0193084 0.0607278
+ 1.264e+11Hz 0.0193314 0.0607707
+ 1.265e+11Hz 0.0193545 0.0608135
+ 1.266e+11Hz 0.0193776 0.0608564
+ 1.267e+11Hz 0.0194007 0.0608992
+ 1.268e+11Hz 0.0194238 0.0609421
+ 1.269e+11Hz 0.019447 0.0609849
+ 1.27e+11Hz 0.0194701 0.0610277
+ 1.271e+11Hz 0.0194933 0.0610705
+ 1.272e+11Hz 0.0195165 0.0611133
+ 1.273e+11Hz 0.0195397 0.061156
+ 1.274e+11Hz 0.0195629 0.0611988
+ 1.275e+11Hz 0.0195861 0.0612415
+ 1.276e+11Hz 0.0196093 0.0612842
+ 1.277e+11Hz 0.0196325 0.0613269
+ 1.278e+11Hz 0.0196558 0.0613696
+ 1.279e+11Hz 0.019679 0.0614123
+ 1.28e+11Hz 0.0197023 0.061455
+ 1.281e+11Hz 0.0197256 0.0614977
+ 1.282e+11Hz 0.0197489 0.0615403
+ 1.283e+11Hz 0.0197722 0.0615829
+ 1.284e+11Hz 0.0197955 0.0616256
+ 1.285e+11Hz 0.0198189 0.0616682
+ 1.286e+11Hz 0.0198422 0.0617108
+ 1.287e+11Hz 0.0198656 0.0617533
+ 1.288e+11Hz 0.0198889 0.0617959
+ 1.289e+11Hz 0.0199123 0.0618385
+ 1.29e+11Hz 0.0199357 0.061881
+ 1.291e+11Hz 0.0199591 0.0619235
+ 1.292e+11Hz 0.0199825 0.0619661
+ 1.293e+11Hz 0.020006 0.0620086
+ 1.294e+11Hz 0.0200294 0.0620511
+ 1.295e+11Hz 0.0200529 0.0620935
+ 1.296e+11Hz 0.0200763 0.062136
+ 1.297e+11Hz 0.0200998 0.0621785
+ 1.298e+11Hz 0.0201233 0.0622209
+ 1.299e+11Hz 0.0201468 0.0622633
+ 1.3e+11Hz 0.0201703 0.0623057
+ 1.301e+11Hz 0.0201938 0.0623481
+ 1.302e+11Hz 0.0202173 0.0623905
+ 1.303e+11Hz 0.0202409 0.0624329
+ 1.304e+11Hz 0.0202644 0.0624753
+ 1.305e+11Hz 0.020288 0.0625176
+ 1.306e+11Hz 0.0203116 0.06256
+ 1.307e+11Hz 0.0203352 0.0626023
+ 1.308e+11Hz 0.0203588 0.0626446
+ 1.309e+11Hz 0.0203824 0.0626869
+ 1.31e+11Hz 0.020406 0.0627292
+ 1.311e+11Hz 0.0204296 0.0627715
+ 1.312e+11Hz 0.0204533 0.0628138
+ 1.313e+11Hz 0.0204769 0.062856
+ 1.314e+11Hz 0.0205006 0.0628983
+ 1.315e+11Hz 0.0205243 0.0629405
+ 1.316e+11Hz 0.0205479 0.0629828
+ 1.317e+11Hz 0.0205717 0.063025
+ 1.318e+11Hz 0.0205954 0.0630672
+ 1.319e+11Hz 0.0206191 0.0631094
+ 1.32e+11Hz 0.0206428 0.0631515
+ 1.321e+11Hz 0.0206666 0.0631937
+ 1.322e+11Hz 0.0206903 0.0632359
+ 1.323e+11Hz 0.0207141 0.063278
+ 1.324e+11Hz 0.0207379 0.0633202
+ 1.325e+11Hz 0.0207616 0.0633623
+ 1.326e+11Hz 0.0207855 0.0634044
+ 1.327e+11Hz 0.0208093 0.0634465
+ 1.328e+11Hz 0.0208331 0.0634886
+ 1.329e+11Hz 0.0208569 0.0635307
+ 1.33e+11Hz 0.0208808 0.0635727
+ 1.331e+11Hz 0.0209046 0.0636148
+ 1.332e+11Hz 0.0209285 0.0636568
+ 1.333e+11Hz 0.0209524 0.0636989
+ 1.334e+11Hz 0.0209762 0.0637409
+ 1.335e+11Hz 0.0210001 0.0637829
+ 1.336e+11Hz 0.021024 0.0638249
+ 1.337e+11Hz 0.021048 0.0638669
+ 1.338e+11Hz 0.0210719 0.0639089
+ 1.339e+11Hz 0.0210958 0.0639509
+ 1.34e+11Hz 0.0211198 0.0639929
+ 1.341e+11Hz 0.0211438 0.0640348
+ 1.342e+11Hz 0.0211678 0.0640768
+ 1.343e+11Hz 0.0211917 0.0641187
+ 1.344e+11Hz 0.0212157 0.0641606
+ 1.345e+11Hz 0.0212398 0.0642026
+ 1.346e+11Hz 0.0212638 0.0642445
+ 1.347e+11Hz 0.0212878 0.0642864
+ 1.348e+11Hz 0.0213119 0.0643283
+ 1.349e+11Hz 0.0213359 0.0643702
+ 1.35e+11Hz 0.02136 0.064412
+ 1.351e+11Hz 0.0213841 0.0644539
+ 1.352e+11Hz 0.0214082 0.0644958
+ 1.353e+11Hz 0.0214323 0.0645376
+ 1.354e+11Hz 0.0214564 0.0645794
+ 1.355e+11Hz 0.0214806 0.0646213
+ 1.356e+11Hz 0.0215047 0.0646631
+ 1.357e+11Hz 0.0215289 0.0647049
+ 1.358e+11Hz 0.021553 0.0647467
+ 1.359e+11Hz 0.0215772 0.0647885
+ 1.36e+11Hz 0.0216014 0.0648303
+ 1.361e+11Hz 0.0216256 0.064872
+ 1.362e+11Hz 0.0216499 0.0649138
+ 1.363e+11Hz 0.0216741 0.0649556
+ 1.364e+11Hz 0.0216983 0.0649973
+ 1.365e+11Hz 0.0217226 0.065039
+ 1.366e+11Hz 0.0217469 0.0650808
+ 1.367e+11Hz 0.0217712 0.0651225
+ 1.368e+11Hz 0.0217955 0.0651642
+ 1.369e+11Hz 0.0218198 0.0652059
+ 1.37e+11Hz 0.0218441 0.0652476
+ 1.371e+11Hz 0.0218685 0.0652893
+ 1.372e+11Hz 0.0218928 0.065331
+ 1.373e+11Hz 0.0219172 0.0653727
+ 1.374e+11Hz 0.0219416 0.0654143
+ 1.375e+11Hz 0.021966 0.065456
+ 1.376e+11Hz 0.0219904 0.0654976
+ 1.377e+11Hz 0.0220148 0.0655393
+ 1.378e+11Hz 0.0220392 0.0655809
+ 1.379e+11Hz 0.0220637 0.0656225
+ 1.38e+11Hz 0.0220882 0.0656641
+ 1.381e+11Hz 0.0221126 0.0657057
+ 1.382e+11Hz 0.0221371 0.0657473
+ 1.383e+11Hz 0.0221616 0.0657889
+ 1.384e+11Hz 0.0221862 0.0658305
+ 1.385e+11Hz 0.0222107 0.0658721
+ 1.386e+11Hz 0.0222353 0.0659137
+ 1.387e+11Hz 0.0222598 0.0659552
+ 1.388e+11Hz 0.0222844 0.0659968
+ 1.389e+11Hz 0.022309 0.0660383
+ 1.39e+11Hz 0.0223337 0.0660798
+ 1.391e+11Hz 0.0223583 0.0661214
+ 1.392e+11Hz 0.0223829 0.0661629
+ 1.393e+11Hz 0.0224076 0.0662044
+ 1.394e+11Hz 0.0224323 0.0662459
+ 1.395e+11Hz 0.022457 0.0662874
+ 1.396e+11Hz 0.0224817 0.0663289
+ 1.397e+11Hz 0.0225064 0.0663704
+ 1.398e+11Hz 0.0225312 0.0664118
+ 1.399e+11Hz 0.0225559 0.0664533
+ 1.4e+11Hz 0.0225807 0.0664947
+ 1.401e+11Hz 0.0226055 0.0665362
+ 1.402e+11Hz 0.0226303 0.0665776
+ 1.403e+11Hz 0.0226552 0.066619
+ 1.404e+11Hz 0.02268 0.0666605
+ 1.405e+11Hz 0.0227049 0.0667019
+ 1.406e+11Hz 0.0227298 0.0667433
+ 1.407e+11Hz 0.0227547 0.0667847
+ 1.408e+11Hz 0.0227796 0.0668261
+ 1.409e+11Hz 0.0228045 0.0668674
+ 1.41e+11Hz 0.0228295 0.0669088
+ 1.411e+11Hz 0.0228545 0.0669502
+ 1.412e+11Hz 0.0228795 0.0669915
+ 1.413e+11Hz 0.0229045 0.0670329
+ 1.414e+11Hz 0.0229295 0.0670742
+ 1.415e+11Hz 0.0229546 0.0671155
+ 1.416e+11Hz 0.0229796 0.0671569
+ 1.417e+11Hz 0.0230047 0.0671982
+ 1.418e+11Hz 0.0230298 0.0672395
+ 1.419e+11Hz 0.0230549 0.0672808
+ 1.42e+11Hz 0.0230801 0.067322
+ 1.421e+11Hz 0.0231053 0.0673633
+ 1.422e+11Hz 0.0231304 0.0674046
+ 1.423e+11Hz 0.0231556 0.0674458
+ 1.424e+11Hz 0.0231808 0.0674871
+ 1.425e+11Hz 0.0232061 0.0675283
+ 1.426e+11Hz 0.0232314 0.0675695
+ 1.427e+11Hz 0.0232566 0.0676107
+ 1.428e+11Hz 0.0232819 0.0676519
+ 1.429e+11Hz 0.0233073 0.0676931
+ 1.43e+11Hz 0.0233326 0.0677343
+ 1.431e+11Hz 0.023358 0.0677755
+ 1.432e+11Hz 0.0233834 0.0678166
+ 1.433e+11Hz 0.0234088 0.0678578
+ 1.434e+11Hz 0.0234342 0.0678989
+ 1.435e+11Hz 0.0234596 0.0679401
+ 1.436e+11Hz 0.0234851 0.0679812
+ 1.437e+11Hz 0.0235106 0.0680223
+ 1.438e+11Hz 0.0235361 0.0680634
+ 1.439e+11Hz 0.0235616 0.0681045
+ 1.44e+11Hz 0.0235872 0.0681455
+ 1.441e+11Hz 0.0236128 0.0681866
+ 1.442e+11Hz 0.0236384 0.0682277
+ 1.443e+11Hz 0.023664 0.0682687
+ 1.444e+11Hz 0.0236896 0.0683097
+ 1.445e+11Hz 0.0237153 0.0683508
+ 1.446e+11Hz 0.023741 0.0683918
+ 1.447e+11Hz 0.0237667 0.0684328
+ 1.448e+11Hz 0.0237924 0.0684737
+ 1.449e+11Hz 0.0238181 0.0685147
+ 1.45e+11Hz 0.0238439 0.0685556
+ 1.451e+11Hz 0.0238697 0.0685966
+ 1.452e+11Hz 0.0238955 0.0686375
+ 1.453e+11Hz 0.0239214 0.0686784
+ 1.454e+11Hz 0.0239472 0.0687193
+ 1.455e+11Hz 0.0239731 0.0687602
+ 1.456e+11Hz 0.023999 0.0688011
+ 1.457e+11Hz 0.0240249 0.068842
+ 1.458e+11Hz 0.0240509 0.0688828
+ 1.459e+11Hz 0.0240769 0.0689236
+ 1.46e+11Hz 0.0241028 0.0689645
+ 1.461e+11Hz 0.0241289 0.0690053
+ 1.462e+11Hz 0.0241549 0.0690461
+ 1.463e+11Hz 0.024181 0.0690868
+ 1.464e+11Hz 0.0242071 0.0691276
+ 1.465e+11Hz 0.0242332 0.0691683
+ 1.466e+11Hz 0.0242593 0.0692091
+ 1.467e+11Hz 0.0242855 0.0692498
+ 1.468e+11Hz 0.0243116 0.0692905
+ 1.469e+11Hz 0.0243378 0.0693312
+ 1.47e+11Hz 0.0243641 0.0693718
+ 1.471e+11Hz 0.0243903 0.0694125
+ 1.472e+11Hz 0.0244166 0.0694531
+ 1.473e+11Hz 0.0244428 0.0694937
+ 1.474e+11Hz 0.0244692 0.0695343
+ 1.475e+11Hz 0.0244955 0.0695749
+ 1.476e+11Hz 0.0245219 0.0696155
+ 1.477e+11Hz 0.0245482 0.069656
+ 1.478e+11Hz 0.0245746 0.0696966
+ 1.479e+11Hz 0.0246011 0.0697371
+ 1.48e+11Hz 0.0246275 0.0697776
+ 1.481e+11Hz 0.024654 0.0698181
+ 1.482e+11Hz 0.0246805 0.0698586
+ 1.483e+11Hz 0.024707 0.069899
+ 1.484e+11Hz 0.0247335 0.0699394
+ 1.485e+11Hz 0.0247601 0.0699798
+ 1.486e+11Hz 0.0247867 0.0700202
+ 1.487e+11Hz 0.0248133 0.0700606
+ 1.488e+11Hz 0.0248399 0.0701009
+ 1.489e+11Hz 0.0248666 0.0701413
+ 1.49e+11Hz 0.0248932 0.0701816
+ 1.491e+11Hz 0.0249199 0.0702219
+ 1.492e+11Hz 0.0249467 0.0702622
+ 1.493e+11Hz 0.0249734 0.0703024
+ 1.494e+11Hz 0.0250001 0.0703427
+ 1.495e+11Hz 0.0250269 0.0703829
+ 1.496e+11Hz 0.0250537 0.0704231
+ 1.497e+11Hz 0.0250806 0.0704633
+ 1.498e+11Hz 0.0251074 0.0705034
+ 1.499e+11Hz 0.0251343 0.0705436
+ 1.5e+11Hz 0.0251612 0.0705837
+ ]

.ENDS
.SUBCKT Sub_SPfile_X7 1 2 3
R1N 1 10 -50
R1P 10 11 100
R2N 2 20 -50
R2P 20 21 100

A11 %vd(10 3) %vd(11, 12) xfer1
.model xfer1 xfer R_I=true table=[
+ 0Hz 0.00397698 0
+ 1e+08Hz 0.00397718 -3.28303e-05
+ 2e+08Hz 0.00397776 -6.56684e-05
+ 3e+08Hz 0.00397872 -9.8522e-05
+ 4e+08Hz 0.00398007 -0.000131399
+ 5e+08Hz 0.00398181 -0.000164307
+ 6e+08Hz 0.00398393 -0.000197254
+ 7e+08Hz 0.00398644 -0.000230247
+ 8e+08Hz 0.00398932 -0.000263294
+ 9e+08Hz 0.00399259 -0.000296403
+ 1e+09Hz 0.00399623 -0.000329581
+ 1.1e+09Hz 0.00400026 -0.000362837
+ 1.2e+09Hz 0.00400466 -0.000396176
+ 1.3e+09Hz 0.00400943 -0.000429608
+ 1.4e+09Hz 0.00401458 -0.000463139
+ 1.5e+09Hz 0.00402009 -0.000496777
+ 1.6e+09Hz 0.00402597 -0.000530528
+ 1.7e+09Hz 0.00403221 -0.000564401
+ 1.8e+09Hz 0.00403882 -0.000598402
+ 1.9e+09Hz 0.00404578 -0.000632539
+ 2e+09Hz 0.00405309 -0.000666817
+ 2.1e+09Hz 0.00406076 -0.000701246
+ 2.2e+09Hz 0.00406878 -0.00073583
+ 2.3e+09Hz 0.00407714 -0.000770577
+ 2.4e+09Hz 0.00408584 -0.000805493
+ 2.5e+09Hz 0.00409487 -0.000840585
+ 2.6e+09Hz 0.00410424 -0.00087586
+ 2.7e+09Hz 0.00411394 -0.000911324
+ 2.8e+09Hz 0.00412396 -0.000946982
+ 2.9e+09Hz 0.00413429 -0.000982842
+ 3e+09Hz 0.00414495 -0.00101891
+ 3.1e+09Hz 0.00415591 -0.00105519
+ 3.2e+09Hz 0.00416718 -0.00109169
+ 3.3e+09Hz 0.00417874 -0.00112841
+ 3.4e+09Hz 0.0041906 -0.00116536
+ 3.5e+09Hz 0.00420275 -0.00120255
+ 3.6e+09Hz 0.00421519 -0.00123997
+ 3.7e+09Hz 0.0042279 -0.00127765
+ 3.8e+09Hz 0.00424088 -0.00131557
+ 3.9e+09Hz 0.00425414 -0.00135375
+ 4e+09Hz 0.00426765 -0.00139219
+ 4.1e+09Hz 0.00428142 -0.00143089
+ 4.2e+09Hz 0.00429544 -0.00146986
+ 4.3e+09Hz 0.0043097 -0.00150911
+ 4.4e+09Hz 0.0043242 -0.00154863
+ 4.5e+09Hz 0.00433893 -0.00158843
+ 4.6e+09Hz 0.00435388 -0.00162852
+ 4.7e+09Hz 0.00436906 -0.00166889
+ 4.8e+09Hz 0.00438444 -0.00170956
+ 4.9e+09Hz 0.00440003 -0.00175052
+ 5e+09Hz 0.00441582 -0.00179179
+ 5.1e+09Hz 0.00443181 -0.00183335
+ 5.2e+09Hz 0.00444798 -0.00187522
+ 5.3e+09Hz 0.00446433 -0.00191739
+ 5.4e+09Hz 0.00448085 -0.00195987
+ 5.5e+09Hz 0.00449754 -0.00200267
+ 5.6e+09Hz 0.00451439 -0.00204578
+ 5.7e+09Hz 0.00453139 -0.00208921
+ 5.8e+09Hz 0.00454853 -0.00213295
+ 5.9e+09Hz 0.00456582 -0.00217702
+ 6e+09Hz 0.00458324 -0.0022214
+ 6.1e+09Hz 0.00460078 -0.00226611
+ 6.2e+09Hz 0.00461844 -0.00231115
+ 6.3e+09Hz 0.00463622 -0.0023565
+ 6.4e+09Hz 0.00465409 -0.00240219
+ 6.5e+09Hz 0.00467207 -0.0024482
+ 6.6e+09Hz 0.00469014 -0.00249454
+ 6.7e+09Hz 0.00470829 -0.00254121
+ 6.8e+09Hz 0.00472652 -0.00258821
+ 6.9e+09Hz 0.00474483 -0.00263553
+ 7e+09Hz 0.00476319 -0.00268319
+ 7.1e+09Hz 0.00478162 -0.00273117
+ 7.2e+09Hz 0.00480009 -0.00277948
+ 7.3e+09Hz 0.00481862 -0.00282812
+ 7.4e+09Hz 0.00483717 -0.00287709
+ 7.5e+09Hz 0.00485576 -0.00292639
+ 7.6e+09Hz 0.00487438 -0.00297601
+ 7.7e+09Hz 0.00489301 -0.00302595
+ 7.8e+09Hz 0.00491166 -0.00307623
+ 7.9e+09Hz 0.00493031 -0.00312682
+ 8e+09Hz 0.00494896 -0.00317774
+ 8.1e+09Hz 0.0049676 -0.00322897
+ 8.2e+09Hz 0.00498623 -0.00328053
+ 8.3e+09Hz 0.00500484 -0.0033324
+ 8.4e+09Hz 0.00502343 -0.00338459
+ 8.5e+09Hz 0.00504199 -0.00343709
+ 8.6e+09Hz 0.00506051 -0.0034899
+ 8.7e+09Hz 0.00507898 -0.00354302
+ 8.8e+09Hz 0.00509741 -0.00359645
+ 8.9e+09Hz 0.00511579 -0.00365018
+ 9e+09Hz 0.0051341 -0.00370421
+ 9.1e+09Hz 0.00515236 -0.00375854
+ 9.2e+09Hz 0.00517054 -0.00381317
+ 9.3e+09Hz 0.00518864 -0.00386809
+ 9.4e+09Hz 0.00520667 -0.00392331
+ 9.5e+09Hz 0.00522461 -0.00397881
+ 9.6e+09Hz 0.00524246 -0.00403459
+ 9.7e+09Hz 0.00526021 -0.00409066
+ 9.8e+09Hz 0.00527787 -0.004147
+ 9.9e+09Hz 0.00529541 -0.00420362
+ 1e+10Hz 0.00531285 -0.00426051
+ 1.01e+10Hz 0.00533018 -0.00431767
+ 1.02e+10Hz 0.00534739 -0.00437509
+ 1.03e+10Hz 0.00536447 -0.00443277
+ 1.04e+10Hz 0.00538143 -0.00449071
+ 1.05e+10Hz 0.00539825 -0.0045489
+ 1.06e+10Hz 0.00541495 -0.00460734
+ 1.07e+10Hz 0.0054315 -0.00466603
+ 1.08e+10Hz 0.00544791 -0.00472496
+ 1.09e+10Hz 0.00546417 -0.00478412
+ 1.1e+10Hz 0.00548029 -0.00484352
+ 1.11e+10Hz 0.00549625 -0.00490315
+ 1.12e+10Hz 0.00551206 -0.004963
+ 1.13e+10Hz 0.0055277 -0.00502307
+ 1.14e+10Hz 0.00554319 -0.00508336
+ 1.15e+10Hz 0.00555851 -0.00514387
+ 1.16e+10Hz 0.00557366 -0.00520458
+ 1.17e+10Hz 0.00558863 -0.00526549
+ 1.18e+10Hz 0.00560344 -0.0053266
+ 1.19e+10Hz 0.00561807 -0.00538791
+ 1.2e+10Hz 0.00563252 -0.00544941
+ 1.21e+10Hz 0.00564679 -0.0055111
+ 1.22e+10Hz 0.00566088 -0.00557297
+ 1.23e+10Hz 0.00567478 -0.00563501
+ 1.24e+10Hz 0.00568849 -0.00569723
+ 1.25e+10Hz 0.00570202 -0.00575961
+ 1.26e+10Hz 0.00571535 -0.00582216
+ 1.27e+10Hz 0.00572849 -0.00588487
+ 1.28e+10Hz 0.00574144 -0.00594773
+ 1.29e+10Hz 0.00575419 -0.00601075
+ 1.3e+10Hz 0.00576675 -0.00607391
+ 1.31e+10Hz 0.00577911 -0.00613721
+ 1.32e+10Hz 0.00579127 -0.00620065
+ 1.33e+10Hz 0.00580323 -0.00626422
+ 1.34e+10Hz 0.00581499 -0.00632792
+ 1.35e+10Hz 0.00582654 -0.00639175
+ 1.36e+10Hz 0.0058379 -0.00645569
+ 1.37e+10Hz 0.00584905 -0.00651975
+ 1.38e+10Hz 0.00586 -0.00658392
+ 1.39e+10Hz 0.00587074 -0.0066482
+ 1.4e+10Hz 0.00588128 -0.00671258
+ 1.41e+10Hz 0.00589162 -0.00677705
+ 1.42e+10Hz 0.00590175 -0.00684162
+ 1.43e+10Hz 0.00591167 -0.00690628
+ 1.44e+10Hz 0.00592139 -0.00697102
+ 1.45e+10Hz 0.00593091 -0.00703585
+ 1.46e+10Hz 0.00594022 -0.00710076
+ 1.47e+10Hz 0.00594933 -0.00716573
+ 1.48e+10Hz 0.00595824 -0.00723078
+ 1.49e+10Hz 0.00596694 -0.00729589
+ 1.5e+10Hz 0.00597544 -0.00736106
+ 1.51e+10Hz 0.00598374 -0.00742629
+ 1.52e+10Hz 0.00599183 -0.00749157
+ 1.53e+10Hz 0.00599973 -0.0075569
+ 1.54e+10Hz 0.00600742 -0.00762228
+ 1.55e+10Hz 0.00601492 -0.0076877
+ 1.56e+10Hz 0.00602222 -0.00775316
+ 1.57e+10Hz 0.00602933 -0.00781865
+ 1.58e+10Hz 0.00603623 -0.00788417
+ 1.59e+10Hz 0.00604295 -0.00794973
+ 1.6e+10Hz 0.00604947 -0.0080153
+ 1.61e+10Hz 0.0060558 -0.0080809
+ 1.62e+10Hz 0.00606193 -0.00814652
+ 1.63e+10Hz 0.00606788 -0.00821215
+ 1.64e+10Hz 0.00607365 -0.00827779
+ 1.65e+10Hz 0.00607922 -0.00834344
+ 1.66e+10Hz 0.00608461 -0.0084091
+ 1.67e+10Hz 0.00608982 -0.00847476
+ 1.68e+10Hz 0.00609485 -0.00854041
+ 1.69e+10Hz 0.0060997 -0.00860607
+ 1.7e+10Hz 0.00610437 -0.00867171
+ 1.71e+10Hz 0.00610887 -0.00873735
+ 1.72e+10Hz 0.00611319 -0.00880298
+ 1.73e+10Hz 0.00611734 -0.00886859
+ 1.74e+10Hz 0.00612133 -0.00893419
+ 1.75e+10Hz 0.00612514 -0.00899976
+ 1.76e+10Hz 0.00612879 -0.00906532
+ 1.77e+10Hz 0.00613227 -0.00913085
+ 1.78e+10Hz 0.00613559 -0.00919635
+ 1.79e+10Hz 0.00613876 -0.00926182
+ 1.8e+10Hz 0.00614176 -0.00932727
+ 1.81e+10Hz 0.00614461 -0.00939268
+ 1.82e+10Hz 0.00614731 -0.00945805
+ 1.83e+10Hz 0.00614986 -0.00952339
+ 1.84e+10Hz 0.00615225 -0.00958869
+ 1.85e+10Hz 0.00615451 -0.00965395
+ 1.86e+10Hz 0.00615661 -0.00971916
+ 1.87e+10Hz 0.00615858 -0.00978433
+ 1.88e+10Hz 0.00616041 -0.00984946
+ 1.89e+10Hz 0.0061621 -0.00991454
+ 1.9e+10Hz 0.00616365 -0.00997957
+ 1.91e+10Hz 0.00616507 -0.0100445
+ 1.92e+10Hz 0.00616637 -0.0101095
+ 1.93e+10Hz 0.00616753 -0.0101744
+ 1.94e+10Hz 0.00616857 -0.0102392
+ 1.95e+10Hz 0.00616949 -0.0103039
+ 1.96e+10Hz 0.00617028 -0.0103686
+ 1.97e+10Hz 0.00617096 -0.0104333
+ 1.98e+10Hz 0.00617152 -0.0104979
+ 1.99e+10Hz 0.00617197 -0.0105624
+ 2e+10Hz 0.00617231 -0.0106269
+ 2.01e+10Hz 0.00617253 -0.0106913
+ 2.02e+10Hz 0.00617266 -0.0107556
+ 2.03e+10Hz 0.00617267 -0.0108199
+ 2.04e+10Hz 0.00617259 -0.0108842
+ 2.05e+10Hz 0.0061724 -0.0109483
+ 2.06e+10Hz 0.00617212 -0.0110124
+ 2.07e+10Hz 0.00617175 -0.0110764
+ 2.08e+10Hz 0.00617128 -0.0111404
+ 2.09e+10Hz 0.00617072 -0.0112043
+ 2.1e+10Hz 0.00617007 -0.0112681
+ 2.11e+10Hz 0.00616934 -0.0113319
+ 2.12e+10Hz 0.00616852 -0.0113956
+ 2.13e+10Hz 0.00616762 -0.0114592
+ 2.14e+10Hz 0.00616665 -0.0115228
+ 2.15e+10Hz 0.00616559 -0.0115863
+ 2.16e+10Hz 0.00616446 -0.0116497
+ 2.17e+10Hz 0.00616326 -0.0117131
+ 2.18e+10Hz 0.00616198 -0.0117764
+ 2.19e+10Hz 0.00616064 -0.0118396
+ 2.2e+10Hz 0.00615923 -0.0119028
+ 2.21e+10Hz 0.00615776 -0.0119659
+ 2.22e+10Hz 0.00615622 -0.0120289
+ 2.23e+10Hz 0.00615463 -0.0120919
+ 2.24e+10Hz 0.00615297 -0.0121548
+ 2.25e+10Hz 0.00615126 -0.0122176
+ 2.26e+10Hz 0.00614949 -0.0122804
+ 2.27e+10Hz 0.00614767 -0.0123431
+ 2.28e+10Hz 0.00614579 -0.0124058
+ 2.29e+10Hz 0.00614387 -0.0124683
+ 2.3e+10Hz 0.0061419 -0.0125309
+ 2.31e+10Hz 0.00613989 -0.0125933
+ 2.32e+10Hz 0.00613783 -0.0126557
+ 2.33e+10Hz 0.00613572 -0.0127181
+ 2.34e+10Hz 0.00613358 -0.0127803
+ 2.35e+10Hz 0.00613139 -0.0128426
+ 2.36e+10Hz 0.00612917 -0.0129047
+ 2.37e+10Hz 0.00612691 -0.0129668
+ 2.38e+10Hz 0.00612461 -0.0130289
+ 2.39e+10Hz 0.00612228 -0.0130909
+ 2.4e+10Hz 0.00611993 -0.0131528
+ 2.41e+10Hz 0.00611753 -0.0132147
+ 2.42e+10Hz 0.00611511 -0.0132765
+ 2.43e+10Hz 0.00611266 -0.0133383
+ 2.44e+10Hz 0.00611018 -0.0134
+ 2.45e+10Hz 0.00610768 -0.0134617
+ 2.46e+10Hz 0.00610516 -0.0135233
+ 2.47e+10Hz 0.0061026 -0.0135849
+ 2.48e+10Hz 0.00610003 -0.0136464
+ 2.49e+10Hz 0.00609744 -0.0137079
+ 2.5e+10Hz 0.00609482 -0.0137694
+ 2.51e+10Hz 0.00609219 -0.0138308
+ 2.52e+10Hz 0.00608953 -0.0138921
+ 2.53e+10Hz 0.00608686 -0.0139534
+ 2.54e+10Hz 0.00608418 -0.0140147
+ 2.55e+10Hz 0.00608147 -0.0140759
+ 2.56e+10Hz 0.00607876 -0.0141371
+ 2.57e+10Hz 0.00607603 -0.0141983
+ 2.58e+10Hz 0.00607328 -0.0142594
+ 2.59e+10Hz 0.00607052 -0.0143205
+ 2.6e+10Hz 0.00606775 -0.0143815
+ 2.61e+10Hz 0.00606497 -0.0144425
+ 2.62e+10Hz 0.00606218 -0.0145035
+ 2.63e+10Hz 0.00605938 -0.0145644
+ 2.64e+10Hz 0.00605657 -0.0146253
+ 2.65e+10Hz 0.00605375 -0.0146862
+ 2.66e+10Hz 0.00605092 -0.0147471
+ 2.67e+10Hz 0.00604808 -0.0148079
+ 2.68e+10Hz 0.00604524 -0.0148687
+ 2.69e+10Hz 0.00604238 -0.0149295
+ 2.7e+10Hz 0.00603952 -0.0149903
+ 2.71e+10Hz 0.00603666 -0.015051
+ 2.72e+10Hz 0.00603378 -0.0151117
+ 2.73e+10Hz 0.0060309 -0.0151724
+ 2.74e+10Hz 0.00602802 -0.0152331
+ 2.75e+10Hz 0.00602513 -0.0152937
+ 2.76e+10Hz 0.00602223 -0.0153544
+ 2.77e+10Hz 0.00601932 -0.015415
+ 2.78e+10Hz 0.00601642 -0.0154756
+ 2.79e+10Hz 0.0060135 -0.0155362
+ 2.8e+10Hz 0.00601058 -0.0155968
+ 2.81e+10Hz 0.00600766 -0.0156574
+ 2.82e+10Hz 0.00600472 -0.0157179
+ 2.83e+10Hz 0.00600179 -0.0157785
+ 2.84e+10Hz 0.00599885 -0.015839
+ 2.85e+10Hz 0.0059959 -0.0158995
+ 2.86e+10Hz 0.00599294 -0.01596
+ 2.87e+10Hz 0.00598998 -0.0160206
+ 2.88e+10Hz 0.00598701 -0.0160811
+ 2.89e+10Hz 0.00598404 -0.0161416
+ 2.9e+10Hz 0.00598106 -0.0162021
+ 2.91e+10Hz 0.00597807 -0.0162626
+ 2.92e+10Hz 0.00597508 -0.0163231
+ 2.93e+10Hz 0.00597208 -0.0163836
+ 2.94e+10Hz 0.00596907 -0.0164441
+ 2.95e+10Hz 0.00596605 -0.0165046
+ 2.96e+10Hz 0.00596303 -0.0165651
+ 2.97e+10Hz 0.00595999 -0.0166256
+ 2.98e+10Hz 0.00595695 -0.0166861
+ 2.99e+10Hz 0.00595389 -0.0167466
+ 3e+10Hz 0.00595083 -0.0168071
+ 3.01e+10Hz 0.00594776 -0.0168676
+ 3.02e+10Hz 0.00594467 -0.0169282
+ 3.03e+10Hz 0.00594158 -0.0169887
+ 3.04e+10Hz 0.00593847 -0.0170492
+ 3.05e+10Hz 0.00593535 -0.0171098
+ 3.06e+10Hz 0.00593221 -0.0171703
+ 3.07e+10Hz 0.00592907 -0.0172309
+ 3.08e+10Hz 0.00592591 -0.0172915
+ 3.09e+10Hz 0.00592273 -0.017352
+ 3.1e+10Hz 0.00591954 -0.0174126
+ 3.11e+10Hz 0.00591634 -0.0174732
+ 3.12e+10Hz 0.00591312 -0.0175338
+ 3.13e+10Hz 0.00590988 -0.0175945
+ 3.14e+10Hz 0.00590663 -0.0176551
+ 3.15e+10Hz 0.00590335 -0.0177157
+ 3.16e+10Hz 0.00590006 -0.0177764
+ 3.17e+10Hz 0.00589675 -0.0178371
+ 3.18e+10Hz 0.00589342 -0.0178978
+ 3.19e+10Hz 0.00589007 -0.0179585
+ 3.2e+10Hz 0.0058867 -0.0180192
+ 3.21e+10Hz 0.00588331 -0.0180799
+ 3.22e+10Hz 0.0058799 -0.0181406
+ 3.23e+10Hz 0.00587646 -0.0182014
+ 3.24e+10Hz 0.005873 -0.0182622
+ 3.25e+10Hz 0.00586952 -0.018323
+ 3.26e+10Hz 0.00586601 -0.0183838
+ 3.27e+10Hz 0.00586248 -0.0184446
+ 3.28e+10Hz 0.00585892 -0.0185054
+ 3.29e+10Hz 0.00585533 -0.0185662
+ 3.3e+10Hz 0.00585172 -0.0186271
+ 3.31e+10Hz 0.00584808 -0.018688
+ 3.32e+10Hz 0.00584441 -0.0187489
+ 3.33e+10Hz 0.00584071 -0.0188098
+ 3.34e+10Hz 0.00583699 -0.0188707
+ 3.35e+10Hz 0.00583323 -0.0189317
+ 3.36e+10Hz 0.00582944 -0.0189926
+ 3.37e+10Hz 0.00582562 -0.0190536
+ 3.38e+10Hz 0.00582177 -0.0191146
+ 3.39e+10Hz 0.00581789 -0.0191756
+ 3.4e+10Hz 0.00581397 -0.0192366
+ 3.41e+10Hz 0.00581002 -0.0192976
+ 3.42e+10Hz 0.00580604 -0.0193587
+ 3.43e+10Hz 0.00580201 -0.0194197
+ 3.44e+10Hz 0.00579796 -0.0194808
+ 3.45e+10Hz 0.00579387 -0.0195419
+ 3.46e+10Hz 0.00578974 -0.019603
+ 3.47e+10Hz 0.00578557 -0.0196641
+ 3.48e+10Hz 0.00578137 -0.0197253
+ 3.49e+10Hz 0.00577713 -0.0197864
+ 3.5e+10Hz 0.00577285 -0.0198476
+ 3.51e+10Hz 0.00576853 -0.0199088
+ 3.52e+10Hz 0.00576417 -0.01997
+ 3.53e+10Hz 0.00575977 -0.0200312
+ 3.54e+10Hz 0.00575533 -0.0200924
+ 3.55e+10Hz 0.00575085 -0.0201536
+ 3.56e+10Hz 0.00574632 -0.0202148
+ 3.57e+10Hz 0.00574176 -0.0202761
+ 3.58e+10Hz 0.00573715 -0.0203373
+ 3.59e+10Hz 0.0057325 -0.0203986
+ 3.6e+10Hz 0.0057278 -0.0204599
+ 3.61e+10Hz 0.00572306 -0.0205211
+ 3.62e+10Hz 0.00571828 -0.0205824
+ 3.63e+10Hz 0.00571345 -0.0206437
+ 3.64e+10Hz 0.00570858 -0.0207051
+ 3.65e+10Hz 0.00570366 -0.0207664
+ 3.66e+10Hz 0.0056987 -0.0208277
+ 3.67e+10Hz 0.00569369 -0.020889
+ 3.68e+10Hz 0.00568863 -0.0209504
+ 3.69e+10Hz 0.00568353 -0.0210117
+ 3.7e+10Hz 0.00567838 -0.0210731
+ 3.71e+10Hz 0.00567318 -0.0211344
+ 3.72e+10Hz 0.00566794 -0.0211958
+ 3.73e+10Hz 0.00566265 -0.0212572
+ 3.74e+10Hz 0.00565731 -0.0213185
+ 3.75e+10Hz 0.00565192 -0.0213799
+ 3.76e+10Hz 0.00564648 -0.0214413
+ 3.77e+10Hz 0.005641 -0.0215026
+ 3.78e+10Hz 0.00563546 -0.021564
+ 3.79e+10Hz 0.00562988 -0.0216254
+ 3.8e+10Hz 0.00562425 -0.0216868
+ 3.81e+10Hz 0.00561856 -0.0217482
+ 3.82e+10Hz 0.00561283 -0.0218095
+ 3.83e+10Hz 0.00560705 -0.0218709
+ 3.84e+10Hz 0.00560122 -0.0219323
+ 3.85e+10Hz 0.00559534 -0.0219936
+ 3.86e+10Hz 0.00558941 -0.022055
+ 3.87e+10Hz 0.00558343 -0.0221164
+ 3.88e+10Hz 0.0055774 -0.0221777
+ 3.89e+10Hz 0.00557132 -0.0222391
+ 3.9e+10Hz 0.00556519 -0.0223004
+ 3.91e+10Hz 0.00555901 -0.0223618
+ 3.92e+10Hz 0.00555278 -0.0224231
+ 3.93e+10Hz 0.0055465 -0.0224844
+ 3.94e+10Hz 0.00554017 -0.0225458
+ 3.95e+10Hz 0.00553379 -0.0226071
+ 3.96e+10Hz 0.00552736 -0.0226684
+ 3.97e+10Hz 0.00552088 -0.0227297
+ 3.98e+10Hz 0.00551435 -0.022791
+ 3.99e+10Hz 0.00550777 -0.0228522
+ 4e+10Hz 0.00550114 -0.0229135
+ 4.01e+10Hz 0.00549446 -0.0229748
+ 4.02e+10Hz 0.00548773 -0.023036
+ 4.03e+10Hz 0.00548096 -0.0230972
+ 4.04e+10Hz 0.00547413 -0.0231585
+ 4.05e+10Hz 0.00546725 -0.0232197
+ 4.06e+10Hz 0.00546033 -0.0232808
+ 4.07e+10Hz 0.00545336 -0.023342
+ 4.08e+10Hz 0.00544634 -0.0234032
+ 4.09e+10Hz 0.00543927 -0.0234643
+ 4.1e+10Hz 0.00543215 -0.0235254
+ 4.11e+10Hz 0.00542499 -0.0235866
+ 4.12e+10Hz 0.00541777 -0.0236477
+ 4.13e+10Hz 0.00541051 -0.0237087
+ 4.14e+10Hz 0.00540321 -0.0237698
+ 4.15e+10Hz 0.00539585 -0.0238309
+ 4.16e+10Hz 0.00538845 -0.0238919
+ 4.17e+10Hz 0.00538101 -0.0239529
+ 4.18e+10Hz 0.00537351 -0.0240139
+ 4.19e+10Hz 0.00536598 -0.0240748
+ 4.2e+10Hz 0.00535839 -0.0241358
+ 4.21e+10Hz 0.00535077 -0.0241967
+ 4.22e+10Hz 0.00534309 -0.0242576
+ 4.23e+10Hz 0.00533537 -0.0243185
+ 4.24e+10Hz 0.00532761 -0.0243793
+ 4.25e+10Hz 0.00531981 -0.0244402
+ 4.26e+10Hz 0.00531196 -0.024501
+ 4.27e+10Hz 0.00530407 -0.0245618
+ 4.28e+10Hz 0.00529613 -0.0246225
+ 4.29e+10Hz 0.00528816 -0.0246833
+ 4.3e+10Hz 0.00528014 -0.024744
+ 4.31e+10Hz 0.00527208 -0.0248047
+ 4.32e+10Hz 0.00526398 -0.0248654
+ 4.33e+10Hz 0.00525584 -0.024926
+ 4.34e+10Hz 0.00524765 -0.0249866
+ 4.35e+10Hz 0.00523943 -0.0250473
+ 4.36e+10Hz 0.00523117 -0.0251078
+ 4.37e+10Hz 0.00522287 -0.0251684
+ 4.38e+10Hz 0.00521453 -0.0252289
+ 4.39e+10Hz 0.00520615 -0.0252894
+ 4.4e+10Hz 0.00519774 -0.0253498
+ 4.41e+10Hz 0.00518928 -0.0254103
+ 4.42e+10Hz 0.00518079 -0.0254707
+ 4.43e+10Hz 0.00517226 -0.025531
+ 4.44e+10Hz 0.0051637 -0.0255914
+ 4.45e+10Hz 0.0051551 -0.0256517
+ 4.46e+10Hz 0.00514647 -0.025712
+ 4.47e+10Hz 0.00513779 -0.0257723
+ 4.48e+10Hz 0.00512909 -0.0258325
+ 4.49e+10Hz 0.00512035 -0.0258927
+ 4.5e+10Hz 0.00511158 -0.0259529
+ 4.51e+10Hz 0.00510277 -0.0260131
+ 4.52e+10Hz 0.00509393 -0.0260732
+ 4.53e+10Hz 0.00508506 -0.0261333
+ 4.54e+10Hz 0.00507616 -0.0261934
+ 4.55e+10Hz 0.00506723 -0.0262534
+ 4.56e+10Hz 0.00505826 -0.0263134
+ 4.57e+10Hz 0.00504926 -0.0263734
+ 4.58e+10Hz 0.00504024 -0.0264334
+ 4.59e+10Hz 0.00503118 -0.0264933
+ 4.6e+10Hz 0.00502209 -0.0265532
+ 4.61e+10Hz 0.00501298 -0.026613
+ 4.62e+10Hz 0.00500384 -0.0266729
+ 4.63e+10Hz 0.00499466 -0.0267327
+ 4.64e+10Hz 0.00498547 -0.0267924
+ 4.65e+10Hz 0.00497624 -0.0268522
+ 4.66e+10Hz 0.00496699 -0.0269119
+ 4.67e+10Hz 0.0049577 -0.0269716
+ 4.68e+10Hz 0.0049484 -0.0270312
+ 4.69e+10Hz 0.00493907 -0.0270908
+ 4.7e+10Hz 0.00492971 -0.0271504
+ 4.71e+10Hz 0.00492032 -0.02721
+ 4.72e+10Hz 0.00491092 -0.0272695
+ 4.73e+10Hz 0.00490149 -0.027329
+ 4.74e+10Hz 0.00489203 -0.0273885
+ 4.75e+10Hz 0.00488255 -0.027448
+ 4.76e+10Hz 0.00487305 -0.0275074
+ 4.77e+10Hz 0.00486353 -0.0275668
+ 4.78e+10Hz 0.00485398 -0.0276261
+ 4.79e+10Hz 0.00484441 -0.0276855
+ 4.8e+10Hz 0.00483482 -0.0277448
+ 4.81e+10Hz 0.00482521 -0.0278041
+ 4.82e+10Hz 0.00481557 -0.0278633
+ 4.83e+10Hz 0.00480592 -0.0279225
+ 4.84e+10Hz 0.00479625 -0.0279817
+ 4.85e+10Hz 0.00478655 -0.0280409
+ 4.86e+10Hz 0.00477684 -0.0281
+ 4.87e+10Hz 0.0047671 -0.0281591
+ 4.88e+10Hz 0.00475735 -0.0282182
+ 4.89e+10Hz 0.00474758 -0.0282772
+ 4.9e+10Hz 0.00473779 -0.0283363
+ 4.91e+10Hz 0.00472798 -0.0283953
+ 4.92e+10Hz 0.00471816 -0.0284542
+ 4.93e+10Hz 0.00470831 -0.0285132
+ 4.94e+10Hz 0.00469845 -0.0285721
+ 4.95e+10Hz 0.00468857 -0.028631
+ 4.96e+10Hz 0.00467868 -0.0286899
+ 4.97e+10Hz 0.00466876 -0.0287487
+ 4.98e+10Hz 0.00465883 -0.0288075
+ 4.99e+10Hz 0.00464889 -0.0288663
+ 5e+10Hz 0.00463893 -0.0289251
+ 5.01e+10Hz 0.00462895 -0.0289838
+ 5.02e+10Hz 0.00461896 -0.0290426
+ 5.03e+10Hz 0.00460895 -0.0291012
+ 5.04e+10Hz 0.00459892 -0.0291599
+ 5.05e+10Hz 0.00458888 -0.0292186
+ 5.06e+10Hz 0.00457883 -0.0292772
+ 5.07e+10Hz 0.00456876 -0.0293358
+ 5.08e+10Hz 0.00455867 -0.0293943
+ 5.09e+10Hz 0.00454858 -0.0294529
+ 5.1e+10Hz 0.00453846 -0.0295114
+ 5.11e+10Hz 0.00452833 -0.0295699
+ 5.12e+10Hz 0.00451819 -0.0296284
+ 5.13e+10Hz 0.00450804 -0.0296869
+ 5.14e+10Hz 0.00449787 -0.0297453
+ 5.15e+10Hz 0.00448768 -0.0298038
+ 5.16e+10Hz 0.00447749 -0.0298622
+ 5.17e+10Hz 0.00446727 -0.0299205
+ 5.18e+10Hz 0.00445705 -0.0299789
+ 5.19e+10Hz 0.00444681 -0.0300372
+ 5.2e+10Hz 0.00443656 -0.0300955
+ 5.21e+10Hz 0.00442629 -0.0301538
+ 5.22e+10Hz 0.00441601 -0.0302121
+ 5.23e+10Hz 0.00440572 -0.0302704
+ 5.24e+10Hz 0.00439542 -0.0303286
+ 5.25e+10Hz 0.0043851 -0.0303868
+ 5.26e+10Hz 0.00437477 -0.030445
+ 5.27e+10Hz 0.00436442 -0.0305032
+ 5.28e+10Hz 0.00435406 -0.0305614
+ 5.29e+10Hz 0.00434369 -0.0306195
+ 5.3e+10Hz 0.0043333 -0.0306777
+ 5.31e+10Hz 0.00432291 -0.0307358
+ 5.32e+10Hz 0.0043125 -0.0307939
+ 5.33e+10Hz 0.00430207 -0.0308519
+ 5.34e+10Hz 0.00429163 -0.03091
+ 5.35e+10Hz 0.00428118 -0.030968
+ 5.36e+10Hz 0.00427071 -0.0310261
+ 5.37e+10Hz 0.00426023 -0.0310841
+ 5.38e+10Hz 0.00424974 -0.0311421
+ 5.39e+10Hz 0.00423924 -0.0312
+ 5.4e+10Hz 0.00422871 -0.031258
+ 5.41e+10Hz 0.00421818 -0.031316
+ 5.42e+10Hz 0.00420763 -0.0313739
+ 5.43e+10Hz 0.00419707 -0.0314318
+ 5.44e+10Hz 0.0041865 -0.0314897
+ 5.45e+10Hz 0.0041759 -0.0315476
+ 5.46e+10Hz 0.0041653 -0.0316055
+ 5.47e+10Hz 0.00415468 -0.0316633
+ 5.48e+10Hz 0.00414405 -0.0317211
+ 5.49e+10Hz 0.0041334 -0.031779
+ 5.5e+10Hz 0.00412274 -0.0318368
+ 5.51e+10Hz 0.00411206 -0.0318946
+ 5.52e+10Hz 0.00410137 -0.0319524
+ 5.53e+10Hz 0.00409066 -0.0320102
+ 5.54e+10Hz 0.00407994 -0.0320679
+ 5.55e+10Hz 0.0040692 -0.0321257
+ 5.56e+10Hz 0.00405845 -0.0321834
+ 5.57e+10Hz 0.00404768 -0.0322411
+ 5.58e+10Hz 0.00403689 -0.0322988
+ 5.59e+10Hz 0.00402609 -0.0323565
+ 5.6e+10Hz 0.00401527 -0.0324142
+ 5.61e+10Hz 0.00400444 -0.0324719
+ 5.62e+10Hz 0.00399359 -0.0325295
+ 5.63e+10Hz 0.00398273 -0.0325872
+ 5.64e+10Hz 0.00397184 -0.0326448
+ 5.65e+10Hz 0.00396094 -0.0327024
+ 5.66e+10Hz 0.00395003 -0.03276
+ 5.67e+10Hz 0.00393909 -0.0328176
+ 5.68e+10Hz 0.00392814 -0.0328752
+ 5.69e+10Hz 0.00391717 -0.0329328
+ 5.7e+10Hz 0.00390618 -0.0329903
+ 5.71e+10Hz 0.00389517 -0.0330479
+ 5.72e+10Hz 0.00388415 -0.0331054
+ 5.73e+10Hz 0.00387311 -0.0331629
+ 5.74e+10Hz 0.00386205 -0.0332204
+ 5.75e+10Hz 0.00385097 -0.0332779
+ 5.76e+10Hz 0.00383987 -0.0333354
+ 5.77e+10Hz 0.00382876 -0.0333929
+ 5.78e+10Hz 0.00381762 -0.0334503
+ 5.79e+10Hz 0.00380646 -0.0335078
+ 5.8e+10Hz 0.00379529 -0.0335652
+ 5.81e+10Hz 0.00378409 -0.0336227
+ 5.82e+10Hz 0.00377288 -0.0336801
+ 5.83e+10Hz 0.00376164 -0.0337375
+ 5.84e+10Hz 0.00375039 -0.0337949
+ 5.85e+10Hz 0.00373911 -0.0338523
+ 5.86e+10Hz 0.00372781 -0.0339096
+ 5.87e+10Hz 0.0037165 -0.033967
+ 5.88e+10Hz 0.00370516 -0.0340243
+ 5.89e+10Hz 0.0036938 -0.0340816
+ 5.9e+10Hz 0.00368242 -0.034139
+ 5.91e+10Hz 0.00367101 -0.0341963
+ 5.92e+10Hz 0.00365959 -0.0342536
+ 5.93e+10Hz 0.00364814 -0.0343108
+ 5.94e+10Hz 0.00363667 -0.0343681
+ 5.95e+10Hz 0.00362518 -0.0344254
+ 5.96e+10Hz 0.00361367 -0.0344826
+ 5.97e+10Hz 0.00360214 -0.0345398
+ 5.98e+10Hz 0.00359058 -0.034597
+ 5.99e+10Hz 0.003579 -0.0346542
+ 6e+10Hz 0.00356739 -0.0347114
+ 6.01e+10Hz 0.00355577 -0.0347686
+ 6.02e+10Hz 0.00354412 -0.0348258
+ 6.03e+10Hz 0.00353244 -0.0348829
+ 6.04e+10Hz 0.00352075 -0.03494
+ 6.05e+10Hz 0.00350902 -0.0349972
+ 6.06e+10Hz 0.00349728 -0.0350543
+ 6.07e+10Hz 0.00348551 -0.0351113
+ 6.08e+10Hz 0.00347372 -0.0351684
+ 6.09e+10Hz 0.0034619 -0.0352255
+ 6.1e+10Hz 0.00345006 -0.0352825
+ 6.11e+10Hz 0.00343819 -0.0353396
+ 6.12e+10Hz 0.00342631 -0.0353966
+ 6.13e+10Hz 0.00341439 -0.0354536
+ 6.14e+10Hz 0.00340245 -0.0355106
+ 6.15e+10Hz 0.00339049 -0.0355675
+ 6.16e+10Hz 0.0033785 -0.0356245
+ 6.17e+10Hz 0.00336648 -0.0356814
+ 6.18e+10Hz 0.00335445 -0.0357384
+ 6.19e+10Hz 0.00334238 -0.0357953
+ 6.2e+10Hz 0.00333029 -0.0358521
+ 6.21e+10Hz 0.00331818 -0.035909
+ 6.22e+10Hz 0.00330604 -0.0359659
+ 6.23e+10Hz 0.00329387 -0.0360227
+ 6.24e+10Hz 0.00328168 -0.0360795
+ 6.25e+10Hz 0.00326947 -0.0361363
+ 6.26e+10Hz 0.00325722 -0.0361931
+ 6.27e+10Hz 0.00324496 -0.0362499
+ 6.28e+10Hz 0.00323266 -0.0363066
+ 6.29e+10Hz 0.00322035 -0.0363634
+ 6.3e+10Hz 0.003208 -0.0364201
+ 6.31e+10Hz 0.00319563 -0.0364768
+ 6.32e+10Hz 0.00318324 -0.0365334
+ 6.33e+10Hz 0.00317081 -0.0365901
+ 6.34e+10Hz 0.00315837 -0.0366467
+ 6.35e+10Hz 0.00314589 -0.0367033
+ 6.36e+10Hz 0.0031334 -0.0367599
+ 6.37e+10Hz 0.00312087 -0.0368165
+ 6.38e+10Hz 0.00310832 -0.0368731
+ 6.39e+10Hz 0.00309575 -0.0369296
+ 6.4e+10Hz 0.00308314 -0.0369861
+ 6.41e+10Hz 0.00307052 -0.0370426
+ 6.42e+10Hz 0.00305786 -0.0370991
+ 6.43e+10Hz 0.00304519 -0.0371555
+ 6.44e+10Hz 0.00303248 -0.0372119
+ 6.45e+10Hz 0.00301975 -0.0372683
+ 6.46e+10Hz 0.003007 -0.0373247
+ 6.47e+10Hz 0.00299422 -0.0373811
+ 6.48e+10Hz 0.00298141 -0.0374374
+ 6.49e+10Hz 0.00296858 -0.0374937
+ 6.5e+10Hz 0.00295573 -0.03755
+ 6.51e+10Hz 0.00294285 -0.0376063
+ 6.52e+10Hz 0.00292994 -0.0376626
+ 6.53e+10Hz 0.00291701 -0.0377188
+ 6.54e+10Hz 0.00290405 -0.037775
+ 6.55e+10Hz 0.00289107 -0.0378312
+ 6.56e+10Hz 0.00287807 -0.0378873
+ 6.57e+10Hz 0.00286504 -0.0379434
+ 6.58e+10Hz 0.00285199 -0.0379995
+ 6.59e+10Hz 0.00283891 -0.0380556
+ 6.6e+10Hz 0.0028258 -0.0381117
+ 6.61e+10Hz 0.00281268 -0.0381677
+ 6.62e+10Hz 0.00279953 -0.0382237
+ 6.63e+10Hz 0.00278635 -0.0382797
+ 6.64e+10Hz 0.00277315 -0.0383356
+ 6.65e+10Hz 0.00275993 -0.0383916
+ 6.66e+10Hz 0.00274669 -0.0384475
+ 6.67e+10Hz 0.00273342 -0.0385033
+ 6.68e+10Hz 0.00272013 -0.0385592
+ 6.69e+10Hz 0.00270681 -0.038615
+ 6.7e+10Hz 0.00269348 -0.0386708
+ 6.71e+10Hz 0.00268012 -0.0387265
+ 6.72e+10Hz 0.00266673 -0.0387823
+ 6.73e+10Hz 0.00265333 -0.038838
+ 6.74e+10Hz 0.0026399 -0.0388937
+ 6.75e+10Hz 0.00262645 -0.0389493
+ 6.76e+10Hz 0.00261298 -0.039005
+ 6.77e+10Hz 0.00259949 -0.0390606
+ 6.78e+10Hz 0.00258598 -0.0391161
+ 6.79e+10Hz 0.00257244 -0.0391717
+ 6.8e+10Hz 0.00255888 -0.0392272
+ 6.81e+10Hz 0.00254531 -0.0392827
+ 6.82e+10Hz 0.00253171 -0.0393382
+ 6.83e+10Hz 0.00251809 -0.0393936
+ 6.84e+10Hz 0.00250445 -0.039449
+ 6.85e+10Hz 0.00249079 -0.0395044
+ 6.86e+10Hz 0.00247711 -0.0395597
+ 6.87e+10Hz 0.00246342 -0.039615
+ 6.88e+10Hz 0.0024497 -0.0396703
+ 6.89e+10Hz 0.00243596 -0.0397256
+ 6.9e+10Hz 0.0024222 -0.0397808
+ 6.91e+10Hz 0.00240843 -0.039836
+ 6.92e+10Hz 0.00239463 -0.0398912
+ 6.93e+10Hz 0.00238082 -0.0399463
+ 6.94e+10Hz 0.00236699 -0.0400014
+ 6.95e+10Hz 0.00235314 -0.0400565
+ 6.96e+10Hz 0.00233927 -0.0401116
+ 6.97e+10Hz 0.00232539 -0.0401666
+ 6.98e+10Hz 0.00231149 -0.0402216
+ 6.99e+10Hz 0.00229757 -0.0402766
+ 7e+10Hz 0.00228363 -0.0403315
+ 7.01e+10Hz 0.00226968 -0.0403864
+ 7.02e+10Hz 0.00225571 -0.0404413
+ 7.03e+10Hz 0.00224172 -0.0404961
+ 7.04e+10Hz 0.00222772 -0.0405509
+ 7.05e+10Hz 0.0022137 -0.0406057
+ 7.06e+10Hz 0.00219966 -0.0406605
+ 7.07e+10Hz 0.00218561 -0.0407152
+ 7.08e+10Hz 0.00217155 -0.0407699
+ 7.09e+10Hz 0.00215747 -0.0408245
+ 7.1e+10Hz 0.00214337 -0.0408792
+ 7.11e+10Hz 0.00212926 -0.0409338
+ 7.12e+10Hz 0.00211514 -0.0409884
+ 7.13e+10Hz 0.002101 -0.0410429
+ 7.14e+10Hz 0.00208685 -0.0410974
+ 7.15e+10Hz 0.00207268 -0.0411519
+ 7.16e+10Hz 0.0020585 -0.0412064
+ 7.17e+10Hz 0.00204431 -0.0412608
+ 7.18e+10Hz 0.0020301 -0.0413152
+ 7.19e+10Hz 0.00201588 -0.0413695
+ 7.2e+10Hz 0.00200165 -0.0414239
+ 7.21e+10Hz 0.0019874 -0.0414782
+ 7.22e+10Hz 0.00197314 -0.0415324
+ 7.23e+10Hz 0.00195887 -0.0415867
+ 7.24e+10Hz 0.00194459 -0.0416409
+ 7.25e+10Hz 0.0019303 -0.0416951
+ 7.26e+10Hz 0.00191599 -0.0417493
+ 7.27e+10Hz 0.00190167 -0.0418034
+ 7.28e+10Hz 0.00188734 -0.0418575
+ 7.29e+10Hz 0.001873 -0.0419115
+ 7.3e+10Hz 0.00185865 -0.0419656
+ 7.31e+10Hz 0.00184429 -0.0420196
+ 7.32e+10Hz 0.00182992 -0.0420736
+ 7.33e+10Hz 0.00181553 -0.0421275
+ 7.34e+10Hz 0.00180114 -0.0421815
+ 7.35e+10Hz 0.00178674 -0.0422353
+ 7.36e+10Hz 0.00177232 -0.0422892
+ 7.37e+10Hz 0.0017579 -0.0423431
+ 7.38e+10Hz 0.00174347 -0.0423969
+ 7.39e+10Hz 0.00172903 -0.0424506
+ 7.4e+10Hz 0.00171458 -0.0425044
+ 7.41e+10Hz 0.00170012 -0.0425581
+ 7.42e+10Hz 0.00168564 -0.0426118
+ 7.43e+10Hz 0.00167117 -0.0426655
+ 7.44e+10Hz 0.00165668 -0.0427191
+ 7.45e+10Hz 0.00164218 -0.0427727
+ 7.46e+10Hz 0.00162768 -0.0428263
+ 7.47e+10Hz 0.00161317 -0.0428799
+ 7.48e+10Hz 0.00159865 -0.0429334
+ 7.49e+10Hz 0.00158412 -0.0429869
+ 7.5e+10Hz 0.00156958 -0.0430404
+ 7.51e+10Hz 0.00155503 -0.0430938
+ 7.52e+10Hz 0.00154048 -0.0431473
+ 7.53e+10Hz 0.00152592 -0.0432007
+ 7.54e+10Hz 0.00151135 -0.043254
+ 7.55e+10Hz 0.00149678 -0.0433074
+ 7.56e+10Hz 0.00148219 -0.0433607
+ 7.57e+10Hz 0.0014676 -0.043414
+ 7.58e+10Hz 0.001453 -0.0434672
+ 7.59e+10Hz 0.0014384 -0.0435205
+ 7.6e+10Hz 0.00142379 -0.0435737
+ 7.61e+10Hz 0.00140917 -0.0436269
+ 7.62e+10Hz 0.00139454 -0.04368
+ 7.63e+10Hz 0.00137991 -0.0437332
+ 7.64e+10Hz 0.00136527 -0.0437863
+ 7.65e+10Hz 0.00135062 -0.0438394
+ 7.66e+10Hz 0.00133597 -0.0438924
+ 7.67e+10Hz 0.00132131 -0.0439455
+ 7.68e+10Hz 0.00130664 -0.0439985
+ 7.69e+10Hz 0.00129197 -0.0440515
+ 7.7e+10Hz 0.00127729 -0.0441045
+ 7.71e+10Hz 0.0012626 -0.0441574
+ 7.72e+10Hz 0.00124791 -0.0442103
+ 7.73e+10Hz 0.00123321 -0.0442632
+ 7.74e+10Hz 0.00121851 -0.0443161
+ 7.75e+10Hz 0.0012038 -0.0443689
+ 7.76e+10Hz 0.00118908 -0.0444217
+ 7.77e+10Hz 0.00117435 -0.0444745
+ 7.78e+10Hz 0.00115962 -0.0445273
+ 7.79e+10Hz 0.00114489 -0.0445801
+ 7.8e+10Hz 0.00113014 -0.0446328
+ 7.81e+10Hz 0.00111539 -0.0446855
+ 7.82e+10Hz 0.00110064 -0.0447382
+ 7.83e+10Hz 0.00108588 -0.0447908
+ 7.84e+10Hz 0.00107111 -0.0448435
+ 7.85e+10Hz 0.00105633 -0.0448961
+ 7.86e+10Hz 0.00104155 -0.0449487
+ 7.87e+10Hz 0.00102676 -0.0450013
+ 7.88e+10Hz 0.00101197 -0.0450538
+ 7.89e+10Hz 0.000997165 -0.0451063
+ 7.9e+10Hz 0.000982358 -0.0451589
+ 7.91e+10Hz 0.000967544 -0.0452113
+ 7.92e+10Hz 0.000952723 -0.0452638
+ 7.93e+10Hz 0.000937896 -0.0453162
+ 7.94e+10Hz 0.000923062 -0.0453687
+ 7.95e+10Hz 0.000908221 -0.0454211
+ 7.96e+10Hz 0.000893374 -0.0454734
+ 7.97e+10Hz 0.000878519 -0.0455258
+ 7.98e+10Hz 0.000863658 -0.0455781
+ 7.99e+10Hz 0.00084879 -0.0456305
+ 8e+10Hz 0.000833915 -0.0456828
+ 8.01e+10Hz 0.000819033 -0.045735
+ 8.02e+10Hz 0.000804144 -0.0457873
+ 8.03e+10Hz 0.000789247 -0.0458395
+ 8.04e+10Hz 0.000774343 -0.0458917
+ 8.05e+10Hz 0.000759432 -0.0459439
+ 8.06e+10Hz 0.000744514 -0.0459961
+ 8.07e+10Hz 0.000729588 -0.0460483
+ 8.08e+10Hz 0.000714655 -0.0461004
+ 8.09e+10Hz 0.000699714 -0.0461525
+ 8.1e+10Hz 0.000684765 -0.0462046
+ 8.11e+10Hz 0.000669809 -0.0462567
+ 8.12e+10Hz 0.000654844 -0.0463087
+ 8.13e+10Hz 0.000639872 -0.0463608
+ 8.14e+10Hz 0.000624892 -0.0464128
+ 8.15e+10Hz 0.000609903 -0.0464648
+ 8.16e+10Hz 0.000594907 -0.0465168
+ 8.17e+10Hz 0.000579902 -0.0465687
+ 8.18e+10Hz 0.000564889 -0.0466206
+ 8.19e+10Hz 0.000549867 -0.0466726
+ 8.2e+10Hz 0.000534837 -0.0467245
+ 8.21e+10Hz 0.000519798 -0.0467763
+ 8.22e+10Hz 0.00050475 -0.0468282
+ 8.23e+10Hz 0.000489694 -0.04688
+ 8.24e+10Hz 0.000474628 -0.0469319
+ 8.25e+10Hz 0.000459554 -0.0469837
+ 8.26e+10Hz 0.000444471 -0.0470354
+ 8.27e+10Hz 0.000429378 -0.0470872
+ 8.28e+10Hz 0.000414276 -0.0471389
+ 8.29e+10Hz 0.000399165 -0.0471907
+ 8.3e+10Hz 0.000384044 -0.0472424
+ 8.31e+10Hz 0.000368914 -0.047294
+ 8.32e+10Hz 0.000353774 -0.0473457
+ 8.33e+10Hz 0.000338624 -0.0473974
+ 8.34e+10Hz 0.000323465 -0.047449
+ 8.35e+10Hz 0.000308296 -0.0475006
+ 8.36e+10Hz 0.000293116 -0.0475522
+ 8.37e+10Hz 0.000277927 -0.0476037
+ 8.38e+10Hz 0.000262727 -0.0476553
+ 8.39e+10Hz 0.000247518 -0.0477068
+ 8.4e+10Hz 0.000232297 -0.0477583
+ 8.41e+10Hz 0.000217067 -0.0478098
+ 8.42e+10Hz 0.000201826 -0.0478613
+ 8.43e+10Hz 0.000186574 -0.0479127
+ 8.44e+10Hz 0.000171312 -0.0479642
+ 8.45e+10Hz 0.000156039 -0.0480156
+ 8.46e+10Hz 0.000140755 -0.0480669
+ 8.47e+10Hz 0.00012546 -0.0481183
+ 8.48e+10Hz 0.000110155 -0.0481697
+ 8.49e+10Hz 9.48382e-05 -0.048221
+ 8.5e+10Hz 7.95105e-05 -0.0482723
+ 8.51e+10Hz 6.41716e-05 -0.0483236
+ 8.52e+10Hz 4.88215e-05 -0.0483748
+ 8.53e+10Hz 3.34602e-05 -0.0484261
+ 8.54e+10Hz 1.80875e-05 -0.0484773
+ 8.55e+10Hz 2.70347e-06 -0.0485285
+ 8.56e+10Hz -1.2692e-05 -0.0485797
+ 8.57e+10Hz -2.8099e-05 -0.0486309
+ 8.58e+10Hz -4.35175e-05 -0.048682
+ 8.59e+10Hz -5.89475e-05 -0.0487331
+ 8.6e+10Hz -7.43892e-05 -0.0487842
+ 8.61e+10Hz -8.98426e-05 -0.0488353
+ 8.62e+10Hz -0.000105308 -0.0488864
+ 8.63e+10Hz -0.000120784 -0.0489374
+ 8.64e+10Hz -0.000136273 -0.0489884
+ 8.65e+10Hz -0.000151773 -0.0490394
+ 8.66e+10Hz -0.000167285 -0.0490903
+ 8.67e+10Hz -0.000182809 -0.0491413
+ 8.68e+10Hz -0.000198345 -0.0491922
+ 8.69e+10Hz -0.000213893 -0.0492431
+ 8.7e+10Hz -0.000229452 -0.049294
+ 8.71e+10Hz -0.000245024 -0.0493449
+ 8.72e+10Hz -0.000260607 -0.0493957
+ 8.73e+10Hz -0.000276202 -0.0494465
+ 8.74e+10Hz -0.000291809 -0.0494973
+ 8.75e+10Hz -0.000307429 -0.049548
+ 8.76e+10Hz -0.00032306 -0.0495988
+ 8.77e+10Hz -0.000338702 -0.0496495
+ 8.78e+10Hz -0.000354357 -0.0497002
+ 8.79e+10Hz -0.000370023 -0.0497508
+ 8.8e+10Hz -0.000385702 -0.0498015
+ 8.81e+10Hz -0.000401392 -0.0498521
+ 8.82e+10Hz -0.000417093 -0.0499027
+ 8.83e+10Hz -0.000432807 -0.0499533
+ 8.84e+10Hz -0.000448532 -0.0500038
+ 8.85e+10Hz -0.000464269 -0.0500543
+ 8.86e+10Hz -0.000480017 -0.0501048
+ 8.87e+10Hz -0.000495777 -0.0501553
+ 8.88e+10Hz -0.000511549 -0.0502058
+ 8.89e+10Hz -0.000527332 -0.0502562
+ 8.9e+10Hz -0.000543126 -0.0503066
+ 8.91e+10Hz -0.000558931 -0.050357
+ 8.92e+10Hz -0.000574748 -0.0504073
+ 8.93e+10Hz -0.000590576 -0.0504576
+ 8.94e+10Hz -0.000606415 -0.0505079
+ 8.95e+10Hz -0.000622266 -0.0505582
+ 8.96e+10Hz -0.000638127 -0.0506084
+ 8.97e+10Hz -0.000653999 -0.0506586
+ 8.98e+10Hz -0.000669881 -0.0507088
+ 8.99e+10Hz -0.000685775 -0.050759
+ 9e+10Hz -0.000701679 -0.0508091
+ 9.01e+10Hz -0.000717593 -0.0508593
+ 9.02e+10Hz -0.000733518 -0.0509093
+ 9.03e+10Hz -0.000749453 -0.0509594
+ 9.04e+10Hz -0.000765398 -0.0510094
+ 9.05e+10Hz -0.000781353 -0.0510594
+ 9.06e+10Hz -0.000797319 -0.0511094
+ 9.07e+10Hz -0.000813294 -0.0511593
+ 9.08e+10Hz -0.000829278 -0.0512093
+ 9.09e+10Hz -0.000845272 -0.0512592
+ 9.1e+10Hz -0.000861276 -0.051309
+ 9.11e+10Hz -0.000877289 -0.0513588
+ 9.12e+10Hz -0.000893311 -0.0514087
+ 9.13e+10Hz -0.000909342 -0.0514584
+ 9.14e+10Hz -0.000925382 -0.0515082
+ 9.15e+10Hz -0.00094143 -0.0515579
+ 9.16e+10Hz -0.000957488 -0.0516076
+ 9.17e+10Hz -0.000973553 -0.0516573
+ 9.18e+10Hz -0.000989627 -0.0517069
+ 9.19e+10Hz -0.00100571 -0.0517565
+ 9.2e+10Hz -0.0010218 -0.0518061
+ 9.21e+10Hz -0.0010379 -0.0518556
+ 9.22e+10Hz -0.001054 -0.0519051
+ 9.23e+10Hz -0.00107011 -0.0519546
+ 9.24e+10Hz -0.00108624 -0.0520041
+ 9.25e+10Hz -0.00110236 -0.0520535
+ 9.26e+10Hz -0.0011185 -0.0521029
+ 9.27e+10Hz -0.00113464 -0.0521523
+ 9.28e+10Hz -0.00115078 -0.0522016
+ 9.29e+10Hz -0.00116694 -0.0522509
+ 9.3e+10Hz -0.0011831 -0.0523002
+ 9.31e+10Hz -0.00119926 -0.0523494
+ 9.32e+10Hz -0.00121543 -0.0523987
+ 9.33e+10Hz -0.00123161 -0.0524479
+ 9.34e+10Hz -0.00124779 -0.052497
+ 9.35e+10Hz -0.00126398 -0.0525461
+ 9.36e+10Hz -0.00128018 -0.0525953
+ 9.37e+10Hz -0.00129637 -0.0526443
+ 9.38e+10Hz -0.00131258 -0.0526934
+ 9.39e+10Hz -0.00132878 -0.0527424
+ 9.4e+10Hz -0.001345 -0.0527913
+ 9.41e+10Hz -0.00136121 -0.0528403
+ 9.42e+10Hz -0.00137743 -0.0528892
+ 9.43e+10Hz -0.00139365 -0.0529381
+ 9.44e+10Hz -0.00140988 -0.0529869
+ 9.45e+10Hz -0.00142611 -0.0530358
+ 9.46e+10Hz -0.00144234 -0.0530846
+ 9.47e+10Hz -0.00145858 -0.0531333
+ 9.48e+10Hz -0.00147482 -0.0531821
+ 9.49e+10Hz -0.00149106 -0.0532308
+ 9.5e+10Hz -0.0015073 -0.0532794
+ 9.51e+10Hz -0.00152355 -0.0533281
+ 9.52e+10Hz -0.00153979 -0.0533767
+ 9.53e+10Hz -0.00155604 -0.0534253
+ 9.54e+10Hz -0.00157229 -0.0534738
+ 9.55e+10Hz -0.00158854 -0.0535223
+ 9.56e+10Hz -0.00160479 -0.0535708
+ 9.57e+10Hz -0.00162105 -0.0536193
+ 9.58e+10Hz -0.0016373 -0.0536677
+ 9.59e+10Hz -0.00165355 -0.0537161
+ 9.6e+10Hz -0.00166981 -0.0537645
+ 9.61e+10Hz -0.00168606 -0.0538128
+ 9.62e+10Hz -0.00170232 -0.0538611
+ 9.63e+10Hz -0.00171857 -0.0539094
+ 9.64e+10Hz -0.00173482 -0.0539576
+ 9.65e+10Hz -0.00175108 -0.0540059
+ 9.66e+10Hz -0.00176733 -0.054054
+ 9.67e+10Hz -0.00178358 -0.0541022
+ 9.68e+10Hz -0.00179983 -0.0541503
+ 9.69e+10Hz -0.00181607 -0.0541984
+ 9.7e+10Hz -0.00183232 -0.0542465
+ 9.71e+10Hz -0.00184856 -0.0542945
+ 9.72e+10Hz -0.0018648 -0.0543425
+ 9.73e+10Hz -0.00188104 -0.0543905
+ 9.74e+10Hz -0.00189728 -0.0544384
+ 9.75e+10Hz -0.00191351 -0.0544864
+ 9.76e+10Hz -0.00192975 -0.0545343
+ 9.77e+10Hz -0.00194597 -0.0545821
+ 9.78e+10Hz -0.0019622 -0.0546299
+ 9.79e+10Hz -0.00197842 -0.0546777
+ 9.8e+10Hz -0.00199464 -0.0547255
+ 9.81e+10Hz -0.00201085 -0.0547733
+ 9.82e+10Hz -0.00202706 -0.054821
+ 9.83e+10Hz -0.00204327 -0.0548687
+ 9.84e+10Hz -0.00205947 -0.0549163
+ 9.85e+10Hz -0.00207567 -0.054964
+ 9.86e+10Hz -0.00209186 -0.0550116
+ 9.87e+10Hz -0.00210805 -0.0550591
+ 9.88e+10Hz -0.00212424 -0.0551067
+ 9.89e+10Hz -0.00214042 -0.0551542
+ 9.9e+10Hz -0.00215659 -0.0552017
+ 9.91e+10Hz -0.00217276 -0.0552492
+ 9.92e+10Hz -0.00218892 -0.0552966
+ 9.93e+10Hz -0.00220508 -0.055344
+ 9.94e+10Hz -0.00222124 -0.0553914
+ 9.95e+10Hz -0.00223738 -0.0554388
+ 9.96e+10Hz -0.00225353 -0.0554861
+ 9.97e+10Hz -0.00226966 -0.0555334
+ 9.98e+10Hz -0.00228579 -0.0555807
+ 9.99e+10Hz -0.00230191 -0.0556279
+ 1e+11Hz -0.00231803 -0.0556751
+ 1.001e+11Hz -0.00233414 -0.0557223
+ 1.002e+11Hz -0.00235025 -0.0557695
+ 1.003e+11Hz -0.00236635 -0.0558167
+ 1.004e+11Hz -0.00238244 -0.0558638
+ 1.005e+11Hz -0.00239852 -0.0559109
+ 1.006e+11Hz -0.0024146 -0.0559579
+ 1.007e+11Hz -0.00243067 -0.056005
+ 1.008e+11Hz -0.00244674 -0.056052
+ 1.009e+11Hz -0.00246279 -0.056099
+ 1.01e+11Hz -0.00247884 -0.056146
+ 1.011e+11Hz -0.00249489 -0.0561929
+ 1.012e+11Hz -0.00251092 -0.0562398
+ 1.013e+11Hz -0.00252695 -0.0562867
+ 1.014e+11Hz -0.00254298 -0.0563336
+ 1.015e+11Hz -0.00255899 -0.0563804
+ 1.016e+11Hz -0.002575 -0.0564273
+ 1.017e+11Hz -0.002591 -0.0564741
+ 1.018e+11Hz -0.00260699 -0.0565209
+ 1.019e+11Hz -0.00262298 -0.0565676
+ 1.02e+11Hz -0.00263895 -0.0566144
+ 1.021e+11Hz -0.00265492 -0.0566611
+ 1.022e+11Hz -0.00267089 -0.0567078
+ 1.023e+11Hz -0.00268684 -0.0567544
+ 1.024e+11Hz -0.00270279 -0.0568011
+ 1.025e+11Hz -0.00271873 -0.0568477
+ 1.026e+11Hz -0.00273466 -0.0568943
+ 1.027e+11Hz -0.00275059 -0.0569409
+ 1.028e+11Hz -0.00276651 -0.0569874
+ 1.029e+11Hz -0.00278242 -0.0570339
+ 1.03e+11Hz -0.00279832 -0.0570804
+ 1.031e+11Hz -0.00281422 -0.0571269
+ 1.032e+11Hz -0.00283011 -0.0571734
+ 1.033e+11Hz -0.00284599 -0.0572199
+ 1.034e+11Hz -0.00286186 -0.0572663
+ 1.035e+11Hz -0.00287773 -0.0573127
+ 1.036e+11Hz -0.00289359 -0.0573591
+ 1.037e+11Hz -0.00290944 -0.0574054
+ 1.038e+11Hz -0.00292529 -0.0574518
+ 1.039e+11Hz -0.00294112 -0.0574981
+ 1.04e+11Hz -0.00295695 -0.0575444
+ 1.041e+11Hz -0.00297278 -0.0575907
+ 1.042e+11Hz -0.00298859 -0.0576369
+ 1.043e+11Hz -0.0030044 -0.0576832
+ 1.044e+11Hz -0.00302021 -0.0577294
+ 1.045e+11Hz -0.003036 -0.0577756
+ 1.046e+11Hz -0.00305179 -0.0578218
+ 1.047e+11Hz -0.00306757 -0.057868
+ 1.048e+11Hz -0.00308335 -0.0579141
+ 1.049e+11Hz -0.00309912 -0.0579602
+ 1.05e+11Hz -0.00311488 -0.0580063
+ 1.051e+11Hz -0.00313064 -0.0580524
+ 1.052e+11Hz -0.00314639 -0.0580985
+ 1.053e+11Hz -0.00316214 -0.0581446
+ 1.054e+11Hz -0.00317787 -0.0581906
+ 1.055e+11Hz -0.00319361 -0.0582366
+ 1.056e+11Hz -0.00320933 -0.0582826
+ 1.057e+11Hz -0.00322505 -0.0583286
+ 1.058e+11Hz -0.00324077 -0.0583745
+ 1.059e+11Hz -0.00325648 -0.0584204
+ 1.06e+11Hz -0.00327218 -0.0584664
+ 1.061e+11Hz -0.00328788 -0.0585123
+ 1.062e+11Hz -0.00330357 -0.0585582
+ 1.063e+11Hz -0.00331926 -0.058604
+ 1.064e+11Hz -0.00333494 -0.0586499
+ 1.065e+11Hz -0.00335062 -0.0586957
+ 1.066e+11Hz -0.0033663 -0.0587415
+ 1.067e+11Hz -0.00338196 -0.0587873
+ 1.068e+11Hz -0.00339763 -0.0588331
+ 1.069e+11Hz -0.00341329 -0.0588788
+ 1.07e+11Hz -0.00342894 -0.0589245
+ 1.071e+11Hz -0.00344459 -0.0589703
+ 1.072e+11Hz -0.00346024 -0.059016
+ 1.073e+11Hz -0.00347588 -0.0590617
+ 1.074e+11Hz -0.00349152 -0.0591073
+ 1.075e+11Hz -0.00350715 -0.059153
+ 1.076e+11Hz -0.00352278 -0.0591986
+ 1.077e+11Hz -0.00353841 -0.0592442
+ 1.078e+11Hz -0.00355403 -0.0592898
+ 1.079e+11Hz -0.00356965 -0.0593354
+ 1.08e+11Hz -0.00358526 -0.0593809
+ 1.081e+11Hz -0.00360088 -0.0594264
+ 1.082e+11Hz -0.00361649 -0.059472
+ 1.083e+11Hz -0.00363209 -0.0595174
+ 1.084e+11Hz -0.0036477 -0.0595629
+ 1.085e+11Hz -0.0036633 -0.0596084
+ 1.086e+11Hz -0.0036789 -0.0596538
+ 1.087e+11Hz -0.00369449 -0.0596993
+ 1.088e+11Hz -0.00371008 -0.0597447
+ 1.089e+11Hz -0.00372567 -0.05979
+ 1.09e+11Hz -0.00374126 -0.0598354
+ 1.091e+11Hz -0.00375685 -0.0598808
+ 1.092e+11Hz -0.00377243 -0.0599261
+ 1.093e+11Hz -0.00378801 -0.0599714
+ 1.094e+11Hz -0.00380359 -0.0600167
+ 1.095e+11Hz -0.00381917 -0.060062
+ 1.096e+11Hz -0.00383475 -0.0601072
+ 1.097e+11Hz -0.00385032 -0.0601524
+ 1.098e+11Hz -0.00386589 -0.0601976
+ 1.099e+11Hz -0.00388147 -0.0602428
+ 1.1e+11Hz -0.00389704 -0.060288
+ 1.101e+11Hz -0.0039126 -0.0603332
+ 1.102e+11Hz -0.00392817 -0.0603783
+ 1.103e+11Hz -0.00394374 -0.0604234
+ 1.104e+11Hz -0.0039593 -0.0604685
+ 1.105e+11Hz -0.00397486 -0.0605136
+ 1.106e+11Hz -0.00399043 -0.0605586
+ 1.107e+11Hz -0.00400599 -0.0606037
+ 1.108e+11Hz -0.00402155 -0.0606486
+ 1.109e+11Hz -0.00403711 -0.0606936
+ 1.11e+11Hz -0.00405266 -0.0607386
+ 1.111e+11Hz -0.00406822 -0.0607835
+ 1.112e+11Hz -0.00408378 -0.0608285
+ 1.113e+11Hz -0.00409933 -0.0608734
+ 1.114e+11Hz -0.00411489 -0.0609183
+ 1.115e+11Hz -0.00413044 -0.0609631
+ 1.116e+11Hz -0.004146 -0.0610079
+ 1.117e+11Hz -0.00416155 -0.0610528
+ 1.118e+11Hz -0.0041771 -0.0610975
+ 1.119e+11Hz -0.00419265 -0.0611423
+ 1.12e+11Hz -0.0042082 -0.061187
+ 1.121e+11Hz -0.00422375 -0.0612318
+ 1.122e+11Hz -0.0042393 -0.0612765
+ 1.123e+11Hz -0.00425485 -0.0613211
+ 1.124e+11Hz -0.0042704 -0.0613658
+ 1.125e+11Hz -0.00428595 -0.0614104
+ 1.126e+11Hz -0.00430149 -0.061455
+ 1.127e+11Hz -0.00431704 -0.0614996
+ 1.128e+11Hz -0.00433258 -0.0615441
+ 1.129e+11Hz -0.00434812 -0.0615887
+ 1.13e+11Hz -0.00436367 -0.0616332
+ 1.131e+11Hz -0.00437921 -0.0616777
+ 1.132e+11Hz -0.00439475 -0.0617221
+ 1.133e+11Hz -0.00441029 -0.0617665
+ 1.134e+11Hz -0.00442583 -0.0618109
+ 1.135e+11Hz -0.00444136 -0.0618553
+ 1.136e+11Hz -0.0044569 -0.0618997
+ 1.137e+11Hz -0.00447243 -0.061944
+ 1.138e+11Hz -0.00448796 -0.0619883
+ 1.139e+11Hz -0.00450349 -0.0620326
+ 1.14e+11Hz -0.00451902 -0.0620768
+ 1.141e+11Hz -0.00453455 -0.062121
+ 1.142e+11Hz -0.00455007 -0.0621652
+ 1.143e+11Hz -0.0045656 -0.0622094
+ 1.144e+11Hz -0.00458112 -0.0622535
+ 1.145e+11Hz -0.00459664 -0.0622976
+ 1.146e+11Hz -0.00461215 -0.0623417
+ 1.147e+11Hz -0.00462767 -0.0623858
+ 1.148e+11Hz -0.00464318 -0.0624298
+ 1.149e+11Hz -0.00465869 -0.0624738
+ 1.15e+11Hz -0.00467419 -0.0625178
+ 1.151e+11Hz -0.0046897 -0.0625617
+ 1.152e+11Hz -0.0047052 -0.0626056
+ 1.153e+11Hz -0.00472069 -0.0626495
+ 1.154e+11Hz -0.00473619 -0.0626933
+ 1.155e+11Hz -0.00475167 -0.0627372
+ 1.156e+11Hz -0.00476716 -0.062781
+ 1.157e+11Hz -0.00478264 -0.0628247
+ 1.158e+11Hz -0.00479812 -0.0628685
+ 1.159e+11Hz -0.00481359 -0.0629122
+ 1.16e+11Hz -0.00482906 -0.0629558
+ 1.161e+11Hz -0.00484452 -0.0629995
+ 1.162e+11Hz -0.00485998 -0.0630431
+ 1.163e+11Hz -0.00487543 -0.0630867
+ 1.164e+11Hz -0.00489088 -0.0631302
+ 1.165e+11Hz -0.00490632 -0.0631738
+ 1.166e+11Hz -0.00492175 -0.0632173
+ 1.167e+11Hz -0.00493718 -0.0632607
+ 1.168e+11Hz -0.00495261 -0.0633042
+ 1.169e+11Hz -0.00496802 -0.0633476
+ 1.17e+11Hz -0.00498343 -0.0633909
+ 1.171e+11Hz -0.00499884 -0.0634342
+ 1.172e+11Hz -0.00501423 -0.0634776
+ 1.173e+11Hz -0.00502962 -0.0635208
+ 1.174e+11Hz -0.005045 -0.0635641
+ 1.175e+11Hz -0.00506037 -0.0636073
+ 1.176e+11Hz -0.00507574 -0.0636505
+ 1.177e+11Hz -0.0050911 -0.0636936
+ 1.178e+11Hz -0.00510644 -0.0637367
+ 1.179e+11Hz -0.00512178 -0.0637798
+ 1.18e+11Hz -0.00513711 -0.0638229
+ 1.181e+11Hz -0.00515243 -0.0638659
+ 1.182e+11Hz -0.00516774 -0.0639089
+ 1.183e+11Hz -0.00518304 -0.0639518
+ 1.184e+11Hz -0.00519833 -0.0639947
+ 1.185e+11Hz -0.00521361 -0.0640376
+ 1.186e+11Hz -0.00522888 -0.0640805
+ 1.187e+11Hz -0.00524414 -0.0641233
+ 1.188e+11Hz -0.00525939 -0.0641661
+ 1.189e+11Hz -0.00527462 -0.0642088
+ 1.19e+11Hz -0.00528984 -0.0642516
+ 1.191e+11Hz -0.00530506 -0.0642942
+ 1.192e+11Hz -0.00532026 -0.0643369
+ 1.193e+11Hz -0.00533544 -0.0643795
+ 1.194e+11Hz -0.00535062 -0.0644221
+ 1.195e+11Hz -0.00536578 -0.0644647
+ 1.196e+11Hz -0.00538092 -0.0645072
+ 1.197e+11Hz -0.00539606 -0.0645497
+ 1.198e+11Hz -0.00541117 -0.0645922
+ 1.199e+11Hz -0.00542628 -0.0646346
+ 1.2e+11Hz -0.00544137 -0.064677
+ 1.201e+11Hz -0.00545644 -0.0647194
+ 1.202e+11Hz -0.00547151 -0.0647617
+ 1.203e+11Hz -0.00548655 -0.064804
+ 1.204e+11Hz -0.00550158 -0.0648463
+ 1.205e+11Hz -0.00551659 -0.0648885
+ 1.206e+11Hz -0.00553159 -0.0649307
+ 1.207e+11Hz -0.00554657 -0.0649729
+ 1.208e+11Hz -0.00556154 -0.0650151
+ 1.209e+11Hz -0.00557648 -0.0650572
+ 1.21e+11Hz -0.00559141 -0.0650992
+ 1.211e+11Hz -0.00560633 -0.0651413
+ 1.212e+11Hz -0.00562122 -0.0651833
+ 1.213e+11Hz -0.0056361 -0.0652253
+ 1.214e+11Hz -0.00565096 -0.0652673
+ 1.215e+11Hz -0.0056658 -0.0653092
+ 1.216e+11Hz -0.00568062 -0.0653511
+ 1.217e+11Hz -0.00569542 -0.065393
+ 1.218e+11Hz -0.00571021 -0.0654348
+ 1.219e+11Hz -0.00572497 -0.0654766
+ 1.22e+11Hz -0.00573972 -0.0655184
+ 1.221e+11Hz -0.00575444 -0.0655601
+ 1.222e+11Hz -0.00576915 -0.0656018
+ 1.223e+11Hz -0.00578383 -0.0656435
+ 1.224e+11Hz -0.0057985 -0.0656852
+ 1.225e+11Hz -0.00581314 -0.0657268
+ 1.226e+11Hz -0.00582776 -0.0657684
+ 1.227e+11Hz -0.00584236 -0.06581
+ 1.228e+11Hz -0.00585694 -0.0658515
+ 1.229e+11Hz -0.0058715 -0.065893
+ 1.23e+11Hz -0.00588604 -0.0659345
+ 1.231e+11Hz -0.00590056 -0.065976
+ 1.232e+11Hz -0.00591505 -0.0660174
+ 1.233e+11Hz -0.00592952 -0.0660588
+ 1.234e+11Hz -0.00594397 -0.0661002
+ 1.235e+11Hz -0.0059584 -0.0661415
+ 1.236e+11Hz -0.0059728 -0.0661829
+ 1.237e+11Hz -0.00598718 -0.0662242
+ 1.238e+11Hz -0.00600154 -0.0662654
+ 1.239e+11Hz -0.00601588 -0.0663067
+ 1.24e+11Hz -0.00603019 -0.0663479
+ 1.241e+11Hz -0.00604448 -0.0663891
+ 1.242e+11Hz -0.00605875 -0.0664303
+ 1.243e+11Hz -0.00607299 -0.0664714
+ 1.244e+11Hz -0.00608721 -0.0665125
+ 1.245e+11Hz -0.0061014 -0.0665536
+ 1.246e+11Hz -0.00611558 -0.0665947
+ 1.247e+11Hz -0.00612972 -0.0666358
+ 1.248e+11Hz -0.00614385 -0.0666768
+ 1.249e+11Hz -0.00615795 -0.0667178
+ 1.25e+11Hz -0.00617203 -0.0667588
+ 1.251e+11Hz -0.00618608 -0.0667997
+ 1.252e+11Hz -0.00620011 -0.0668407
+ 1.253e+11Hz -0.00621411 -0.0668816
+ 1.254e+11Hz -0.00622809 -0.0669225
+ 1.255e+11Hz -0.00624205 -0.0669634
+ 1.256e+11Hz -0.00625598 -0.0670042
+ 1.257e+11Hz -0.00626989 -0.067045
+ 1.258e+11Hz -0.00628377 -0.0670858
+ 1.259e+11Hz -0.00629763 -0.0671266
+ 1.26e+11Hz -0.00631147 -0.0671674
+ 1.261e+11Hz -0.00632528 -0.0672081
+ 1.262e+11Hz -0.00633906 -0.0672489
+ 1.263e+11Hz -0.00635283 -0.0672896
+ 1.264e+11Hz -0.00636657 -0.0673303
+ 1.265e+11Hz -0.00638029 -0.067371
+ 1.266e+11Hz -0.00639398 -0.0674116
+ 1.267e+11Hz -0.00640765 -0.0674523
+ 1.268e+11Hz -0.00642129 -0.0674929
+ 1.269e+11Hz -0.00643491 -0.0675335
+ 1.27e+11Hz -0.00644851 -0.0675741
+ 1.271e+11Hz -0.00646209 -0.0676146
+ 1.272e+11Hz -0.00647564 -0.0676552
+ 1.273e+11Hz -0.00648916 -0.0676957
+ 1.274e+11Hz -0.00650267 -0.0677362
+ 1.275e+11Hz -0.00651615 -0.0677767
+ 1.276e+11Hz -0.00652961 -0.0678172
+ 1.277e+11Hz -0.00654305 -0.0678577
+ 1.278e+11Hz -0.00655647 -0.0678982
+ 1.279e+11Hz -0.00656986 -0.0679386
+ 1.28e+11Hz -0.00658323 -0.0679791
+ 1.281e+11Hz -0.00659658 -0.0680195
+ 1.282e+11Hz -0.00660991 -0.0680599
+ 1.283e+11Hz -0.00662321 -0.0681003
+ 1.284e+11Hz -0.0066365 -0.0681406
+ 1.285e+11Hz -0.00664976 -0.068181
+ 1.286e+11Hz -0.006663 -0.0682214
+ 1.287e+11Hz -0.00667623 -0.0682617
+ 1.288e+11Hz -0.00668943 -0.068302
+ 1.289e+11Hz -0.00670261 -0.0683423
+ 1.29e+11Hz -0.00671577 -0.0683826
+ 1.291e+11Hz -0.00672891 -0.0684229
+ 1.292e+11Hz -0.00674204 -0.0684632
+ 1.293e+11Hz -0.00675514 -0.0685035
+ 1.294e+11Hz -0.00676822 -0.0685437
+ 1.295e+11Hz -0.00678129 -0.068584
+ 1.296e+11Hz -0.00679434 -0.0686242
+ 1.297e+11Hz -0.00680737 -0.0686644
+ 1.298e+11Hz -0.00682038 -0.0687046
+ 1.299e+11Hz -0.00683337 -0.0687448
+ 1.3e+11Hz -0.00684635 -0.068785
+ 1.301e+11Hz -0.00685931 -0.0688252
+ 1.302e+11Hz -0.00687225 -0.0688654
+ 1.303e+11Hz -0.00688518 -0.0689055
+ 1.304e+11Hz -0.00689809 -0.0689457
+ 1.305e+11Hz -0.00691098 -0.0689858
+ 1.306e+11Hz -0.00692386 -0.069026
+ 1.307e+11Hz -0.00693672 -0.0690661
+ 1.308e+11Hz -0.00694957 -0.0691062
+ 1.309e+11Hz -0.00696241 -0.0691463
+ 1.31e+11Hz -0.00697523 -0.0691864
+ 1.311e+11Hz -0.00698803 -0.0692265
+ 1.312e+11Hz -0.00700083 -0.0692665
+ 1.313e+11Hz -0.00701361 -0.0693066
+ 1.314e+11Hz -0.00702637 -0.0693466
+ 1.315e+11Hz -0.00703913 -0.0693867
+ 1.316e+11Hz -0.00705187 -0.0694267
+ 1.317e+11Hz -0.0070646 -0.0694667
+ 1.318e+11Hz -0.00707732 -0.0695068
+ 1.319e+11Hz -0.00709002 -0.0695468
+ 1.32e+11Hz -0.00710272 -0.0695868
+ 1.321e+11Hz -0.00711541 -0.0696267
+ 1.322e+11Hz -0.00712808 -0.0696667
+ 1.323e+11Hz -0.00714075 -0.0697067
+ 1.324e+11Hz -0.0071534 -0.0697466
+ 1.325e+11Hz -0.00716605 -0.0697866
+ 1.326e+11Hz -0.00717869 -0.0698265
+ 1.327e+11Hz -0.00719132 -0.0698664
+ 1.328e+11Hz -0.00720394 -0.0699064
+ 1.329e+11Hz -0.00721655 -0.0699463
+ 1.33e+11Hz -0.00722916 -0.0699862
+ 1.331e+11Hz -0.00724175 -0.070026
+ 1.332e+11Hz -0.00725434 -0.0700659
+ 1.333e+11Hz -0.00726693 -0.0701058
+ 1.334e+11Hz -0.00727951 -0.0701456
+ 1.335e+11Hz -0.00729208 -0.0701855
+ 1.336e+11Hz -0.00730464 -0.0702253
+ 1.337e+11Hz -0.0073172 -0.0702651
+ 1.338e+11Hz -0.00732976 -0.0703049
+ 1.339e+11Hz -0.00734231 -0.0703447
+ 1.34e+11Hz -0.00735485 -0.0703845
+ 1.341e+11Hz -0.00736739 -0.0704243
+ 1.342e+11Hz -0.00737993 -0.070464
+ 1.343e+11Hz -0.00739246 -0.0705038
+ 1.344e+11Hz -0.00740499 -0.0705435
+ 1.345e+11Hz -0.00741752 -0.0705832
+ 1.346e+11Hz -0.00743004 -0.0706229
+ 1.347e+11Hz -0.00744256 -0.0706626
+ 1.348e+11Hz -0.00745508 -0.0707023
+ 1.349e+11Hz -0.00746759 -0.0707419
+ 1.35e+11Hz -0.0074801 -0.0707816
+ 1.351e+11Hz -0.00749261 -0.0708212
+ 1.352e+11Hz -0.00750512 -0.0708608
+ 1.353e+11Hz -0.00751763 -0.0709004
+ 1.354e+11Hz -0.00753013 -0.07094
+ 1.355e+11Hz -0.00754264 -0.0709796
+ 1.356e+11Hz -0.00755514 -0.0710191
+ 1.357e+11Hz -0.00756764 -0.0710586
+ 1.358e+11Hz -0.00758014 -0.0710981
+ 1.359e+11Hz -0.00759265 -0.0711376
+ 1.36e+11Hz -0.00760515 -0.0711771
+ 1.361e+11Hz -0.00761765 -0.0712166
+ 1.362e+11Hz -0.00763014 -0.071256
+ 1.363e+11Hz -0.00764264 -0.0712954
+ 1.364e+11Hz -0.00765514 -0.0713348
+ 1.365e+11Hz -0.00766764 -0.0713742
+ 1.366e+11Hz -0.00768014 -0.0714136
+ 1.367e+11Hz -0.00769264 -0.0714529
+ 1.368e+11Hz -0.00770514 -0.0714922
+ 1.369e+11Hz -0.00771764 -0.0715315
+ 1.37e+11Hz -0.00773014 -0.0715708
+ 1.371e+11Hz -0.00774264 -0.0716101
+ 1.372e+11Hz -0.00775514 -0.0716493
+ 1.373e+11Hz -0.00776764 -0.0716885
+ 1.374e+11Hz -0.00778014 -0.0717277
+ 1.375e+11Hz -0.00779264 -0.0717668
+ 1.376e+11Hz -0.00780514 -0.071806
+ 1.377e+11Hz -0.00781764 -0.0718451
+ 1.378e+11Hz -0.00783014 -0.0718842
+ 1.379e+11Hz -0.00784264 -0.0719232
+ 1.38e+11Hz -0.00785514 -0.0719623
+ 1.381e+11Hz -0.00786764 -0.0720013
+ 1.382e+11Hz -0.00788014 -0.0720402
+ 1.383e+11Hz -0.00789264 -0.0720792
+ 1.384e+11Hz -0.00790513 -0.0721181
+ 1.385e+11Hz -0.00791763 -0.072157
+ 1.386e+11Hz -0.00793012 -0.0721959
+ 1.387e+11Hz -0.00794262 -0.0722347
+ 1.388e+11Hz -0.00795511 -0.0722735
+ 1.389e+11Hz -0.0079676 -0.0723123
+ 1.39e+11Hz -0.00798009 -0.0723511
+ 1.391e+11Hz -0.00799258 -0.0723898
+ 1.392e+11Hz -0.00800506 -0.0724285
+ 1.393e+11Hz -0.00801754 -0.0724671
+ 1.394e+11Hz -0.00803002 -0.0725057
+ 1.395e+11Hz -0.0080425 -0.0725443
+ 1.396e+11Hz -0.00805497 -0.0725829
+ 1.397e+11Hz -0.00806744 -0.0726214
+ 1.398e+11Hz -0.0080799 -0.0726599
+ 1.399e+11Hz -0.00809236 -0.0726984
+ 1.4e+11Hz -0.00810481 -0.0727368
+ 1.401e+11Hz -0.00811726 -0.0727752
+ 1.402e+11Hz -0.00812971 -0.0728136
+ 1.403e+11Hz -0.00814214 -0.0728519
+ 1.404e+11Hz -0.00815458 -0.0728902
+ 1.405e+11Hz -0.008167 -0.0729284
+ 1.406e+11Hz -0.00817942 -0.0729666
+ 1.407e+11Hz -0.00819182 -0.0730048
+ 1.408e+11Hz -0.00820423 -0.073043
+ 1.409e+11Hz -0.00821662 -0.0730811
+ 1.41e+11Hz -0.008229 -0.0731192
+ 1.411e+11Hz -0.00824138 -0.0731572
+ 1.412e+11Hz -0.00825374 -0.0731952
+ 1.413e+11Hz -0.00826609 -0.0732332
+ 1.414e+11Hz -0.00827844 -0.0732711
+ 1.415e+11Hz -0.00829077 -0.073309
+ 1.416e+11Hz -0.00830308 -0.0733468
+ 1.417e+11Hz -0.00831539 -0.0733846
+ 1.418e+11Hz -0.00832768 -0.0734224
+ 1.419e+11Hz -0.00833996 -0.0734602
+ 1.42e+11Hz -0.00835223 -0.0734979
+ 1.421e+11Hz -0.00836448 -0.0735355
+ 1.422e+11Hz -0.00837672 -0.0735732
+ 1.423e+11Hz -0.00838894 -0.0736107
+ 1.424e+11Hz -0.00840114 -0.0736483
+ 1.425e+11Hz -0.00841332 -0.0736858
+ 1.426e+11Hz -0.00842549 -0.0737233
+ 1.427e+11Hz -0.00843764 -0.0737607
+ 1.428e+11Hz -0.00844977 -0.0737981
+ 1.429e+11Hz -0.00846188 -0.0738354
+ 1.43e+11Hz -0.00847397 -0.0738728
+ 1.431e+11Hz -0.00848604 -0.07391
+ 1.432e+11Hz -0.00849809 -0.0739473
+ 1.433e+11Hz -0.00851012 -0.0739845
+ 1.434e+11Hz -0.00852212 -0.0740216
+ 1.435e+11Hz -0.0085341 -0.0740587
+ 1.436e+11Hz -0.00854606 -0.0740958
+ 1.437e+11Hz -0.00855799 -0.0741329
+ 1.438e+11Hz -0.0085699 -0.0741699
+ 1.439e+11Hz -0.00858178 -0.0742069
+ 1.44e+11Hz -0.00859363 -0.0742438
+ 1.441e+11Hz -0.00860546 -0.0742807
+ 1.442e+11Hz -0.00861725 -0.0743175
+ 1.443e+11Hz -0.00862902 -0.0743544
+ 1.444e+11Hz -0.00864076 -0.0743912
+ 1.445e+11Hz -0.00865247 -0.0744279
+ 1.446e+11Hz -0.00866415 -0.0744646
+ 1.447e+11Hz -0.0086758 -0.0745013
+ 1.448e+11Hz -0.00868742 -0.074538
+ 1.449e+11Hz -0.008699 -0.0745746
+ 1.45e+11Hz -0.00871056 -0.0746111
+ 1.451e+11Hz -0.00872207 -0.0746477
+ 1.452e+11Hz -0.00873356 -0.0746842
+ 1.453e+11Hz -0.00874501 -0.0747207
+ 1.454e+11Hz -0.00875642 -0.0747571
+ 1.455e+11Hz -0.00876779 -0.0747935
+ 1.456e+11Hz -0.00877913 -0.0748299
+ 1.457e+11Hz -0.00879043 -0.0748662
+ 1.458e+11Hz -0.0088017 -0.0749026
+ 1.459e+11Hz -0.00881292 -0.0749389
+ 1.46e+11Hz -0.00882411 -0.0749751
+ 1.461e+11Hz -0.00883525 -0.0750114
+ 1.462e+11Hz -0.00884636 -0.0750476
+ 1.463e+11Hz -0.00885742 -0.0750837
+ 1.464e+11Hz -0.00886845 -0.0751199
+ 1.465e+11Hz -0.00887943 -0.075156
+ 1.466e+11Hz -0.00889036 -0.0751921
+ 1.467e+11Hz -0.00890126 -0.0752282
+ 1.468e+11Hz -0.00891211 -0.0752642
+ 1.469e+11Hz -0.00892292 -0.0753002
+ 1.47e+11Hz -0.00893368 -0.0753362
+ 1.471e+11Hz -0.0089444 -0.0753722
+ 1.472e+11Hz -0.00895507 -0.0754082
+ 1.473e+11Hz -0.0089657 -0.0754441
+ 1.474e+11Hz -0.00897628 -0.07548
+ 1.475e+11Hz -0.00898681 -0.0755159
+ 1.476e+11Hz -0.0089973 -0.0755518
+ 1.477e+11Hz -0.00900773 -0.0755877
+ 1.478e+11Hz -0.00901812 -0.0756235
+ 1.479e+11Hz -0.00902847 -0.0756593
+ 1.48e+11Hz -0.00903876 -0.0756951
+ 1.481e+11Hz -0.00904901 -0.0757309
+ 1.482e+11Hz -0.0090592 -0.0757667
+ 1.483e+11Hz -0.00906935 -0.0758025
+ 1.484e+11Hz -0.00907945 -0.0758383
+ 1.485e+11Hz -0.00908949 -0.075874
+ 1.486e+11Hz -0.00909949 -0.0759098
+ 1.487e+11Hz -0.00910944 -0.0759455
+ 1.488e+11Hz -0.00911933 -0.0759813
+ 1.489e+11Hz -0.00912918 -0.076017
+ 1.49e+11Hz -0.00913897 -0.0760527
+ 1.491e+11Hz -0.00914872 -0.0760884
+ 1.492e+11Hz -0.00915841 -0.0761241
+ 1.493e+11Hz -0.00916805 -0.0761598
+ 1.494e+11Hz -0.00917764 -0.0761955
+ 1.495e+11Hz -0.00918718 -0.0762312
+ 1.496e+11Hz -0.00919667 -0.076267
+ 1.497e+11Hz -0.00920611 -0.0763027
+ 1.498e+11Hz -0.0092155 -0.0763384
+ 1.499e+11Hz -0.00922483 -0.0763741
+ 1.5e+11Hz -0.00923411 -0.0764098
+ ]

A12 %vd(20 3) %vd(12, 3) xfer2
.model xfer2 xfer R_I=true table=[
+ 0Hz 0.996062 0
+ 1e+08Hz 0.996062 -0.000713128
+ 2e+08Hz 0.99606 -0.00142625
+ 3e+08Hz 0.996058 -0.00213934
+ 4e+08Hz 0.996054 -0.0028524
+ 5e+08Hz 0.99605 -0.00356542
+ 6e+08Hz 0.996045 -0.00427839
+ 7e+08Hz 0.996039 -0.00499129
+ 8e+08Hz 0.996031 -0.00570411
+ 9e+08Hz 0.996023 -0.00641685
+ 1e+09Hz 0.996014 -0.0071295
+ 1.1e+09Hz 0.996004 -0.00784203
+ 1.2e+09Hz 0.995993 -0.00855445
+ 1.3e+09Hz 0.995981 -0.00926674
+ 1.4e+09Hz 0.995968 -0.00997889
+ 1.5e+09Hz 0.995954 -0.0106909
+ 1.6e+09Hz 0.99594 -0.0114027
+ 1.7e+09Hz 0.995924 -0.0121144
+ 1.8e+09Hz 0.995907 -0.0128259
+ 1.9e+09Hz 0.99589 -0.0135372
+ 2e+09Hz 0.995872 -0.0142483
+ 2.1e+09Hz 0.995852 -0.0149593
+ 2.2e+09Hz 0.995832 -0.0156699
+ 2.3e+09Hz 0.995811 -0.0163804
+ 2.4e+09Hz 0.995789 -0.0170906
+ 2.5e+09Hz 0.995766 -0.0178006
+ 2.6e+09Hz 0.995742 -0.0185103
+ 2.7e+09Hz 0.995718 -0.0192198
+ 2.8e+09Hz 0.995692 -0.019929
+ 2.9e+09Hz 0.995665 -0.0206379
+ 3e+09Hz 0.995638 -0.0213466
+ 3.1e+09Hz 0.99561 -0.0220549
+ 3.2e+09Hz 0.995581 -0.022763
+ 3.3e+09Hz 0.995551 -0.0234707
+ 3.4e+09Hz 0.995521 -0.0241781
+ 3.5e+09Hz 0.995489 -0.0248852
+ 3.6e+09Hz 0.995457 -0.025592
+ 3.7e+09Hz 0.995424 -0.0262984
+ 3.8e+09Hz 0.99539 -0.0270045
+ 3.9e+09Hz 0.995355 -0.0277102
+ 4e+09Hz 0.99532 -0.0284156
+ 4.1e+09Hz 0.995283 -0.0291206
+ 4.2e+09Hz 0.995247 -0.0298253
+ 4.3e+09Hz 0.995209 -0.0305296
+ 4.4e+09Hz 0.99517 -0.0312334
+ 4.5e+09Hz 0.995131 -0.031937
+ 4.6e+09Hz 0.995091 -0.0326401
+ 4.7e+09Hz 0.99505 -0.0333428
+ 4.8e+09Hz 0.995009 -0.0340452
+ 4.9e+09Hz 0.994966 -0.0347471
+ 5e+09Hz 0.994924 -0.0354486
+ 5.1e+09Hz 0.99488 -0.0361498
+ 5.2e+09Hz 0.994836 -0.0368504
+ 5.3e+09Hz 0.994791 -0.0375508
+ 5.4e+09Hz 0.994745 -0.0382506
+ 5.5e+09Hz 0.994699 -0.0389501
+ 5.6e+09Hz 0.994652 -0.0396491
+ 5.7e+09Hz 0.994605 -0.0403477
+ 5.8e+09Hz 0.994557 -0.0410459
+ 5.9e+09Hz 0.994508 -0.0417437
+ 6e+09Hz 0.994459 -0.042441
+ 6.1e+09Hz 0.994409 -0.0431379
+ 6.2e+09Hz 0.994358 -0.0438343
+ 6.3e+09Hz 0.994307 -0.0445303
+ 6.4e+09Hz 0.994255 -0.0452259
+ 6.5e+09Hz 0.994203 -0.0459211
+ 6.6e+09Hz 0.99415 -0.0466158
+ 6.7e+09Hz 0.994097 -0.0473101
+ 6.8e+09Hz 0.994043 -0.0480039
+ 6.9e+09Hz 0.993988 -0.0486973
+ 7e+09Hz 0.993933 -0.0493903
+ 7.1e+09Hz 0.993878 -0.0500829
+ 7.2e+09Hz 0.993822 -0.050775
+ 7.3e+09Hz 0.993765 -0.0514667
+ 7.4e+09Hz 0.993708 -0.0521579
+ 7.5e+09Hz 0.993651 -0.0528487
+ 7.6e+09Hz 0.993593 -0.0535392
+ 7.7e+09Hz 0.993534 -0.0542291
+ 7.8e+09Hz 0.993476 -0.0549187
+ 7.9e+09Hz 0.993416 -0.0556078
+ 8e+09Hz 0.993357 -0.0562966
+ 8.1e+09Hz 0.993297 -0.0569849
+ 8.2e+09Hz 0.993236 -0.0576728
+ 8.3e+09Hz 0.993175 -0.0583603
+ 8.4e+09Hz 0.993113 -0.0590473
+ 8.5e+09Hz 0.993052 -0.059734
+ 8.6e+09Hz 0.992989 -0.0604203
+ 8.7e+09Hz 0.992927 -0.0611062
+ 8.8e+09Hz 0.992864 -0.0617917
+ 8.9e+09Hz 0.992801 -0.0624769
+ 9e+09Hz 0.992737 -0.0631616
+ 9.1e+09Hz 0.992673 -0.0638459
+ 9.2e+09Hz 0.992608 -0.0645299
+ 9.3e+09Hz 0.992544 -0.0652136
+ 9.4e+09Hz 0.992478 -0.0658968
+ 9.5e+09Hz 0.992413 -0.0665797
+ 9.6e+09Hz 0.992347 -0.0672623
+ 9.7e+09Hz 0.992281 -0.0679445
+ 9.8e+09Hz 0.992215 -0.0686263
+ 9.9e+09Hz 0.992148 -0.0693078
+ 1e+10Hz 0.992081 -0.069989
+ 1.01e+10Hz 0.992013 -0.0706699
+ 1.02e+10Hz 0.991946 -0.0713504
+ 1.03e+10Hz 0.991878 -0.0720306
+ 1.04e+10Hz 0.991809 -0.0727105
+ 1.05e+10Hz 0.991741 -0.0733901
+ 1.06e+10Hz 0.991672 -0.0740694
+ 1.07e+10Hz 0.991603 -0.0747484
+ 1.08e+10Hz 0.991533 -0.0754271
+ 1.09e+10Hz 0.991464 -0.0761055
+ 1.1e+10Hz 0.991394 -0.0767837
+ 1.11e+10Hz 0.991323 -0.0774616
+ 1.12e+10Hz 0.991253 -0.0781392
+ 1.13e+10Hz 0.991182 -0.0788165
+ 1.14e+10Hz 0.991111 -0.0794936
+ 1.15e+10Hz 0.99104 -0.0801705
+ 1.16e+10Hz 0.990968 -0.0808471
+ 1.17e+10Hz 0.990896 -0.0815234
+ 1.18e+10Hz 0.990824 -0.0821996
+ 1.19e+10Hz 0.990752 -0.0828755
+ 1.2e+10Hz 0.99068 -0.0835512
+ 1.21e+10Hz 0.990607 -0.0842267
+ 1.22e+10Hz 0.990534 -0.0849019
+ 1.23e+10Hz 0.99046 -0.085577
+ 1.24e+10Hz 0.990387 -0.0862519
+ 1.25e+10Hz 0.990313 -0.0869266
+ 1.26e+10Hz 0.990239 -0.0876011
+ 1.27e+10Hz 0.990165 -0.0882754
+ 1.28e+10Hz 0.99009 -0.0889496
+ 1.29e+10Hz 0.990015 -0.0896235
+ 1.3e+10Hz 0.98994 -0.0902974
+ 1.31e+10Hz 0.989865 -0.0909711
+ 1.32e+10Hz 0.98979 -0.0916446
+ 1.33e+10Hz 0.989714 -0.092318
+ 1.34e+10Hz 0.989638 -0.0929912
+ 1.35e+10Hz 0.989562 -0.0936643
+ 1.36e+10Hz 0.989485 -0.0943373
+ 1.37e+10Hz 0.989409 -0.0950102
+ 1.38e+10Hz 0.989332 -0.0956829
+ 1.39e+10Hz 0.989254 -0.0963556
+ 1.4e+10Hz 0.989177 -0.0970281
+ 1.41e+10Hz 0.989099 -0.0977005
+ 1.42e+10Hz 0.989021 -0.0983729
+ 1.43e+10Hz 0.988943 -0.0990451
+ 1.44e+10Hz 0.988864 -0.0997173
+ 1.45e+10Hz 0.988786 -0.100389
+ 1.46e+10Hz 0.988707 -0.101061
+ 1.47e+10Hz 0.988627 -0.101733
+ 1.48e+10Hz 0.988548 -0.102405
+ 1.49e+10Hz 0.988468 -0.103077
+ 1.5e+10Hz 0.988388 -0.103749
+ 1.51e+10Hz 0.988308 -0.10442
+ 1.52e+10Hz 0.988227 -0.105092
+ 1.53e+10Hz 0.988146 -0.105763
+ 1.54e+10Hz 0.988065 -0.106435
+ 1.55e+10Hz 0.987984 -0.107106
+ 1.56e+10Hz 0.987902 -0.107778
+ 1.57e+10Hz 0.98782 -0.108449
+ 1.58e+10Hz 0.987737 -0.109121
+ 1.59e+10Hz 0.987655 -0.109792
+ 1.6e+10Hz 0.987572 -0.110463
+ 1.61e+10Hz 0.987489 -0.111135
+ 1.62e+10Hz 0.987405 -0.111806
+ 1.63e+10Hz 0.987321 -0.112477
+ 1.64e+10Hz 0.987237 -0.113149
+ 1.65e+10Hz 0.987153 -0.11382
+ 1.66e+10Hz 0.987068 -0.114491
+ 1.67e+10Hz 0.986983 -0.115162
+ 1.68e+10Hz 0.986897 -0.115834
+ 1.69e+10Hz 0.986812 -0.116505
+ 1.7e+10Hz 0.986726 -0.117176
+ 1.71e+10Hz 0.986639 -0.117847
+ 1.72e+10Hz 0.986553 -0.118519
+ 1.73e+10Hz 0.986466 -0.11919
+ 1.74e+10Hz 0.986378 -0.119861
+ 1.75e+10Hz 0.98629 -0.120532
+ 1.76e+10Hz 0.986202 -0.121204
+ 1.77e+10Hz 0.986114 -0.121875
+ 1.78e+10Hz 0.986025 -0.122546
+ 1.79e+10Hz 0.985936 -0.123218
+ 1.8e+10Hz 0.985846 -0.123889
+ 1.81e+10Hz 0.985756 -0.12456
+ 1.82e+10Hz 0.985666 -0.125232
+ 1.83e+10Hz 0.985575 -0.125903
+ 1.84e+10Hz 0.985484 -0.126575
+ 1.85e+10Hz 0.985393 -0.127246
+ 1.86e+10Hz 0.985301 -0.127918
+ 1.87e+10Hz 0.985209 -0.128589
+ 1.88e+10Hz 0.985116 -0.129261
+ 1.89e+10Hz 0.985023 -0.129932
+ 1.9e+10Hz 0.98493 -0.130604
+ 1.91e+10Hz 0.984836 -0.131275
+ 1.92e+10Hz 0.984742 -0.131947
+ 1.93e+10Hz 0.984647 -0.132619
+ 1.94e+10Hz 0.984552 -0.13329
+ 1.95e+10Hz 0.984457 -0.133962
+ 1.96e+10Hz 0.984361 -0.134633
+ 1.97e+10Hz 0.984265 -0.135305
+ 1.98e+10Hz 0.984168 -0.135977
+ 1.99e+10Hz 0.984071 -0.136649
+ 2e+10Hz 0.983973 -0.137321
+ 2.01e+10Hz 0.983875 -0.137992
+ 2.02e+10Hz 0.983777 -0.138664
+ 2.03e+10Hz 0.983678 -0.139336
+ 2.04e+10Hz 0.983579 -0.140008
+ 2.05e+10Hz 0.983479 -0.14068
+ 2.06e+10Hz 0.983379 -0.141351
+ 2.07e+10Hz 0.983278 -0.142023
+ 2.08e+10Hz 0.983177 -0.142695
+ 2.09e+10Hz 0.983075 -0.143367
+ 2.1e+10Hz 0.982973 -0.144039
+ 2.11e+10Hz 0.982871 -0.144711
+ 2.12e+10Hz 0.982768 -0.145383
+ 2.13e+10Hz 0.982664 -0.146055
+ 2.14e+10Hz 0.98256 -0.146727
+ 2.15e+10Hz 0.982456 -0.147398
+ 2.16e+10Hz 0.982351 -0.14807
+ 2.17e+10Hz 0.982246 -0.148742
+ 2.18e+10Hz 0.98214 -0.149414
+ 2.19e+10Hz 0.982034 -0.150086
+ 2.2e+10Hz 0.981927 -0.150758
+ 2.21e+10Hz 0.98182 -0.15143
+ 2.22e+10Hz 0.981712 -0.152101
+ 2.23e+10Hz 0.981604 -0.152773
+ 2.24e+10Hz 0.981495 -0.153445
+ 2.25e+10Hz 0.981386 -0.154117
+ 2.26e+10Hz 0.981276 -0.154788
+ 2.27e+10Hz 0.981166 -0.15546
+ 2.28e+10Hz 0.981055 -0.156132
+ 2.29e+10Hz 0.980944 -0.156804
+ 2.3e+10Hz 0.980832 -0.157475
+ 2.31e+10Hz 0.98072 -0.158147
+ 2.32e+10Hz 0.980607 -0.158818
+ 2.33e+10Hz 0.980494 -0.15949
+ 2.34e+10Hz 0.980381 -0.160161
+ 2.35e+10Hz 0.980267 -0.160833
+ 2.36e+10Hz 0.980152 -0.161504
+ 2.37e+10Hz 0.980037 -0.162176
+ 2.38e+10Hz 0.979921 -0.162847
+ 2.39e+10Hz 0.979805 -0.163518
+ 2.4e+10Hz 0.979688 -0.164189
+ 2.41e+10Hz 0.979571 -0.16486
+ 2.42e+10Hz 0.979453 -0.165531
+ 2.43e+10Hz 0.979335 -0.166202
+ 2.44e+10Hz 0.979216 -0.166873
+ 2.45e+10Hz 0.979097 -0.167544
+ 2.46e+10Hz 0.978977 -0.168215
+ 2.47e+10Hz 0.978857 -0.168886
+ 2.48e+10Hz 0.978736 -0.169556
+ 2.49e+10Hz 0.978615 -0.170227
+ 2.5e+10Hz 0.978493 -0.170898
+ 2.51e+10Hz 0.978371 -0.171568
+ 2.52e+10Hz 0.978248 -0.172238
+ 2.53e+10Hz 0.978125 -0.172909
+ 2.54e+10Hz 0.978001 -0.173579
+ 2.55e+10Hz 0.977877 -0.174249
+ 2.56e+10Hz 0.977752 -0.174919
+ 2.57e+10Hz 0.977627 -0.175589
+ 2.58e+10Hz 0.977501 -0.176259
+ 2.59e+10Hz 0.977375 -0.176928
+ 2.6e+10Hz 0.977248 -0.177598
+ 2.61e+10Hz 0.977121 -0.178267
+ 2.62e+10Hz 0.976993 -0.178937
+ 2.63e+10Hz 0.976865 -0.179606
+ 2.64e+10Hz 0.976736 -0.180276
+ 2.65e+10Hz 0.976606 -0.180945
+ 2.66e+10Hz 0.976477 -0.181614
+ 2.67e+10Hz 0.976346 -0.182282
+ 2.68e+10Hz 0.976215 -0.182951
+ 2.69e+10Hz 0.976084 -0.18362
+ 2.7e+10Hz 0.975952 -0.184288
+ 2.71e+10Hz 0.97582 -0.184957
+ 2.72e+10Hz 0.975687 -0.185625
+ 2.73e+10Hz 0.975554 -0.186294
+ 2.74e+10Hz 0.97542 -0.186962
+ 2.75e+10Hz 0.975286 -0.18763
+ 2.76e+10Hz 0.975151 -0.188297
+ 2.77e+10Hz 0.975016 -0.188965
+ 2.78e+10Hz 0.97488 -0.189633
+ 2.79e+10Hz 0.974744 -0.1903
+ 2.8e+10Hz 0.974607 -0.190967
+ 2.81e+10Hz 0.97447 -0.191635
+ 2.82e+10Hz 0.974332 -0.192302
+ 2.83e+10Hz 0.974194 -0.192969
+ 2.84e+10Hz 0.974056 -0.193635
+ 2.85e+10Hz 0.973917 -0.194302
+ 2.86e+10Hz 0.973777 -0.194968
+ 2.87e+10Hz 0.973637 -0.195635
+ 2.88e+10Hz 0.973496 -0.196301
+ 2.89e+10Hz 0.973355 -0.196967
+ 2.9e+10Hz 0.973214 -0.197633
+ 2.91e+10Hz 0.973072 -0.198299
+ 2.92e+10Hz 0.97293 -0.198965
+ 2.93e+10Hz 0.972787 -0.19963
+ 2.94e+10Hz 0.972643 -0.200296
+ 2.95e+10Hz 0.9725 -0.200961
+ 2.96e+10Hz 0.972355 -0.201626
+ 2.97e+10Hz 0.972211 -0.202291
+ 2.98e+10Hz 0.972066 -0.202956
+ 2.99e+10Hz 0.97192 -0.203621
+ 3e+10Hz 0.971774 -0.204285
+ 3.01e+10Hz 0.971627 -0.20495
+ 3.02e+10Hz 0.97148 -0.205614
+ 3.03e+10Hz 0.971333 -0.206278
+ 3.04e+10Hz 0.971185 -0.206942
+ 3.05e+10Hz 0.971036 -0.207606
+ 3.06e+10Hz 0.970888 -0.208269
+ 3.07e+10Hz 0.970738 -0.208933
+ 3.08e+10Hz 0.970589 -0.209596
+ 3.09e+10Hz 0.970438 -0.21026
+ 3.1e+10Hz 0.970288 -0.210923
+ 3.11e+10Hz 0.970137 -0.211586
+ 3.12e+10Hz 0.969985 -0.212249
+ 3.13e+10Hz 0.969834 -0.212911
+ 3.14e+10Hz 0.969681 -0.213574
+ 3.15e+10Hz 0.969528 -0.214236
+ 3.16e+10Hz 0.969375 -0.214898
+ 3.17e+10Hz 0.969221 -0.21556
+ 3.18e+10Hz 0.969067 -0.216222
+ 3.19e+10Hz 0.968913 -0.216884
+ 3.2e+10Hz 0.968758 -0.217546
+ 3.21e+10Hz 0.968603 -0.218207
+ 3.22e+10Hz 0.968447 -0.218869
+ 3.23e+10Hz 0.96829 -0.21953
+ 3.24e+10Hz 0.968134 -0.220191
+ 3.25e+10Hz 0.967977 -0.220852
+ 3.26e+10Hz 0.967819 -0.221513
+ 3.27e+10Hz 0.967661 -0.222173
+ 3.28e+10Hz 0.967503 -0.222834
+ 3.29e+10Hz 0.967344 -0.223494
+ 3.3e+10Hz 0.967185 -0.224154
+ 3.31e+10Hz 0.967025 -0.224814
+ 3.32e+10Hz 0.966865 -0.225474
+ 3.33e+10Hz 0.966705 -0.226134
+ 3.34e+10Hz 0.966544 -0.226794
+ 3.35e+10Hz 0.966382 -0.227453
+ 3.36e+10Hz 0.966221 -0.228113
+ 3.37e+10Hz 0.966059 -0.228772
+ 3.38e+10Hz 0.965896 -0.229431
+ 3.39e+10Hz 0.965733 -0.23009
+ 3.4e+10Hz 0.96557 -0.230749
+ 3.41e+10Hz 0.965406 -0.231407
+ 3.42e+10Hz 0.965242 -0.232066
+ 3.43e+10Hz 0.965077 -0.232725
+ 3.44e+10Hz 0.964912 -0.233383
+ 3.45e+10Hz 0.964746 -0.234041
+ 3.46e+10Hz 0.964581 -0.234699
+ 3.47e+10Hz 0.964414 -0.235357
+ 3.48e+10Hz 0.964248 -0.236015
+ 3.49e+10Hz 0.964081 -0.236673
+ 3.5e+10Hz 0.963913 -0.23733
+ 3.51e+10Hz 0.963745 -0.237987
+ 3.52e+10Hz 0.963577 -0.238645
+ 3.53e+10Hz 0.963408 -0.239302
+ 3.54e+10Hz 0.963239 -0.239959
+ 3.55e+10Hz 0.963069 -0.240616
+ 3.56e+10Hz 0.962899 -0.241273
+ 3.57e+10Hz 0.962729 -0.241929
+ 3.58e+10Hz 0.962558 -0.242586
+ 3.59e+10Hz 0.962387 -0.243242
+ 3.6e+10Hz 0.962216 -0.243899
+ 3.61e+10Hz 0.962044 -0.244555
+ 3.62e+10Hz 0.961871 -0.245211
+ 3.63e+10Hz 0.961698 -0.245867
+ 3.64e+10Hz 0.961525 -0.246523
+ 3.65e+10Hz 0.961351 -0.247179
+ 3.66e+10Hz 0.961177 -0.247834
+ 3.67e+10Hz 0.961003 -0.24849
+ 3.68e+10Hz 0.960828 -0.249145
+ 3.69e+10Hz 0.960653 -0.2498
+ 3.7e+10Hz 0.960477 -0.250455
+ 3.71e+10Hz 0.960301 -0.251111
+ 3.72e+10Hz 0.960124 -0.251765
+ 3.73e+10Hz 0.959947 -0.25242
+ 3.74e+10Hz 0.95977 -0.253075
+ 3.75e+10Hz 0.959592 -0.25373
+ 3.76e+10Hz 0.959414 -0.254384
+ 3.77e+10Hz 0.959236 -0.255039
+ 3.78e+10Hz 0.959057 -0.255693
+ 3.79e+10Hz 0.958877 -0.256347
+ 3.8e+10Hz 0.958697 -0.257001
+ 3.81e+10Hz 0.958517 -0.257655
+ 3.82e+10Hz 0.958337 -0.258309
+ 3.83e+10Hz 0.958156 -0.258963
+ 3.84e+10Hz 0.957974 -0.259616
+ 3.85e+10Hz 0.957792 -0.26027
+ 3.86e+10Hz 0.95761 -0.260923
+ 3.87e+10Hz 0.957427 -0.261577
+ 3.88e+10Hz 0.957244 -0.26223
+ 3.89e+10Hz 0.95706 -0.262883
+ 3.9e+10Hz 0.956876 -0.263536
+ 3.91e+10Hz 0.956692 -0.264189
+ 3.92e+10Hz 0.956507 -0.264842
+ 3.93e+10Hz 0.956322 -0.265494
+ 3.94e+10Hz 0.956136 -0.266147
+ 3.95e+10Hz 0.95595 -0.266799
+ 3.96e+10Hz 0.955764 -0.267452
+ 3.97e+10Hz 0.955577 -0.268104
+ 3.98e+10Hz 0.955389 -0.268756
+ 3.99e+10Hz 0.955202 -0.269408
+ 4e+10Hz 0.955013 -0.27006
+ 4.01e+10Hz 0.954825 -0.270712
+ 4.02e+10Hz 0.954636 -0.271364
+ 4.03e+10Hz 0.954446 -0.272016
+ 4.04e+10Hz 0.954256 -0.272667
+ 4.05e+10Hz 0.954066 -0.273319
+ 4.06e+10Hz 0.953875 -0.27397
+ 4.07e+10Hz 0.953684 -0.274621
+ 4.08e+10Hz 0.953492 -0.275272
+ 4.09e+10Hz 0.9533 -0.275924
+ 4.1e+10Hz 0.953107 -0.276575
+ 4.11e+10Hz 0.952914 -0.277225
+ 4.12e+10Hz 0.952721 -0.277876
+ 4.13e+10Hz 0.952527 -0.278527
+ 4.14e+10Hz 0.952333 -0.279177
+ 4.15e+10Hz 0.952138 -0.279828
+ 4.16e+10Hz 0.951943 -0.280478
+ 4.17e+10Hz 0.951748 -0.281128
+ 4.18e+10Hz 0.951552 -0.281778
+ 4.19e+10Hz 0.951355 -0.282428
+ 4.2e+10Hz 0.951158 -0.283078
+ 4.21e+10Hz 0.950961 -0.283728
+ 4.22e+10Hz 0.950763 -0.284378
+ 4.23e+10Hz 0.950565 -0.285027
+ 4.24e+10Hz 0.950366 -0.285677
+ 4.25e+10Hz 0.950167 -0.286326
+ 4.26e+10Hz 0.949967 -0.286975
+ 4.27e+10Hz 0.949767 -0.287625
+ 4.28e+10Hz 0.949567 -0.288274
+ 4.29e+10Hz 0.949366 -0.288923
+ 4.3e+10Hz 0.949165 -0.289571
+ 4.31e+10Hz 0.948963 -0.29022
+ 4.32e+10Hz 0.948761 -0.290869
+ 4.33e+10Hz 0.948558 -0.291517
+ 4.34e+10Hz 0.948355 -0.292165
+ 4.35e+10Hz 0.948151 -0.292814
+ 4.36e+10Hz 0.947947 -0.293462
+ 4.37e+10Hz 0.947743 -0.29411
+ 4.38e+10Hz 0.947538 -0.294758
+ 4.39e+10Hz 0.947332 -0.295405
+ 4.4e+10Hz 0.947126 -0.296053
+ 4.41e+10Hz 0.94692 -0.296701
+ 4.42e+10Hz 0.946713 -0.297348
+ 4.43e+10Hz 0.946506 -0.297995
+ 4.44e+10Hz 0.946299 -0.298642
+ 4.45e+10Hz 0.94609 -0.299289
+ 4.46e+10Hz 0.945882 -0.299936
+ 4.47e+10Hz 0.945673 -0.300583
+ 4.48e+10Hz 0.945463 -0.30123
+ 4.49e+10Hz 0.945253 -0.301876
+ 4.5e+10Hz 0.945043 -0.302523
+ 4.51e+10Hz 0.944832 -0.303169
+ 4.52e+10Hz 0.944621 -0.303815
+ 4.53e+10Hz 0.944409 -0.304461
+ 4.54e+10Hz 0.944196 -0.305107
+ 4.55e+10Hz 0.943984 -0.305753
+ 4.56e+10Hz 0.943771 -0.306399
+ 4.57e+10Hz 0.943557 -0.307044
+ 4.58e+10Hz 0.943343 -0.307689
+ 4.59e+10Hz 0.943128 -0.308335
+ 4.6e+10Hz 0.942913 -0.30898
+ 4.61e+10Hz 0.942698 -0.309625
+ 4.62e+10Hz 0.942482 -0.310269
+ 4.63e+10Hz 0.942266 -0.310914
+ 4.64e+10Hz 0.942049 -0.311559
+ 4.65e+10Hz 0.941831 -0.312203
+ 4.66e+10Hz 0.941614 -0.312847
+ 4.67e+10Hz 0.941395 -0.313491
+ 4.68e+10Hz 0.941177 -0.314135
+ 4.69e+10Hz 0.940958 -0.314779
+ 4.7e+10Hz 0.940738 -0.315423
+ 4.71e+10Hz 0.940518 -0.316066
+ 4.72e+10Hz 0.940297 -0.31671
+ 4.73e+10Hz 0.940076 -0.317353
+ 4.74e+10Hz 0.939855 -0.317996
+ 4.75e+10Hz 0.939633 -0.318639
+ 4.76e+10Hz 0.939411 -0.319281
+ 4.77e+10Hz 0.939188 -0.319924
+ 4.78e+10Hz 0.938964 -0.320567
+ 4.79e+10Hz 0.938741 -0.321209
+ 4.8e+10Hz 0.938516 -0.321851
+ 4.81e+10Hz 0.938292 -0.322493
+ 4.82e+10Hz 0.938067 -0.323135
+ 4.83e+10Hz 0.937841 -0.323777
+ 4.84e+10Hz 0.937615 -0.324418
+ 4.85e+10Hz 0.937389 -0.325059
+ 4.86e+10Hz 0.937162 -0.325701
+ 4.87e+10Hz 0.936934 -0.326342
+ 4.88e+10Hz 0.936706 -0.326982
+ 4.89e+10Hz 0.936478 -0.327623
+ 4.9e+10Hz 0.936249 -0.328263
+ 4.91e+10Hz 0.93602 -0.328904
+ 4.92e+10Hz 0.93579 -0.329544
+ 4.93e+10Hz 0.93556 -0.330184
+ 4.94e+10Hz 0.93533 -0.330824
+ 4.95e+10Hz 0.935099 -0.331464
+ 4.96e+10Hz 0.934867 -0.332103
+ 4.97e+10Hz 0.934635 -0.332742
+ 4.98e+10Hz 0.934403 -0.333382
+ 4.99e+10Hz 0.93417 -0.334021
+ 5e+10Hz 0.933936 -0.334659
+ 5.01e+10Hz 0.933703 -0.335298
+ 5.02e+10Hz 0.933469 -0.335937
+ 5.03e+10Hz 0.933234 -0.336575
+ 5.04e+10Hz 0.932999 -0.337213
+ 5.05e+10Hz 0.932763 -0.337851
+ 5.06e+10Hz 0.932527 -0.338489
+ 5.07e+10Hz 0.932291 -0.339126
+ 5.08e+10Hz 0.932054 -0.339764
+ 5.09e+10Hz 0.931816 -0.340401
+ 5.1e+10Hz 0.931579 -0.341038
+ 5.11e+10Hz 0.93134 -0.341675
+ 5.12e+10Hz 0.931102 -0.342311
+ 5.13e+10Hz 0.930863 -0.342948
+ 5.14e+10Hz 0.930623 -0.343584
+ 5.15e+10Hz 0.930383 -0.34422
+ 5.16e+10Hz 0.930143 -0.344856
+ 5.17e+10Hz 0.929902 -0.345492
+ 5.18e+10Hz 0.92966 -0.346128
+ 5.19e+10Hz 0.929419 -0.346763
+ 5.2e+10Hz 0.929176 -0.347398
+ 5.21e+10Hz 0.928934 -0.348033
+ 5.22e+10Hz 0.928691 -0.348668
+ 5.23e+10Hz 0.928447 -0.349303
+ 5.24e+10Hz 0.928203 -0.349937
+ 5.25e+10Hz 0.927959 -0.350571
+ 5.26e+10Hz 0.927714 -0.351206
+ 5.27e+10Hz 0.927469 -0.351839
+ 5.28e+10Hz 0.927223 -0.352473
+ 5.29e+10Hz 0.926977 -0.353107
+ 5.3e+10Hz 0.92673 -0.35374
+ 5.31e+10Hz 0.926483 -0.354373
+ 5.32e+10Hz 0.926236 -0.355006
+ 5.33e+10Hz 0.925988 -0.355639
+ 5.34e+10Hz 0.92574 -0.356271
+ 5.35e+10Hz 0.925491 -0.356904
+ 5.36e+10Hz 0.925242 -0.357536
+ 5.37e+10Hz 0.924992 -0.358168
+ 5.38e+10Hz 0.924742 -0.3588
+ 5.39e+10Hz 0.924492 -0.359431
+ 5.4e+10Hz 0.924241 -0.360063
+ 5.41e+10Hz 0.92399 -0.360694
+ 5.42e+10Hz 0.923738 -0.361325
+ 5.43e+10Hz 0.923486 -0.361956
+ 5.44e+10Hz 0.923233 -0.362586
+ 5.45e+10Hz 0.92298 -0.363217
+ 5.46e+10Hz 0.922727 -0.363847
+ 5.47e+10Hz 0.922473 -0.364477
+ 5.48e+10Hz 0.922219 -0.365107
+ 5.49e+10Hz 0.921964 -0.365737
+ 5.5e+10Hz 0.921709 -0.366366
+ 5.51e+10Hz 0.921454 -0.366995
+ 5.52e+10Hz 0.921198 -0.367625
+ 5.53e+10Hz 0.920941 -0.368253
+ 5.54e+10Hz 0.920685 -0.368882
+ 5.55e+10Hz 0.920427 -0.369511
+ 5.56e+10Hz 0.92017 -0.370139
+ 5.57e+10Hz 0.919912 -0.370767
+ 5.58e+10Hz 0.919653 -0.371395
+ 5.59e+10Hz 0.919395 -0.372023
+ 5.6e+10Hz 0.919135 -0.37265
+ 5.61e+10Hz 0.918875 -0.373278
+ 5.62e+10Hz 0.918616 -0.373905
+ 5.63e+10Hz 0.918355 -0.374532
+ 5.64e+10Hz 0.918094 -0.375159
+ 5.65e+10Hz 0.917833 -0.375785
+ 5.66e+10Hz 0.917571 -0.376412
+ 5.67e+10Hz 0.917309 -0.377038
+ 5.68e+10Hz 0.917046 -0.377664
+ 5.69e+10Hz 0.916783 -0.37829
+ 5.7e+10Hz 0.91652 -0.378915
+ 5.71e+10Hz 0.916256 -0.379541
+ 5.72e+10Hz 0.915992 -0.380166
+ 5.73e+10Hz 0.915727 -0.380791
+ 5.74e+10Hz 0.915462 -0.381416
+ 5.75e+10Hz 0.915197 -0.382041
+ 5.76e+10Hz 0.914931 -0.382665
+ 5.77e+10Hz 0.914665 -0.383289
+ 5.78e+10Hz 0.914398 -0.383913
+ 5.79e+10Hz 0.914131 -0.384537
+ 5.8e+10Hz 0.913864 -0.385161
+ 5.81e+10Hz 0.913596 -0.385785
+ 5.82e+10Hz 0.913327 -0.386408
+ 5.83e+10Hz 0.913059 -0.387031
+ 5.84e+10Hz 0.91279 -0.387654
+ 5.85e+10Hz 0.91252 -0.388277
+ 5.86e+10Hz 0.91225 -0.388899
+ 5.87e+10Hz 0.91198 -0.389522
+ 5.88e+10Hz 0.911709 -0.390144
+ 5.89e+10Hz 0.911438 -0.390766
+ 5.9e+10Hz 0.911167 -0.391388
+ 5.91e+10Hz 0.910895 -0.39201
+ 5.92e+10Hz 0.910622 -0.392631
+ 5.93e+10Hz 0.91035 -0.393252
+ 5.94e+10Hz 0.910076 -0.393873
+ 5.95e+10Hz 0.909803 -0.394494
+ 5.96e+10Hz 0.909529 -0.395115
+ 5.97e+10Hz 0.909254 -0.395736
+ 5.98e+10Hz 0.90898 -0.396356
+ 5.99e+10Hz 0.908704 -0.396976
+ 6e+10Hz 0.908429 -0.397596
+ 6.01e+10Hz 0.908153 -0.398216
+ 6.02e+10Hz 0.907876 -0.398835
+ 6.03e+10Hz 0.9076 -0.399455
+ 6.04e+10Hz 0.907322 -0.400074
+ 6.05e+10Hz 0.907045 -0.400693
+ 6.06e+10Hz 0.906767 -0.401312
+ 6.07e+10Hz 0.906488 -0.401931
+ 6.08e+10Hz 0.906209 -0.402549
+ 6.09e+10Hz 0.90593 -0.403168
+ 6.1e+10Hz 0.90565 -0.403786
+ 6.11e+10Hz 0.90537 -0.404404
+ 6.12e+10Hz 0.90509 -0.405021
+ 6.13e+10Hz 0.904809 -0.405639
+ 6.14e+10Hz 0.904528 -0.406256
+ 6.15e+10Hz 0.904246 -0.406873
+ 6.16e+10Hz 0.903964 -0.40749
+ 6.17e+10Hz 0.903681 -0.408107
+ 6.18e+10Hz 0.903398 -0.408724
+ 6.19e+10Hz 0.903115 -0.40934
+ 6.2e+10Hz 0.902831 -0.409957
+ 6.21e+10Hz 0.902547 -0.410573
+ 6.22e+10Hz 0.902262 -0.411189
+ 6.23e+10Hz 0.901977 -0.411804
+ 6.24e+10Hz 0.901692 -0.41242
+ 6.25e+10Hz 0.901406 -0.413035
+ 6.26e+10Hz 0.90112 -0.41365
+ 6.27e+10Hz 0.900833 -0.414265
+ 6.28e+10Hz 0.900546 -0.41488
+ 6.29e+10Hz 0.900259 -0.415495
+ 6.3e+10Hz 0.899971 -0.416109
+ 6.31e+10Hz 0.899683 -0.416724
+ 6.32e+10Hz 0.899394 -0.417337
+ 6.33e+10Hz 0.899105 -0.417951
+ 6.34e+10Hz 0.898815 -0.418565
+ 6.35e+10Hz 0.898525 -0.419179
+ 6.36e+10Hz 0.898235 -0.419792
+ 6.37e+10Hz 0.897944 -0.420405
+ 6.38e+10Hz 0.897653 -0.421018
+ 6.39e+10Hz 0.897362 -0.421631
+ 6.4e+10Hz 0.89707 -0.422243
+ 6.41e+10Hz 0.896777 -0.422856
+ 6.42e+10Hz 0.896484 -0.423468
+ 6.43e+10Hz 0.896191 -0.42408
+ 6.44e+10Hz 0.895897 -0.424692
+ 6.45e+10Hz 0.895603 -0.425303
+ 6.46e+10Hz 0.895309 -0.425915
+ 6.47e+10Hz 0.895014 -0.426526
+ 6.48e+10Hz 0.894718 -0.427137
+ 6.49e+10Hz 0.894423 -0.427748
+ 6.5e+10Hz 0.894127 -0.428359
+ 6.51e+10Hz 0.89383 -0.428969
+ 6.52e+10Hz 0.893533 -0.42958
+ 6.53e+10Hz 0.893235 -0.43019
+ 6.54e+10Hz 0.892938 -0.4308
+ 6.55e+10Hz 0.892639 -0.431409
+ 6.56e+10Hz 0.892341 -0.432019
+ 6.57e+10Hz 0.892042 -0.432628
+ 6.58e+10Hz 0.891742 -0.433237
+ 6.59e+10Hz 0.891442 -0.433846
+ 6.6e+10Hz 0.891142 -0.434455
+ 6.61e+10Hz 0.890841 -0.435064
+ 6.62e+10Hz 0.89054 -0.435672
+ 6.63e+10Hz 0.890238 -0.43628
+ 6.64e+10Hz 0.889936 -0.436888
+ 6.65e+10Hz 0.889633 -0.437496
+ 6.66e+10Hz 0.889331 -0.438104
+ 6.67e+10Hz 0.889027 -0.438711
+ 6.68e+10Hz 0.888723 -0.439318
+ 6.69e+10Hz 0.888419 -0.439925
+ 6.7e+10Hz 0.888115 -0.440532
+ 6.71e+10Hz 0.88781 -0.441139
+ 6.72e+10Hz 0.887504 -0.441745
+ 6.73e+10Hz 0.887198 -0.442352
+ 6.74e+10Hz 0.886892 -0.442958
+ 6.75e+10Hz 0.886585 -0.443563
+ 6.76e+10Hz 0.886278 -0.444169
+ 6.77e+10Hz 0.88597 -0.444774
+ 6.78e+10Hz 0.885662 -0.445379
+ 6.79e+10Hz 0.885354 -0.445985
+ 6.8e+10Hz 0.885045 -0.446589
+ 6.81e+10Hz 0.884736 -0.447194
+ 6.82e+10Hz 0.884426 -0.447798
+ 6.83e+10Hz 0.884116 -0.448402
+ 6.84e+10Hz 0.883805 -0.449006
+ 6.85e+10Hz 0.883494 -0.44961
+ 6.86e+10Hz 0.883183 -0.450214
+ 6.87e+10Hz 0.882871 -0.450817
+ 6.88e+10Hz 0.882559 -0.45142
+ 6.89e+10Hz 0.882246 -0.452023
+ 6.9e+10Hz 0.881933 -0.452626
+ 6.91e+10Hz 0.881619 -0.453228
+ 6.92e+10Hz 0.881305 -0.453831
+ 6.93e+10Hz 0.880991 -0.454433
+ 6.94e+10Hz 0.880676 -0.455035
+ 6.95e+10Hz 0.880361 -0.455636
+ 6.96e+10Hz 0.880045 -0.456238
+ 6.97e+10Hz 0.879729 -0.456839
+ 6.98e+10Hz 0.879412 -0.45744
+ 6.99e+10Hz 0.879095 -0.458041
+ 7e+10Hz 0.878778 -0.458641
+ 7.01e+10Hz 0.87846 -0.459242
+ 7.02e+10Hz 0.878142 -0.459842
+ 7.03e+10Hz 0.877823 -0.460442
+ 7.04e+10Hz 0.877504 -0.461041
+ 7.05e+10Hz 0.877185 -0.461641
+ 7.06e+10Hz 0.876865 -0.46224
+ 7.07e+10Hz 0.876544 -0.462839
+ 7.08e+10Hz 0.876224 -0.463438
+ 7.09e+10Hz 0.875902 -0.464036
+ 7.1e+10Hz 0.875581 -0.464635
+ 7.11e+10Hz 0.875259 -0.465233
+ 7.12e+10Hz 0.874936 -0.465831
+ 7.13e+10Hz 0.874613 -0.466428
+ 7.14e+10Hz 0.87429 -0.467026
+ 7.15e+10Hz 0.873966 -0.467623
+ 7.16e+10Hz 0.873642 -0.46822
+ 7.17e+10Hz 0.873317 -0.468817
+ 7.18e+10Hz 0.872992 -0.469413
+ 7.19e+10Hz 0.872667 -0.47001
+ 7.2e+10Hz 0.872341 -0.470606
+ 7.21e+10Hz 0.872014 -0.471201
+ 7.22e+10Hz 0.871688 -0.471797
+ 7.23e+10Hz 0.87136 -0.472392
+ 7.24e+10Hz 0.871033 -0.472987
+ 7.25e+10Hz 0.870705 -0.473582
+ 7.26e+10Hz 0.870377 -0.474177
+ 7.27e+10Hz 0.870048 -0.474771
+ 7.28e+10Hz 0.869718 -0.475365
+ 7.29e+10Hz 0.869389 -0.475959
+ 7.3e+10Hz 0.869059 -0.476553
+ 7.31e+10Hz 0.868728 -0.477147
+ 7.32e+10Hz 0.868397 -0.47774
+ 7.33e+10Hz 0.868066 -0.478333
+ 7.34e+10Hz 0.867734 -0.478926
+ 7.35e+10Hz 0.867402 -0.479518
+ 7.36e+10Hz 0.867069 -0.48011
+ 7.37e+10Hz 0.866736 -0.480702
+ 7.38e+10Hz 0.866403 -0.481294
+ 7.39e+10Hz 0.866069 -0.481886
+ 7.4e+10Hz 0.865735 -0.482477
+ 7.41e+10Hz 0.8654 -0.483068
+ 7.42e+10Hz 0.865065 -0.483659
+ 7.43e+10Hz 0.86473 -0.484249
+ 7.44e+10Hz 0.864394 -0.484839
+ 7.45e+10Hz 0.864058 -0.485429
+ 7.46e+10Hz 0.863721 -0.486019
+ 7.47e+10Hz 0.863384 -0.486609
+ 7.48e+10Hz 0.863046 -0.487198
+ 7.49e+10Hz 0.862708 -0.487787
+ 7.5e+10Hz 0.86237 -0.488376
+ 7.51e+10Hz 0.862031 -0.488965
+ 7.52e+10Hz 0.861692 -0.489553
+ 7.53e+10Hz 0.861352 -0.490141
+ 7.54e+10Hz 0.861012 -0.490729
+ 7.55e+10Hz 0.860672 -0.491316
+ 7.56e+10Hz 0.860331 -0.491903
+ 7.57e+10Hz 0.85999 -0.492491
+ 7.58e+10Hz 0.859648 -0.493077
+ 7.59e+10Hz 0.859306 -0.493664
+ 7.6e+10Hz 0.858964 -0.49425
+ 7.61e+10Hz 0.858621 -0.494836
+ 7.62e+10Hz 0.858278 -0.495422
+ 7.63e+10Hz 0.857934 -0.496008
+ 7.64e+10Hz 0.85759 -0.496593
+ 7.65e+10Hz 0.857246 -0.497178
+ 7.66e+10Hz 0.856901 -0.497763
+ 7.67e+10Hz 0.856556 -0.498347
+ 7.68e+10Hz 0.85621 -0.498932
+ 7.69e+10Hz 0.855864 -0.499516
+ 7.7e+10Hz 0.855518 -0.500099
+ 7.71e+10Hz 0.855171 -0.500683
+ 7.72e+10Hz 0.854824 -0.501266
+ 7.73e+10Hz 0.854476 -0.501849
+ 7.74e+10Hz 0.854128 -0.502432
+ 7.75e+10Hz 0.85378 -0.503014
+ 7.76e+10Hz 0.853431 -0.503597
+ 7.77e+10Hz 0.853082 -0.504178
+ 7.78e+10Hz 0.852733 -0.50476
+ 7.79e+10Hz 0.852383 -0.505342
+ 7.8e+10Hz 0.852032 -0.505923
+ 7.81e+10Hz 0.851681 -0.506504
+ 7.82e+10Hz 0.85133 -0.507085
+ 7.83e+10Hz 0.850979 -0.507665
+ 7.84e+10Hz 0.850627 -0.508245
+ 7.85e+10Hz 0.850275 -0.508825
+ 7.86e+10Hz 0.849922 -0.509405
+ 7.87e+10Hz 0.849569 -0.509984
+ 7.88e+10Hz 0.849216 -0.510563
+ 7.89e+10Hz 0.848862 -0.511142
+ 7.9e+10Hz 0.848507 -0.511721
+ 7.91e+10Hz 0.848153 -0.512299
+ 7.92e+10Hz 0.847798 -0.512878
+ 7.93e+10Hz 0.847442 -0.513455
+ 7.94e+10Hz 0.847087 -0.514033
+ 7.95e+10Hz 0.846731 -0.51461
+ 7.96e+10Hz 0.846374 -0.515188
+ 7.97e+10Hz 0.846017 -0.515764
+ 7.98e+10Hz 0.84566 -0.516341
+ 7.99e+10Hz 0.845302 -0.516917
+ 8e+10Hz 0.844944 -0.517494
+ 8.01e+10Hz 0.844586 -0.518069
+ 8.02e+10Hz 0.844227 -0.518645
+ 8.03e+10Hz 0.843868 -0.51922
+ 8.04e+10Hz 0.843508 -0.519795
+ 8.05e+10Hz 0.843148 -0.52037
+ 8.06e+10Hz 0.842788 -0.520945
+ 8.07e+10Hz 0.842427 -0.521519
+ 8.08e+10Hz 0.842066 -0.522093
+ 8.09e+10Hz 0.841704 -0.522667
+ 8.1e+10Hz 0.841342 -0.52324
+ 8.11e+10Hz 0.84098 -0.523814
+ 8.12e+10Hz 0.840618 -0.524387
+ 8.13e+10Hz 0.840255 -0.52496
+ 8.14e+10Hz 0.839891 -0.525532
+ 8.15e+10Hz 0.839527 -0.526104
+ 8.16e+10Hz 0.839163 -0.526676
+ 8.17e+10Hz 0.838799 -0.527248
+ 8.18e+10Hz 0.838434 -0.52782
+ 8.19e+10Hz 0.838069 -0.528391
+ 8.2e+10Hz 0.837703 -0.528962
+ 8.21e+10Hz 0.837337 -0.529533
+ 8.22e+10Hz 0.836971 -0.530103
+ 8.23e+10Hz 0.836604 -0.530674
+ 8.24e+10Hz 0.836237 -0.531244
+ 8.25e+10Hz 0.835869 -0.531813
+ 8.26e+10Hz 0.835501 -0.532383
+ 8.27e+10Hz 0.835133 -0.532952
+ 8.28e+10Hz 0.834764 -0.533521
+ 8.29e+10Hz 0.834395 -0.53409
+ 8.3e+10Hz 0.834026 -0.534659
+ 8.31e+10Hz 0.833656 -0.535227
+ 8.32e+10Hz 0.833286 -0.535795
+ 8.33e+10Hz 0.832916 -0.536362
+ 8.34e+10Hz 0.832545 -0.53693
+ 8.35e+10Hz 0.832173 -0.537497
+ 8.36e+10Hz 0.831802 -0.538064
+ 8.37e+10Hz 0.83143 -0.538631
+ 8.38e+10Hz 0.831057 -0.539198
+ 8.39e+10Hz 0.830685 -0.539764
+ 8.4e+10Hz 0.830311 -0.54033
+ 8.41e+10Hz 0.829938 -0.540896
+ 8.42e+10Hz 0.829564 -0.541461
+ 8.43e+10Hz 0.82919 -0.542026
+ 8.44e+10Hz 0.828815 -0.542591
+ 8.45e+10Hz 0.82844 -0.543156
+ 8.46e+10Hz 0.828064 -0.543721
+ 8.47e+10Hz 0.827689 -0.544285
+ 8.48e+10Hz 0.827313 -0.544849
+ 8.49e+10Hz 0.826936 -0.545413
+ 8.5e+10Hz 0.826559 -0.545976
+ 8.51e+10Hz 0.826182 -0.546539
+ 8.52e+10Hz 0.825804 -0.547103
+ 8.53e+10Hz 0.825426 -0.547665
+ 8.54e+10Hz 0.825048 -0.548228
+ 8.55e+10Hz 0.824669 -0.54879
+ 8.56e+10Hz 0.82429 -0.549352
+ 8.57e+10Hz 0.82391 -0.549914
+ 8.58e+10Hz 0.82353 -0.550476
+ 8.59e+10Hz 0.82315 -0.551037
+ 8.6e+10Hz 0.822769 -0.551598
+ 8.61e+10Hz 0.822388 -0.552159
+ 8.62e+10Hz 0.822007 -0.552719
+ 8.63e+10Hz 0.821625 -0.55328
+ 8.64e+10Hz 0.821243 -0.55384
+ 8.65e+10Hz 0.82086 -0.554399
+ 8.66e+10Hz 0.820477 -0.554959
+ 8.67e+10Hz 0.820094 -0.555518
+ 8.68e+10Hz 0.81971 -0.556077
+ 8.69e+10Hz 0.819326 -0.556636
+ 8.7e+10Hz 0.818942 -0.557195
+ 8.71e+10Hz 0.818557 -0.557753
+ 8.72e+10Hz 0.818172 -0.558311
+ 8.73e+10Hz 0.817786 -0.558869
+ 8.74e+10Hz 0.8174 -0.559426
+ 8.75e+10Hz 0.817013 -0.559984
+ 8.76e+10Hz 0.816627 -0.560541
+ 8.77e+10Hz 0.81624 -0.561097
+ 8.78e+10Hz 0.815852 -0.561654
+ 8.79e+10Hz 0.815464 -0.56221
+ 8.8e+10Hz 0.815076 -0.562766
+ 8.81e+10Hz 0.814687 -0.563322
+ 8.82e+10Hz 0.814298 -0.563878
+ 8.83e+10Hz 0.813909 -0.564433
+ 8.84e+10Hz 0.813519 -0.564988
+ 8.85e+10Hz 0.813129 -0.565543
+ 8.86e+10Hz 0.812738 -0.566097
+ 8.87e+10Hz 0.812347 -0.566652
+ 8.88e+10Hz 0.811956 -0.567206
+ 8.89e+10Hz 0.811564 -0.567759
+ 8.9e+10Hz 0.811172 -0.568313
+ 8.91e+10Hz 0.810779 -0.568866
+ 8.92e+10Hz 0.810387 -0.569419
+ 8.93e+10Hz 0.809993 -0.569972
+ 8.94e+10Hz 0.8096 -0.570524
+ 8.95e+10Hz 0.809206 -0.571077
+ 8.96e+10Hz 0.808811 -0.571629
+ 8.97e+10Hz 0.808416 -0.57218
+ 8.98e+10Hz 0.808021 -0.572732
+ 8.99e+10Hz 0.807625 -0.573283
+ 9e+10Hz 0.807229 -0.573834
+ 9.01e+10Hz 0.806833 -0.574385
+ 9.02e+10Hz 0.806436 -0.574935
+ 9.03e+10Hz 0.806039 -0.575485
+ 9.04e+10Hz 0.805642 -0.576035
+ 9.05e+10Hz 0.805244 -0.576585
+ 9.06e+10Hz 0.804845 -0.577134
+ 9.07e+10Hz 0.804447 -0.577683
+ 9.08e+10Hz 0.804048 -0.578232
+ 9.09e+10Hz 0.803648 -0.578781
+ 9.1e+10Hz 0.803248 -0.579329
+ 9.11e+10Hz 0.802848 -0.579877
+ 9.12e+10Hz 0.802447 -0.580425
+ 9.13e+10Hz 0.802046 -0.580973
+ 9.14e+10Hz 0.801645 -0.58152
+ 9.15e+10Hz 0.801243 -0.582067
+ 9.16e+10Hz 0.800841 -0.582614
+ 9.17e+10Hz 0.800438 -0.58316
+ 9.18e+10Hz 0.800035 -0.583706
+ 9.19e+10Hz 0.799632 -0.584252
+ 9.2e+10Hz 0.799228 -0.584798
+ 9.21e+10Hz 0.798824 -0.585343
+ 9.22e+10Hz 0.798419 -0.585889
+ 9.23e+10Hz 0.798014 -0.586433
+ 9.24e+10Hz 0.797609 -0.586978
+ 9.25e+10Hz 0.797203 -0.587522
+ 9.26e+10Hz 0.796797 -0.588066
+ 9.27e+10Hz 0.796391 -0.58861
+ 9.28e+10Hz 0.795984 -0.589153
+ 9.29e+10Hz 0.795577 -0.589697
+ 9.3e+10Hz 0.795169 -0.59024
+ 9.31e+10Hz 0.794761 -0.590782
+ 9.32e+10Hz 0.794352 -0.591325
+ 9.33e+10Hz 0.793944 -0.591867
+ 9.34e+10Hz 0.793534 -0.592409
+ 9.35e+10Hz 0.793125 -0.59295
+ 9.36e+10Hz 0.792715 -0.593491
+ 9.37e+10Hz 0.792304 -0.594032
+ 9.38e+10Hz 0.791893 -0.594573
+ 9.39e+10Hz 0.791482 -0.595113
+ 9.4e+10Hz 0.791071 -0.595653
+ 9.41e+10Hz 0.790659 -0.596193
+ 9.42e+10Hz 0.790246 -0.596733
+ 9.43e+10Hz 0.789834 -0.597272
+ 9.44e+10Hz 0.789421 -0.597811
+ 9.45e+10Hz 0.789007 -0.59835
+ 9.46e+10Hz 0.788593 -0.598888
+ 9.47e+10Hz 0.788179 -0.599426
+ 9.48e+10Hz 0.787764 -0.599964
+ 9.49e+10Hz 0.787349 -0.600502
+ 9.5e+10Hz 0.786934 -0.601039
+ 9.51e+10Hz 0.786518 -0.601576
+ 9.52e+10Hz 0.786102 -0.602112
+ 9.53e+10Hz 0.785685 -0.602649
+ 9.54e+10Hz 0.785268 -0.603185
+ 9.55e+10Hz 0.784851 -0.603721
+ 9.56e+10Hz 0.784433 -0.604256
+ 9.57e+10Hz 0.784015 -0.604791
+ 9.58e+10Hz 0.783597 -0.605326
+ 9.59e+10Hz 0.783178 -0.605861
+ 9.6e+10Hz 0.782759 -0.606395
+ 9.61e+10Hz 0.782339 -0.606929
+ 9.62e+10Hz 0.781919 -0.607463
+ 9.63e+10Hz 0.781499 -0.607996
+ 9.64e+10Hz 0.781078 -0.608529
+ 9.65e+10Hz 0.780657 -0.609062
+ 9.66e+10Hz 0.780235 -0.609595
+ 9.67e+10Hz 0.779813 -0.610127
+ 9.68e+10Hz 0.779391 -0.610659
+ 9.69e+10Hz 0.778968 -0.61119
+ 9.7e+10Hz 0.778546 -0.611721
+ 9.71e+10Hz 0.778122 -0.612252
+ 9.72e+10Hz 0.777698 -0.612783
+ 9.73e+10Hz 0.777274 -0.613313
+ 9.74e+10Hz 0.77685 -0.613843
+ 9.75e+10Hz 0.776425 -0.614373
+ 9.76e+10Hz 0.775999 -0.614903
+ 9.77e+10Hz 0.775574 -0.615432
+ 9.78e+10Hz 0.775148 -0.615961
+ 9.79e+10Hz 0.774721 -0.616489
+ 9.8e+10Hz 0.774295 -0.617017
+ 9.81e+10Hz 0.773868 -0.617545
+ 9.82e+10Hz 0.77344 -0.618073
+ 9.83e+10Hz 0.773012 -0.6186
+ 9.84e+10Hz 0.772584 -0.619127
+ 9.85e+10Hz 0.772156 -0.619654
+ 9.86e+10Hz 0.771727 -0.62018
+ 9.87e+10Hz 0.771297 -0.620706
+ 9.88e+10Hz 0.770868 -0.621232
+ 9.89e+10Hz 0.770438 -0.621757
+ 9.9e+10Hz 0.770007 -0.622282
+ 9.91e+10Hz 0.769576 -0.622807
+ 9.92e+10Hz 0.769145 -0.623332
+ 9.93e+10Hz 0.768714 -0.623856
+ 9.94e+10Hz 0.768282 -0.62438
+ 9.95e+10Hz 0.76785 -0.624903
+ 9.96e+10Hz 0.767417 -0.625426
+ 9.97e+10Hz 0.766984 -0.625949
+ 9.98e+10Hz 0.766551 -0.626472
+ 9.99e+10Hz 0.766118 -0.626994
+ 1e+11Hz 0.765684 -0.627516
+ 1.001e+11Hz 0.765249 -0.628038
+ 1.002e+11Hz 0.764815 -0.628559
+ 1.003e+11Hz 0.764379 -0.62908
+ 1.004e+11Hz 0.763944 -0.629601
+ 1.005e+11Hz 0.763508 -0.630121
+ 1.006e+11Hz 0.763072 -0.630641
+ 1.007e+11Hz 0.762636 -0.631161
+ 1.008e+11Hz 0.762199 -0.63168
+ 1.009e+11Hz 0.761762 -0.6322
+ 1.01e+11Hz 0.761324 -0.632718
+ 1.011e+11Hz 0.760887 -0.633237
+ 1.012e+11Hz 0.760448 -0.633755
+ 1.013e+11Hz 0.76001 -0.634273
+ 1.014e+11Hz 0.759571 -0.63479
+ 1.015e+11Hz 0.759132 -0.635308
+ 1.016e+11Hz 0.758692 -0.635825
+ 1.017e+11Hz 0.758252 -0.636341
+ 1.018e+11Hz 0.757812 -0.636857
+ 1.019e+11Hz 0.757372 -0.637373
+ 1.02e+11Hz 0.756931 -0.637889
+ 1.021e+11Hz 0.756489 -0.638404
+ 1.022e+11Hz 0.756048 -0.638919
+ 1.023e+11Hz 0.755606 -0.639434
+ 1.024e+11Hz 0.755164 -0.639948
+ 1.025e+11Hz 0.754721 -0.640462
+ 1.026e+11Hz 0.754278 -0.640976
+ 1.027e+11Hz 0.753835 -0.64149
+ 1.028e+11Hz 0.753391 -0.642003
+ 1.029e+11Hz 0.752947 -0.642516
+ 1.03e+11Hz 0.752503 -0.643028
+ 1.031e+11Hz 0.752058 -0.64354
+ 1.032e+11Hz 0.751613 -0.644052
+ 1.033e+11Hz 0.751168 -0.644563
+ 1.034e+11Hz 0.750722 -0.645075
+ 1.035e+11Hz 0.750276 -0.645586
+ 1.036e+11Hz 0.74983 -0.646096
+ 1.037e+11Hz 0.749383 -0.646606
+ 1.038e+11Hz 0.748937 -0.647116
+ 1.039e+11Hz 0.748489 -0.647626
+ 1.04e+11Hz 0.748042 -0.648135
+ 1.041e+11Hz 0.747594 -0.648644
+ 1.042e+11Hz 0.747146 -0.649153
+ 1.043e+11Hz 0.746697 -0.649662
+ 1.044e+11Hz 0.746248 -0.65017
+ 1.045e+11Hz 0.745799 -0.650678
+ 1.046e+11Hz 0.745349 -0.651185
+ 1.047e+11Hz 0.744899 -0.651692
+ 1.048e+11Hz 0.744449 -0.652199
+ 1.049e+11Hz 0.743998 -0.652706
+ 1.05e+11Hz 0.743548 -0.653212
+ 1.051e+11Hz 0.743096 -0.653718
+ 1.052e+11Hz 0.742645 -0.654223
+ 1.053e+11Hz 0.742193 -0.654729
+ 1.054e+11Hz 0.741741 -0.655234
+ 1.055e+11Hz 0.741288 -0.655738
+ 1.056e+11Hz 0.740835 -0.656243
+ 1.057e+11Hz 0.740382 -0.656747
+ 1.058e+11Hz 0.739929 -0.657251
+ 1.059e+11Hz 0.739475 -0.657754
+ 1.06e+11Hz 0.739021 -0.658257
+ 1.061e+11Hz 0.738566 -0.65876
+ 1.062e+11Hz 0.738112 -0.659263
+ 1.063e+11Hz 0.737657 -0.659765
+ 1.064e+11Hz 0.737201 -0.660267
+ 1.065e+11Hz 0.736745 -0.660769
+ 1.066e+11Hz 0.736289 -0.66127
+ 1.067e+11Hz 0.735833 -0.661771
+ 1.068e+11Hz 0.735376 -0.662272
+ 1.069e+11Hz 0.734919 -0.662772
+ 1.07e+11Hz 0.734462 -0.663272
+ 1.071e+11Hz 0.734004 -0.663772
+ 1.072e+11Hz 0.733546 -0.664272
+ 1.073e+11Hz 0.733088 -0.664771
+ 1.074e+11Hz 0.732629 -0.66527
+ 1.075e+11Hz 0.73217 -0.665768
+ 1.076e+11Hz 0.731711 -0.666267
+ 1.077e+11Hz 0.731251 -0.666765
+ 1.078e+11Hz 0.730791 -0.667263
+ 1.079e+11Hz 0.730331 -0.66776
+ 1.08e+11Hz 0.729871 -0.668257
+ 1.081e+11Hz 0.72941 -0.668754
+ 1.082e+11Hz 0.728948 -0.66925
+ 1.083e+11Hz 0.728487 -0.669747
+ 1.084e+11Hz 0.728025 -0.670243
+ 1.085e+11Hz 0.727563 -0.670738
+ 1.086e+11Hz 0.7271 -0.671234
+ 1.087e+11Hz 0.726637 -0.671729
+ 1.088e+11Hz 0.726174 -0.672223
+ 1.089e+11Hz 0.725711 -0.672718
+ 1.09e+11Hz 0.725247 -0.673212
+ 1.091e+11Hz 0.724783 -0.673706
+ 1.092e+11Hz 0.724318 -0.674199
+ 1.093e+11Hz 0.723853 -0.674693
+ 1.094e+11Hz 0.723388 -0.675186
+ 1.095e+11Hz 0.722923 -0.675678
+ 1.096e+11Hz 0.722457 -0.676171
+ 1.097e+11Hz 0.721991 -0.676663
+ 1.098e+11Hz 0.721525 -0.677155
+ 1.099e+11Hz 0.721058 -0.677646
+ 1.1e+11Hz 0.720591 -0.678137
+ 1.101e+11Hz 0.720123 -0.678628
+ 1.102e+11Hz 0.719655 -0.679119
+ 1.103e+11Hz 0.719187 -0.679609
+ 1.104e+11Hz 0.718719 -0.680099
+ 1.105e+11Hz 0.71825 -0.680589
+ 1.106e+11Hz 0.717781 -0.681078
+ 1.107e+11Hz 0.717312 -0.681567
+ 1.108e+11Hz 0.716842 -0.682056
+ 1.109e+11Hz 0.716372 -0.682545
+ 1.11e+11Hz 0.715901 -0.683033
+ 1.111e+11Hz 0.715431 -0.683521
+ 1.112e+11Hz 0.714959 -0.684009
+ 1.113e+11Hz 0.714488 -0.684496
+ 1.114e+11Hz 0.714016 -0.684983
+ 1.115e+11Hz 0.713544 -0.68547
+ 1.116e+11Hz 0.713072 -0.685956
+ 1.117e+11Hz 0.712599 -0.686442
+ 1.118e+11Hz 0.712126 -0.686928
+ 1.119e+11Hz 0.711653 -0.687414
+ 1.12e+11Hz 0.711179 -0.687899
+ 1.121e+11Hz 0.710705 -0.688384
+ 1.122e+11Hz 0.71023 -0.688869
+ 1.123e+11Hz 0.709755 -0.689353
+ 1.124e+11Hz 0.70928 -0.689837
+ 1.125e+11Hz 0.708805 -0.690321
+ 1.126e+11Hz 0.708329 -0.690805
+ 1.127e+11Hz 0.707853 -0.691288
+ 1.128e+11Hz 0.707376 -0.69177
+ 1.129e+11Hz 0.706899 -0.692253
+ 1.13e+11Hz 0.706422 -0.692735
+ 1.131e+11Hz 0.705945 -0.693217
+ 1.132e+11Hz 0.705467 -0.693699
+ 1.133e+11Hz 0.704989 -0.69418
+ 1.134e+11Hz 0.70451 -0.694661
+ 1.135e+11Hz 0.704031 -0.695142
+ 1.136e+11Hz 0.703552 -0.695623
+ 1.137e+11Hz 0.703072 -0.696103
+ 1.138e+11Hz 0.702592 -0.696582
+ 1.139e+11Hz 0.702112 -0.697062
+ 1.14e+11Hz 0.701631 -0.697541
+ 1.141e+11Hz 0.70115 -0.69802
+ 1.142e+11Hz 0.700669 -0.698499
+ 1.143e+11Hz 0.700187 -0.698977
+ 1.144e+11Hz 0.699705 -0.699455
+ 1.145e+11Hz 0.699223 -0.699932
+ 1.146e+11Hz 0.69874 -0.70041
+ 1.147e+11Hz 0.698257 -0.700887
+ 1.148e+11Hz 0.697774 -0.701363
+ 1.149e+11Hz 0.69729 -0.70184
+ 1.15e+11Hz 0.696806 -0.702316
+ 1.151e+11Hz 0.696322 -0.702792
+ 1.152e+11Hz 0.695837 -0.703267
+ 1.153e+11Hz 0.695352 -0.703742
+ 1.154e+11Hz 0.694866 -0.704217
+ 1.155e+11Hz 0.69438 -0.704691
+ 1.156e+11Hz 0.693894 -0.705166
+ 1.157e+11Hz 0.693407 -0.705639
+ 1.158e+11Hz 0.69292 -0.706113
+ 1.159e+11Hz 0.692433 -0.706586
+ 1.16e+11Hz 0.691945 -0.707059
+ 1.161e+11Hz 0.691458 -0.707531
+ 1.162e+11Hz 0.690969 -0.708004
+ 1.163e+11Hz 0.690481 -0.708475
+ 1.164e+11Hz 0.689992 -0.708947
+ 1.165e+11Hz 0.689502 -0.709418
+ 1.166e+11Hz 0.689013 -0.709889
+ 1.167e+11Hz 0.688522 -0.71036
+ 1.168e+11Hz 0.688032 -0.71083
+ 1.169e+11Hz 0.687541 -0.711299
+ 1.17e+11Hz 0.68705 -0.711769
+ 1.171e+11Hz 0.686559 -0.712238
+ 1.172e+11Hz 0.686067 -0.712707
+ 1.173e+11Hz 0.685575 -0.713176
+ 1.174e+11Hz 0.685082 -0.713644
+ 1.175e+11Hz 0.684589 -0.714112
+ 1.176e+11Hz 0.684096 -0.714579
+ 1.177e+11Hz 0.683602 -0.715046
+ 1.178e+11Hz 0.683109 -0.715513
+ 1.179e+11Hz 0.682614 -0.715979
+ 1.18e+11Hz 0.68212 -0.716445
+ 1.181e+11Hz 0.681625 -0.716911
+ 1.182e+11Hz 0.681129 -0.717377
+ 1.183e+11Hz 0.680634 -0.717842
+ 1.184e+11Hz 0.680138 -0.718306
+ 1.185e+11Hz 0.679641 -0.718771
+ 1.186e+11Hz 0.679145 -0.719235
+ 1.187e+11Hz 0.678648 -0.719698
+ 1.188e+11Hz 0.67815 -0.720162
+ 1.189e+11Hz 0.677652 -0.720625
+ 1.19e+11Hz 0.677154 -0.721087
+ 1.191e+11Hz 0.676656 -0.721549
+ 1.192e+11Hz 0.676157 -0.722011
+ 1.193e+11Hz 0.675658 -0.722473
+ 1.194e+11Hz 0.675159 -0.722934
+ 1.195e+11Hz 0.674659 -0.723395
+ 1.196e+11Hz 0.674159 -0.723855
+ 1.197e+11Hz 0.673658 -0.724315
+ 1.198e+11Hz 0.673158 -0.724775
+ 1.199e+11Hz 0.672656 -0.725234
+ 1.2e+11Hz 0.672155 -0.725693
+ 1.201e+11Hz 0.671653 -0.726151
+ 1.202e+11Hz 0.671151 -0.72661
+ 1.203e+11Hz 0.670649 -0.727068
+ 1.204e+11Hz 0.670146 -0.727525
+ 1.205e+11Hz 0.669643 -0.727982
+ 1.206e+11Hz 0.669139 -0.728439
+ 1.207e+11Hz 0.668636 -0.728895
+ 1.208e+11Hz 0.668131 -0.729351
+ 1.209e+11Hz 0.667627 -0.729807
+ 1.21e+11Hz 0.667122 -0.730262
+ 1.211e+11Hz 0.666617 -0.730717
+ 1.212e+11Hz 0.666112 -0.731171
+ 1.213e+11Hz 0.665606 -0.731625
+ 1.214e+11Hz 0.6651 -0.732079
+ 1.215e+11Hz 0.664593 -0.732532
+ 1.216e+11Hz 0.664087 -0.732985
+ 1.217e+11Hz 0.66358 -0.733438
+ 1.218e+11Hz 0.663072 -0.73389
+ 1.219e+11Hz 0.662565 -0.734342
+ 1.22e+11Hz 0.662057 -0.734793
+ 1.221e+11Hz 0.661549 -0.735244
+ 1.222e+11Hz 0.66104 -0.735695
+ 1.223e+11Hz 0.660531 -0.736145
+ 1.224e+11Hz 0.660022 -0.736595
+ 1.225e+11Hz 0.659512 -0.737044
+ 1.226e+11Hz 0.659003 -0.737493
+ 1.227e+11Hz 0.658492 -0.737942
+ 1.228e+11Hz 0.657982 -0.73839
+ 1.229e+11Hz 0.657471 -0.738838
+ 1.23e+11Hz 0.65696 -0.739286
+ 1.231e+11Hz 0.656449 -0.739733
+ 1.232e+11Hz 0.655937 -0.74018
+ 1.233e+11Hz 0.655425 -0.740626
+ 1.234e+11Hz 0.654913 -0.741072
+ 1.235e+11Hz 0.6544 -0.741518
+ 1.236e+11Hz 0.653887 -0.741963
+ 1.237e+11Hz 0.653374 -0.742408
+ 1.238e+11Hz 0.652861 -0.742852
+ 1.239e+11Hz 0.652347 -0.743296
+ 1.24e+11Hz 0.651833 -0.74374
+ 1.241e+11Hz 0.651319 -0.744183
+ 1.242e+11Hz 0.650804 -0.744626
+ 1.243e+11Hz 0.650289 -0.745069
+ 1.244e+11Hz 0.649774 -0.745511
+ 1.245e+11Hz 0.649259 -0.745953
+ 1.246e+11Hz 0.648743 -0.746394
+ 1.247e+11Hz 0.648227 -0.746835
+ 1.248e+11Hz 0.647711 -0.747275
+ 1.249e+11Hz 0.647194 -0.747715
+ 1.25e+11Hz 0.646677 -0.748155
+ 1.251e+11Hz 0.64616 -0.748595
+ 1.252e+11Hz 0.645643 -0.749034
+ 1.253e+11Hz 0.645125 -0.749472
+ 1.254e+11Hz 0.644607 -0.74991
+ 1.255e+11Hz 0.644089 -0.750348
+ 1.256e+11Hz 0.64357 -0.750786
+ 1.257e+11Hz 0.643052 -0.751223
+ 1.258e+11Hz 0.642533 -0.751659
+ 1.259e+11Hz 0.642013 -0.752096
+ 1.26e+11Hz 0.641494 -0.752532
+ 1.261e+11Hz 0.640974 -0.752967
+ 1.262e+11Hz 0.640454 -0.753402
+ 1.263e+11Hz 0.639933 -0.753837
+ 1.264e+11Hz 0.639413 -0.754271
+ 1.265e+11Hz 0.638892 -0.754705
+ 1.266e+11Hz 0.638371 -0.755139
+ 1.267e+11Hz 0.637849 -0.755572
+ 1.268e+11Hz 0.637328 -0.756005
+ 1.269e+11Hz 0.636806 -0.756438
+ 1.27e+11Hz 0.636284 -0.75687
+ 1.271e+11Hz 0.635761 -0.757301
+ 1.272e+11Hz 0.635239 -0.757733
+ 1.273e+11Hz 0.634716 -0.758164
+ 1.274e+11Hz 0.634192 -0.758594
+ 1.275e+11Hz 0.633669 -0.759024
+ 1.276e+11Hz 0.633145 -0.759454
+ 1.277e+11Hz 0.632621 -0.759884
+ 1.278e+11Hz 0.632097 -0.760313
+ 1.279e+11Hz 0.631573 -0.760742
+ 1.28e+11Hz 0.631048 -0.76117
+ 1.281e+11Hz 0.630523 -0.761598
+ 1.282e+11Hz 0.629998 -0.762026
+ 1.283e+11Hz 0.629472 -0.762453
+ 1.284e+11Hz 0.628947 -0.76288
+ 1.285e+11Hz 0.628421 -0.763306
+ 1.286e+11Hz 0.627895 -0.763733
+ 1.287e+11Hz 0.627368 -0.764158
+ 1.288e+11Hz 0.626842 -0.764584
+ 1.289e+11Hz 0.626315 -0.765009
+ 1.29e+11Hz 0.625787 -0.765434
+ 1.291e+11Hz 0.62526 -0.765858
+ 1.292e+11Hz 0.624732 -0.766282
+ 1.293e+11Hz 0.624205 -0.766706
+ 1.294e+11Hz 0.623676 -0.767129
+ 1.295e+11Hz 0.623148 -0.767552
+ 1.296e+11Hz 0.622619 -0.767975
+ 1.297e+11Hz 0.62209 -0.768397
+ 1.298e+11Hz 0.621561 -0.768819
+ 1.299e+11Hz 0.621032 -0.76924
+ 1.3e+11Hz 0.620502 -0.769661
+ 1.301e+11Hz 0.619973 -0.770082
+ 1.302e+11Hz 0.619443 -0.770503
+ 1.303e+11Hz 0.618912 -0.770923
+ 1.304e+11Hz 0.618382 -0.771343
+ 1.305e+11Hz 0.617851 -0.771762
+ 1.306e+11Hz 0.61732 -0.772181
+ 1.307e+11Hz 0.616788 -0.7726
+ 1.308e+11Hz 0.616257 -0.773019
+ 1.309e+11Hz 0.615725 -0.773437
+ 1.31e+11Hz 0.615193 -0.773855
+ 1.311e+11Hz 0.614661 -0.774272
+ 1.312e+11Hz 0.614128 -0.774689
+ 1.313e+11Hz 0.613595 -0.775106
+ 1.314e+11Hz 0.613062 -0.775522
+ 1.315e+11Hz 0.612529 -0.775938
+ 1.316e+11Hz 0.611996 -0.776354
+ 1.317e+11Hz 0.611462 -0.77677
+ 1.318e+11Hz 0.610928 -0.777185
+ 1.319e+11Hz 0.610394 -0.7776
+ 1.32e+11Hz 0.609859 -0.778014
+ 1.321e+11Hz 0.609324 -0.778428
+ 1.322e+11Hz 0.608789 -0.778842
+ 1.323e+11Hz 0.608254 -0.779255
+ 1.324e+11Hz 0.607718 -0.779669
+ 1.325e+11Hz 0.607182 -0.780081
+ 1.326e+11Hz 0.606646 -0.780494
+ 1.327e+11Hz 0.60611 -0.780906
+ 1.328e+11Hz 0.605573 -0.781318
+ 1.329e+11Hz 0.605037 -0.78173
+ 1.33e+11Hz 0.6045 -0.782141
+ 1.331e+11Hz 0.603962 -0.782552
+ 1.332e+11Hz 0.603425 -0.782962
+ 1.333e+11Hz 0.602887 -0.783373
+ 1.334e+11Hz 0.602348 -0.783783
+ 1.335e+11Hz 0.60181 -0.784192
+ 1.336e+11Hz 0.601271 -0.784602
+ 1.337e+11Hz 0.600732 -0.785011
+ 1.338e+11Hz 0.600193 -0.785419
+ 1.339e+11Hz 0.599654 -0.785828
+ 1.34e+11Hz 0.599114 -0.786236
+ 1.341e+11Hz 0.598574 -0.786644
+ 1.342e+11Hz 0.598033 -0.787051
+ 1.343e+11Hz 0.597493 -0.787458
+ 1.344e+11Hz 0.596952 -0.787865
+ 1.345e+11Hz 0.596411 -0.788271
+ 1.346e+11Hz 0.595869 -0.788678
+ 1.347e+11Hz 0.595327 -0.789083
+ 1.348e+11Hz 0.594785 -0.789489
+ 1.349e+11Hz 0.594243 -0.789894
+ 1.35e+11Hz 0.5937 -0.790299
+ 1.351e+11Hz 0.593158 -0.790704
+ 1.352e+11Hz 0.592614 -0.791108
+ 1.353e+11Hz 0.592071 -0.791512
+ 1.354e+11Hz 0.591527 -0.791915
+ 1.355e+11Hz 0.590983 -0.792319
+ 1.356e+11Hz 0.590438 -0.792722
+ 1.357e+11Hz 0.589894 -0.793125
+ 1.358e+11Hz 0.589349 -0.793527
+ 1.359e+11Hz 0.588804 -0.793929
+ 1.36e+11Hz 0.588258 -0.794331
+ 1.361e+11Hz 0.587712 -0.794732
+ 1.362e+11Hz 0.587166 -0.795133
+ 1.363e+11Hz 0.586619 -0.795534
+ 1.364e+11Hz 0.586072 -0.795934
+ 1.365e+11Hz 0.585525 -0.796334
+ 1.366e+11Hz 0.584978 -0.796734
+ 1.367e+11Hz 0.58443 -0.797134
+ 1.368e+11Hz 0.583882 -0.797533
+ 1.369e+11Hz 0.583333 -0.797932
+ 1.37e+11Hz 0.582785 -0.79833
+ 1.371e+11Hz 0.582236 -0.798728
+ 1.372e+11Hz 0.581686 -0.799126
+ 1.373e+11Hz 0.581137 -0.799524
+ 1.374e+11Hz 0.580587 -0.799921
+ 1.375e+11Hz 0.580036 -0.800318
+ 1.376e+11Hz 0.579485 -0.800714
+ 1.377e+11Hz 0.578935 -0.80111
+ 1.378e+11Hz 0.578383 -0.801506
+ 1.379e+11Hz 0.577832 -0.801902
+ 1.38e+11Hz 0.577279 -0.802297
+ 1.381e+11Hz 0.576727 -0.802692
+ 1.382e+11Hz 0.576174 -0.803086
+ 1.383e+11Hz 0.575621 -0.80348
+ 1.384e+11Hz 0.575068 -0.803874
+ 1.385e+11Hz 0.574514 -0.804267
+ 1.386e+11Hz 0.57396 -0.80466
+ 1.387e+11Hz 0.573406 -0.805053
+ 1.388e+11Hz 0.572851 -0.805445
+ 1.389e+11Hz 0.572296 -0.805837
+ 1.39e+11Hz 0.571741 -0.806229
+ 1.391e+11Hz 0.571185 -0.80662
+ 1.392e+11Hz 0.570629 -0.807011
+ 1.393e+11Hz 0.570072 -0.807402
+ 1.394e+11Hz 0.569516 -0.807792
+ 1.395e+11Hz 0.568958 -0.808182
+ 1.396e+11Hz 0.568401 -0.808571
+ 1.397e+11Hz 0.567843 -0.80896
+ 1.398e+11Hz 0.567285 -0.809349
+ 1.399e+11Hz 0.566726 -0.809737
+ 1.4e+11Hz 0.566167 -0.810125
+ 1.401e+11Hz 0.565608 -0.810512
+ 1.402e+11Hz 0.565049 -0.810899
+ 1.403e+11Hz 0.564489 -0.811286
+ 1.404e+11Hz 0.563928 -0.811673
+ 1.405e+11Hz 0.563368 -0.812059
+ 1.406e+11Hz 0.562807 -0.812444
+ 1.407e+11Hz 0.562245 -0.812829
+ 1.408e+11Hz 0.561684 -0.813214
+ 1.409e+11Hz 0.561122 -0.813598
+ 1.41e+11Hz 0.560559 -0.813982
+ 1.411e+11Hz 0.559996 -0.814366
+ 1.412e+11Hz 0.559433 -0.814749
+ 1.413e+11Hz 0.55887 -0.815132
+ 1.414e+11Hz 0.558306 -0.815514
+ 1.415e+11Hz 0.557742 -0.815896
+ 1.416e+11Hz 0.557177 -0.816277
+ 1.417e+11Hz 0.556612 -0.816658
+ 1.418e+11Hz 0.556047 -0.817039
+ 1.419e+11Hz 0.555481 -0.817419
+ 1.42e+11Hz 0.554916 -0.817799
+ 1.421e+11Hz 0.554349 -0.818178
+ 1.422e+11Hz 0.553783 -0.818557
+ 1.423e+11Hz 0.553216 -0.818936
+ 1.424e+11Hz 0.552648 -0.819314
+ 1.425e+11Hz 0.552081 -0.819691
+ 1.426e+11Hz 0.551513 -0.820068
+ 1.427e+11Hz 0.550944 -0.820445
+ 1.428e+11Hz 0.550376 -0.820821
+ 1.429e+11Hz 0.549807 -0.821197
+ 1.43e+11Hz 0.549237 -0.821572
+ 1.431e+11Hz 0.548668 -0.821947
+ 1.432e+11Hz 0.548098 -0.822321
+ 1.433e+11Hz 0.547527 -0.822695
+ 1.434e+11Hz 0.546957 -0.823069
+ 1.435e+11Hz 0.546386 -0.823442
+ 1.436e+11Hz 0.545814 -0.823814
+ 1.437e+11Hz 0.545243 -0.824186
+ 1.438e+11Hz 0.544671 -0.824558
+ 1.439e+11Hz 0.544099 -0.824929
+ 1.44e+11Hz 0.543526 -0.825299
+ 1.441e+11Hz 0.542953 -0.825669
+ 1.442e+11Hz 0.54238 -0.826039
+ 1.443e+11Hz 0.541806 -0.826408
+ 1.444e+11Hz 0.541232 -0.826777
+ 1.445e+11Hz 0.540658 -0.827145
+ 1.446e+11Hz 0.540084 -0.827513
+ 1.447e+11Hz 0.539509 -0.82788
+ 1.448e+11Hz 0.538934 -0.828247
+ 1.449e+11Hz 0.538359 -0.828613
+ 1.45e+11Hz 0.537783 -0.828979
+ 1.451e+11Hz 0.537207 -0.829344
+ 1.452e+11Hz 0.536631 -0.829708
+ 1.453e+11Hz 0.536054 -0.830073
+ 1.454e+11Hz 0.535478 -0.830436
+ 1.455e+11Hz 0.534901 -0.8308
+ 1.456e+11Hz 0.534323 -0.831162
+ 1.457e+11Hz 0.533746 -0.831524
+ 1.458e+11Hz 0.533168 -0.831886
+ 1.459e+11Hz 0.53259 -0.832247
+ 1.46e+11Hz 0.532011 -0.832608
+ 1.461e+11Hz 0.531432 -0.832968
+ 1.462e+11Hz 0.530853 -0.833328
+ 1.463e+11Hz 0.530274 -0.833687
+ 1.464e+11Hz 0.529695 -0.834046
+ 1.465e+11Hz 0.529115 -0.834404
+ 1.466e+11Hz 0.528535 -0.834761
+ 1.467e+11Hz 0.527955 -0.835118
+ 1.468e+11Hz 0.527375 -0.835475
+ 1.469e+11Hz 0.526794 -0.835831
+ 1.47e+11Hz 0.526213 -0.836187
+ 1.471e+11Hz 0.525632 -0.836542
+ 1.472e+11Hz 0.525051 -0.836896
+ 1.473e+11Hz 0.524469 -0.83725
+ 1.474e+11Hz 0.523887 -0.837604
+ 1.475e+11Hz 0.523306 -0.837957
+ 1.476e+11Hz 0.522723 -0.838309
+ 1.477e+11Hz 0.522141 -0.838661
+ 1.478e+11Hz 0.521558 -0.839012
+ 1.479e+11Hz 0.520976 -0.839363
+ 1.48e+11Hz 0.520393 -0.839714
+ 1.481e+11Hz 0.51981 -0.840064
+ 1.482e+11Hz 0.519226 -0.840413
+ 1.483e+11Hz 0.518643 -0.840762
+ 1.484e+11Hz 0.518059 -0.84111
+ 1.485e+11Hz 0.517475 -0.841458
+ 1.486e+11Hz 0.516891 -0.841806
+ 1.487e+11Hz 0.516307 -0.842153
+ 1.488e+11Hz 0.515722 -0.842499
+ 1.489e+11Hz 0.515138 -0.842845
+ 1.49e+11Hz 0.514553 -0.84319
+ 1.491e+11Hz 0.513968 -0.843535
+ 1.492e+11Hz 0.513383 -0.84388
+ 1.493e+11Hz 0.512798 -0.844224
+ 1.494e+11Hz 0.512212 -0.844567
+ 1.495e+11Hz 0.511627 -0.84491
+ 1.496e+11Hz 0.511041 -0.845253
+ 1.497e+11Hz 0.510455 -0.845595
+ 1.498e+11Hz 0.509869 -0.845936
+ 1.499e+11Hz 0.509283 -0.846277
+ 1.5e+11Hz 0.508697 -0.846618
+ ]

A21 %vd(10 3) %vd(21, 22) xfer3
.model xfer3 xfer R_I=true table=[
+ 0Hz 0.996076 0
+ 1e+08Hz 0.996075 -0.000713666
+ 2e+08Hz 0.996074 -0.00142732
+ 3e+08Hz 0.996071 -0.00214095
+ 4e+08Hz 0.996068 -0.00285455
+ 5e+08Hz 0.996064 -0.0035681
+ 6e+08Hz 0.996058 -0.0042816
+ 7e+08Hz 0.996052 -0.00499503
+ 8e+08Hz 0.996045 -0.00570838
+ 9e+08Hz 0.996036 -0.00642164
+ 1e+09Hz 0.996027 -0.0071348
+ 1.1e+09Hz 0.996017 -0.00784785
+ 1.2e+09Hz 0.996006 -0.00856077
+ 1.3e+09Hz 0.995994 -0.00927357
+ 1.4e+09Hz 0.995981 -0.00998621
+ 1.5e+09Hz 0.995967 -0.0106987
+ 1.6e+09Hz 0.995952 -0.011411
+ 1.7e+09Hz 0.995936 -0.0121232
+ 1.8e+09Hz 0.995919 -0.0128352
+ 1.9e+09Hz 0.995901 -0.0135469
+ 2e+09Hz 0.995882 -0.0142585
+ 2.1e+09Hz 0.995863 -0.0149698
+ 2.2e+09Hz 0.995842 -0.015681
+ 2.3e+09Hz 0.995821 -0.0163918
+ 2.4e+09Hz 0.995798 -0.0171025
+ 2.5e+09Hz 0.995775 -0.0178129
+ 2.6e+09Hz 0.995751 -0.018523
+ 2.7e+09Hz 0.995726 -0.0192329
+ 2.8e+09Hz 0.9957 -0.0199424
+ 2.9e+09Hz 0.995673 -0.0206517
+ 3e+09Hz 0.995646 -0.0213607
+ 3.1e+09Hz 0.995617 -0.0220694
+ 3.2e+09Hz 0.995588 -0.0227777
+ 3.3e+09Hz 0.995557 -0.0234858
+ 3.4e+09Hz 0.995526 -0.0241935
+ 3.5e+09Hz 0.995494 -0.0249009
+ 3.6e+09Hz 0.995462 -0.0256079
+ 3.7e+09Hz 0.995428 -0.0263146
+ 3.8e+09Hz 0.995394 -0.0270209
+ 3.9e+09Hz 0.995359 -0.0277269
+ 4e+09Hz 0.995323 -0.0284325
+ 4.1e+09Hz 0.995286 -0.0291377
+ 4.2e+09Hz 0.995248 -0.0298426
+ 4.3e+09Hz 0.99521 -0.030547
+ 4.4e+09Hz 0.995171 -0.0312511
+ 4.5e+09Hz 0.995131 -0.0319547
+ 4.6e+09Hz 0.995091 -0.032658
+ 4.7e+09Hz 0.99505 -0.0333609
+ 4.8e+09Hz 0.995008 -0.0340633
+ 4.9e+09Hz 0.994965 -0.0347653
+ 5e+09Hz 0.994922 -0.0354669
+ 5.1e+09Hz 0.994878 -0.0361681
+ 5.2e+09Hz 0.994833 -0.0368689
+ 5.3e+09Hz 0.994788 -0.0375692
+ 5.4e+09Hz 0.994742 -0.0382691
+ 5.5e+09Hz 0.994695 -0.0389686
+ 5.6e+09Hz 0.994648 -0.0396676
+ 5.7e+09Hz 0.994599 -0.0403662
+ 5.8e+09Hz 0.994551 -0.0410643
+ 5.9e+09Hz 0.994502 -0.041762
+ 6e+09Hz 0.994452 -0.0424593
+ 6.1e+09Hz 0.994401 -0.0431561
+ 6.2e+09Hz 0.99435 -0.0438525
+ 6.3e+09Hz 0.994299 -0.0445484
+ 6.4e+09Hz 0.994247 -0.0452439
+ 6.5e+09Hz 0.994194 -0.0459389
+ 6.6e+09Hz 0.99414 -0.0466335
+ 6.7e+09Hz 0.994087 -0.0473276
+ 6.8e+09Hz 0.994032 -0.0480213
+ 6.9e+09Hz 0.993977 -0.0487146
+ 7e+09Hz 0.993922 -0.0494074
+ 7.1e+09Hz 0.993866 -0.0500997
+ 7.2e+09Hz 0.99381 -0.0507916
+ 7.3e+09Hz 0.993753 -0.0514831
+ 7.4e+09Hz 0.993695 -0.0521741
+ 7.5e+09Hz 0.993638 -0.0528647
+ 7.6e+09Hz 0.993579 -0.0535549
+ 7.7e+09Hz 0.993521 -0.0542446
+ 7.8e+09Hz 0.993461 -0.0549339
+ 7.9e+09Hz 0.993402 -0.0556228
+ 8e+09Hz 0.993342 -0.0563113
+ 8.1e+09Hz 0.993281 -0.0569993
+ 8.2e+09Hz 0.99322 -0.0576869
+ 8.3e+09Hz 0.993159 -0.0583741
+ 8.4e+09Hz 0.993097 -0.0590609
+ 8.5e+09Hz 0.993035 -0.0597473
+ 8.6e+09Hz 0.992973 -0.0604333
+ 8.7e+09Hz 0.99291 -0.0611188
+ 8.8e+09Hz 0.992847 -0.061804
+ 8.9e+09Hz 0.992783 -0.0624888
+ 9e+09Hz 0.992719 -0.0631732
+ 9.1e+09Hz 0.992655 -0.0638573
+ 9.2e+09Hz 0.99259 -0.0645409
+ 9.3e+09Hz 0.992525 -0.0652242
+ 9.4e+09Hz 0.99246 -0.0659071
+ 9.5e+09Hz 0.992394 -0.0665897
+ 9.6e+09Hz 0.992328 -0.0672719
+ 9.7e+09Hz 0.992262 -0.0679537
+ 9.8e+09Hz 0.992195 -0.0686352
+ 9.9e+09Hz 0.992128 -0.0693164
+ 1e+10Hz 0.992061 -0.0699972
+ 1.01e+10Hz 0.991994 -0.0706777
+ 1.02e+10Hz 0.991926 -0.0713579
+ 1.03e+10Hz 0.991858 -0.0720378
+ 1.04e+10Hz 0.99179 -0.0727174
+ 1.05e+10Hz 0.991721 -0.0733966
+ 1.06e+10Hz 0.991652 -0.0740756
+ 1.07e+10Hz 0.991583 -0.0747542
+ 1.08e+10Hz 0.991514 -0.0754326
+ 1.09e+10Hz 0.991444 -0.0761107
+ 1.1e+10Hz 0.991374 -0.0767885
+ 1.11e+10Hz 0.991304 -0.0774661
+ 1.12e+10Hz 0.991233 -0.0781434
+ 1.13e+10Hz 0.991162 -0.0788204
+ 1.14e+10Hz 0.991091 -0.0794972
+ 1.15e+10Hz 0.99102 -0.0801738
+ 1.16e+10Hz 0.990949 -0.0808501
+ 1.17e+10Hz 0.990877 -0.0815261
+ 1.18e+10Hz 0.990805 -0.082202
+ 1.19e+10Hz 0.990733 -0.0828776
+ 1.2e+10Hz 0.99066 -0.0835531
+ 1.21e+10Hz 0.990587 -0.0842283
+ 1.22e+10Hz 0.990514 -0.0849033
+ 1.23e+10Hz 0.990441 -0.0855781
+ 1.24e+10Hz 0.990368 -0.0862528
+ 1.25e+10Hz 0.990294 -0.0869272
+ 1.26e+10Hz 0.99022 -0.0876015
+ 1.27e+10Hz 0.990146 -0.0882757
+ 1.28e+10Hz 0.990072 -0.0889496
+ 1.29e+10Hz 0.989997 -0.0896234
+ 1.3e+10Hz 0.989922 -0.0902971
+ 1.31e+10Hz 0.989847 -0.0909706
+ 1.32e+10Hz 0.989772 -0.0916439
+ 1.33e+10Hz 0.989696 -0.0923172
+ 1.34e+10Hz 0.98962 -0.0929903
+ 1.35e+10Hz 0.989544 -0.0936633
+ 1.36e+10Hz 0.989468 -0.0943361
+ 1.37e+10Hz 0.989392 -0.0950089
+ 1.38e+10Hz 0.989315 -0.0956815
+ 1.39e+10Hz 0.989238 -0.0963541
+ 1.4e+10Hz 0.98916 -0.0970265
+ 1.41e+10Hz 0.989083 -0.0976989
+ 1.42e+10Hz 0.989005 -0.0983712
+ 1.43e+10Hz 0.988927 -0.0990434
+ 1.44e+10Hz 0.988849 -0.0997155
+ 1.45e+10Hz 0.98877 -0.100388
+ 1.46e+10Hz 0.988691 -0.101059
+ 1.47e+10Hz 0.988612 -0.101732
+ 1.48e+10Hz 0.988533 -0.102403
+ 1.49e+10Hz 0.988453 -0.103075
+ 1.5e+10Hz 0.988374 -0.103747
+ 1.51e+10Hz 0.988293 -0.104419
+ 1.52e+10Hz 0.988213 -0.10509
+ 1.53e+10Hz 0.988132 -0.105762
+ 1.54e+10Hz 0.988051 -0.106434
+ 1.55e+10Hz 0.98797 -0.107105
+ 1.56e+10Hz 0.987888 -0.107777
+ 1.57e+10Hz 0.987807 -0.108448
+ 1.58e+10Hz 0.987724 -0.10912
+ 1.59e+10Hz 0.987642 -0.109791
+ 1.6e+10Hz 0.987559 -0.110463
+ 1.61e+10Hz 0.987476 -0.111134
+ 1.62e+10Hz 0.987393 -0.111806
+ 1.63e+10Hz 0.987309 -0.112477
+ 1.64e+10Hz 0.987225 -0.113148
+ 1.65e+10Hz 0.987141 -0.11382
+ 1.66e+10Hz 0.987056 -0.114491
+ 1.67e+10Hz 0.986971 -0.115163
+ 1.68e+10Hz 0.986886 -0.115834
+ 1.69e+10Hz 0.9868 -0.116506
+ 1.7e+10Hz 0.986714 -0.117177
+ 1.71e+10Hz 0.986628 -0.117849
+ 1.72e+10Hz 0.986541 -0.11852
+ 1.73e+10Hz 0.986454 -0.119192
+ 1.74e+10Hz 0.986367 -0.119863
+ 1.75e+10Hz 0.986279 -0.120535
+ 1.76e+10Hz 0.986191 -0.121206
+ 1.77e+10Hz 0.986103 -0.121878
+ 1.78e+10Hz 0.986014 -0.12255
+ 1.79e+10Hz 0.985925 -0.123221
+ 1.8e+10Hz 0.985835 -0.123893
+ 1.81e+10Hz 0.985745 -0.124565
+ 1.82e+10Hz 0.985655 -0.125236
+ 1.83e+10Hz 0.985564 -0.125908
+ 1.84e+10Hz 0.985473 -0.12658
+ 1.85e+10Hz 0.985382 -0.127252
+ 1.86e+10Hz 0.98529 -0.127923
+ 1.87e+10Hz 0.985198 -0.128595
+ 1.88e+10Hz 0.985105 -0.129267
+ 1.89e+10Hz 0.985012 -0.129939
+ 1.9e+10Hz 0.984918 -0.130611
+ 1.91e+10Hz 0.984824 -0.131283
+ 1.92e+10Hz 0.98473 -0.131955
+ 1.93e+10Hz 0.984635 -0.132627
+ 1.94e+10Hz 0.98454 -0.133299
+ 1.95e+10Hz 0.984444 -0.133971
+ 1.96e+10Hz 0.984348 -0.134643
+ 1.97e+10Hz 0.984252 -0.135315
+ 1.98e+10Hz 0.984155 -0.135987
+ 1.99e+10Hz 0.984058 -0.136659
+ 2e+10Hz 0.98396 -0.137331
+ 2.01e+10Hz 0.983862 -0.138004
+ 2.02e+10Hz 0.983763 -0.138676
+ 2.03e+10Hz 0.983664 -0.139348
+ 2.04e+10Hz 0.983564 -0.14002
+ 2.05e+10Hz 0.983464 -0.140692
+ 2.06e+10Hz 0.983364 -0.141365
+ 2.07e+10Hz 0.983263 -0.142037
+ 2.08e+10Hz 0.983161 -0.142709
+ 2.09e+10Hz 0.983059 -0.143381
+ 2.1e+10Hz 0.982957 -0.144054
+ 2.11e+10Hz 0.982854 -0.144726
+ 2.12e+10Hz 0.982751 -0.145398
+ 2.13e+10Hz 0.982647 -0.14607
+ 2.14e+10Hz 0.982542 -0.146742
+ 2.15e+10Hz 0.982438 -0.147415
+ 2.16e+10Hz 0.982332 -0.148087
+ 2.17e+10Hz 0.982227 -0.148759
+ 2.18e+10Hz 0.98212 -0.149431
+ 2.19e+10Hz 0.982014 -0.150104
+ 2.2e+10Hz 0.981907 -0.150776
+ 2.21e+10Hz 0.981799 -0.151448
+ 2.22e+10Hz 0.981691 -0.15212
+ 2.23e+10Hz 0.981582 -0.152792
+ 2.24e+10Hz 0.981473 -0.153464
+ 2.25e+10Hz 0.981363 -0.154136
+ 2.26e+10Hz 0.981253 -0.154808
+ 2.27e+10Hz 0.981142 -0.15548
+ 2.28e+10Hz 0.981031 -0.156152
+ 2.29e+10Hz 0.980919 -0.156824
+ 2.3e+10Hz 0.980807 -0.157496
+ 2.31e+10Hz 0.980694 -0.158168
+ 2.32e+10Hz 0.980581 -0.158839
+ 2.33e+10Hz 0.980467 -0.159511
+ 2.34e+10Hz 0.980353 -0.160183
+ 2.35e+10Hz 0.980238 -0.160855
+ 2.36e+10Hz 0.980123 -0.161526
+ 2.37e+10Hz 0.980007 -0.162198
+ 2.38e+10Hz 0.979891 -0.162869
+ 2.39e+10Hz 0.979774 -0.163541
+ 2.4e+10Hz 0.979657 -0.164212
+ 2.41e+10Hz 0.979539 -0.164883
+ 2.42e+10Hz 0.979421 -0.165554
+ 2.43e+10Hz 0.979302 -0.166225
+ 2.44e+10Hz 0.979182 -0.166897
+ 2.45e+10Hz 0.979062 -0.167568
+ 2.46e+10Hz 0.978942 -0.168238
+ 2.47e+10Hz 0.978821 -0.168909
+ 2.48e+10Hz 0.9787 -0.16958
+ 2.49e+10Hz 0.978578 -0.170251
+ 2.5e+10Hz 0.978456 -0.170921
+ 2.51e+10Hz 0.978333 -0.171592
+ 2.52e+10Hz 0.978209 -0.172262
+ 2.53e+10Hz 0.978085 -0.172932
+ 2.54e+10Hz 0.977961 -0.173603
+ 2.55e+10Hz 0.977836 -0.174273
+ 2.56e+10Hz 0.97771 -0.174943
+ 2.57e+10Hz 0.977584 -0.175613
+ 2.58e+10Hz 0.977458 -0.176283
+ 2.59e+10Hz 0.977331 -0.176952
+ 2.6e+10Hz 0.977204 -0.177622
+ 2.61e+10Hz 0.977075 -0.178291
+ 2.62e+10Hz 0.976947 -0.178961
+ 2.63e+10Hz 0.976818 -0.17963
+ 2.64e+10Hz 0.976689 -0.180299
+ 2.65e+10Hz 0.976559 -0.180968
+ 2.66e+10Hz 0.976428 -0.181637
+ 2.67e+10Hz 0.976297 -0.182306
+ 2.68e+10Hz 0.976166 -0.182975
+ 2.69e+10Hz 0.976034 -0.183643
+ 2.7e+10Hz 0.975901 -0.184311
+ 2.71e+10Hz 0.975768 -0.18498
+ 2.72e+10Hz 0.975635 -0.185648
+ 2.73e+10Hz 0.975501 -0.186316
+ 2.74e+10Hz 0.975367 -0.186984
+ 2.75e+10Hz 0.975232 -0.187652
+ 2.76e+10Hz 0.975096 -0.188319
+ 2.77e+10Hz 0.97496 -0.188987
+ 2.78e+10Hz 0.974824 -0.189654
+ 2.79e+10Hz 0.974687 -0.190322
+ 2.8e+10Hz 0.97455 -0.190989
+ 2.81e+10Hz 0.974412 -0.191656
+ 2.82e+10Hz 0.974274 -0.192323
+ 2.83e+10Hz 0.974135 -0.192989
+ 2.84e+10Hz 0.973996 -0.193656
+ 2.85e+10Hz 0.973856 -0.194322
+ 2.86e+10Hz 0.973716 -0.194989
+ 2.87e+10Hz 0.973575 -0.195655
+ 2.88e+10Hz 0.973434 -0.196321
+ 2.89e+10Hz 0.973292 -0.196987
+ 2.9e+10Hz 0.97315 -0.197652
+ 2.91e+10Hz 0.973008 -0.198318
+ 2.92e+10Hz 0.972865 -0.198983
+ 2.93e+10Hz 0.972722 -0.199649
+ 2.94e+10Hz 0.972578 -0.200314
+ 2.95e+10Hz 0.972433 -0.200979
+ 2.96e+10Hz 0.972288 -0.201644
+ 2.97e+10Hz 0.972143 -0.202308
+ 2.98e+10Hz 0.971997 -0.202973
+ 2.99e+10Hz 0.971851 -0.203637
+ 3e+10Hz 0.971705 -0.204301
+ 3.01e+10Hz 0.971558 -0.204966
+ 3.02e+10Hz 0.97141 -0.205629
+ 3.03e+10Hz 0.971262 -0.206293
+ 3.04e+10Hz 0.971114 -0.206957
+ 3.05e+10Hz 0.970965 -0.207621
+ 3.06e+10Hz 0.970816 -0.208284
+ 3.07e+10Hz 0.970666 -0.208947
+ 3.08e+10Hz 0.970516 -0.20961
+ 3.09e+10Hz 0.970365 -0.210273
+ 3.1e+10Hz 0.970214 -0.210936
+ 3.11e+10Hz 0.970063 -0.211598
+ 3.12e+10Hz 0.969911 -0.212261
+ 3.13e+10Hz 0.969758 -0.212923
+ 3.14e+10Hz 0.969606 -0.213586
+ 3.15e+10Hz 0.969452 -0.214248
+ 3.16e+10Hz 0.969299 -0.21491
+ 3.17e+10Hz 0.969145 -0.215571
+ 3.18e+10Hz 0.96899 -0.216233
+ 3.19e+10Hz 0.968835 -0.216894
+ 3.2e+10Hz 0.96868 -0.217556
+ 3.21e+10Hz 0.968524 -0.218217
+ 3.22e+10Hz 0.968368 -0.218878
+ 3.23e+10Hz 0.968211 -0.219539
+ 3.24e+10Hz 0.968054 -0.2202
+ 3.25e+10Hz 0.967897 -0.22086
+ 3.26e+10Hz 0.967739 -0.221521
+ 3.27e+10Hz 0.967581 -0.222181
+ 3.28e+10Hz 0.967422 -0.222841
+ 3.29e+10Hz 0.967263 -0.223501
+ 3.3e+10Hz 0.967103 -0.224161
+ 3.31e+10Hz 0.966943 -0.224821
+ 3.32e+10Hz 0.966783 -0.225481
+ 3.33e+10Hz 0.966622 -0.22614
+ 3.34e+10Hz 0.966461 -0.2268
+ 3.35e+10Hz 0.966299 -0.227459
+ 3.36e+10Hz 0.966137 -0.228118
+ 3.37e+10Hz 0.965975 -0.228777
+ 3.38e+10Hz 0.965812 -0.229436
+ 3.39e+10Hz 0.965649 -0.230095
+ 3.4e+10Hz 0.965485 -0.230753
+ 3.41e+10Hz 0.965321 -0.231412
+ 3.42e+10Hz 0.965156 -0.23207
+ 3.43e+10Hz 0.964991 -0.232729
+ 3.44e+10Hz 0.964826 -0.233387
+ 3.45e+10Hz 0.96466 -0.234045
+ 3.46e+10Hz 0.964494 -0.234702
+ 3.47e+10Hz 0.964328 -0.23536
+ 3.48e+10Hz 0.964161 -0.236018
+ 3.49e+10Hz 0.963993 -0.236675
+ 3.5e+10Hz 0.963826 -0.237333
+ 3.51e+10Hz 0.963657 -0.23799
+ 3.52e+10Hz 0.963489 -0.238647
+ 3.53e+10Hz 0.96332 -0.239304
+ 3.54e+10Hz 0.96315 -0.239961
+ 3.55e+10Hz 0.962981 -0.240618
+ 3.56e+10Hz 0.96281 -0.241274
+ 3.57e+10Hz 0.96264 -0.241931
+ 3.58e+10Hz 0.962469 -0.242587
+ 3.59e+10Hz 0.962297 -0.243244
+ 3.6e+10Hz 0.962125 -0.2439
+ 3.61e+10Hz 0.961953 -0.244556
+ 3.62e+10Hz 0.96178 -0.245212
+ 3.63e+10Hz 0.961607 -0.245868
+ 3.64e+10Hz 0.961434 -0.246524
+ 3.65e+10Hz 0.96126 -0.247179
+ 3.66e+10Hz 0.961085 -0.247835
+ 3.67e+10Hz 0.960911 -0.24849
+ 3.68e+10Hz 0.960735 -0.249145
+ 3.69e+10Hz 0.96056 -0.249801
+ 3.7e+10Hz 0.960384 -0.250456
+ 3.71e+10Hz 0.960208 -0.251111
+ 3.72e+10Hz 0.960031 -0.251766
+ 3.73e+10Hz 0.959854 -0.252421
+ 3.74e+10Hz 0.959676 -0.253075
+ 3.75e+10Hz 0.959498 -0.25373
+ 3.76e+10Hz 0.959319 -0.254384
+ 3.77e+10Hz 0.95914 -0.255039
+ 3.78e+10Hz 0.958961 -0.255693
+ 3.79e+10Hz 0.958781 -0.256347
+ 3.8e+10Hz 0.958601 -0.257001
+ 3.81e+10Hz 0.958421 -0.257655
+ 3.82e+10Hz 0.95824 -0.258309
+ 3.83e+10Hz 0.958058 -0.258963
+ 3.84e+10Hz 0.957877 -0.259616
+ 3.85e+10Hz 0.957694 -0.26027
+ 3.86e+10Hz 0.957512 -0.260923
+ 3.87e+10Hz 0.957329 -0.261577
+ 3.88e+10Hz 0.957145 -0.26223
+ 3.89e+10Hz 0.956961 -0.262883
+ 3.9e+10Hz 0.956777 -0.263536
+ 3.91e+10Hz 0.956592 -0.264189
+ 3.92e+10Hz 0.956407 -0.264842
+ 3.93e+10Hz 0.956221 -0.265495
+ 3.94e+10Hz 0.956035 -0.266148
+ 3.95e+10Hz 0.955849 -0.2668
+ 3.96e+10Hz 0.955662 -0.267453
+ 3.97e+10Hz 0.955474 -0.268105
+ 3.98e+10Hz 0.955287 -0.268757
+ 3.99e+10Hz 0.955098 -0.26941
+ 4e+10Hz 0.95491 -0.270062
+ 4.01e+10Hz 0.95472 -0.270713
+ 4.02e+10Hz 0.954531 -0.271365
+ 4.03e+10Hz 0.954341 -0.272017
+ 4.04e+10Hz 0.954151 -0.272669
+ 4.05e+10Hz 0.95396 -0.27332
+ 4.06e+10Hz 0.953768 -0.273972
+ 4.07e+10Hz 0.953577 -0.274623
+ 4.08e+10Hz 0.953384 -0.275274
+ 4.09e+10Hz 0.953192 -0.275926
+ 4.1e+10Hz 0.952999 -0.276577
+ 4.11e+10Hz 0.952805 -0.277228
+ 4.12e+10Hz 0.952612 -0.277878
+ 4.13e+10Hz 0.952417 -0.278529
+ 4.14e+10Hz 0.952222 -0.27918
+ 4.15e+10Hz 0.952027 -0.27983
+ 4.16e+10Hz 0.951831 -0.280481
+ 4.17e+10Hz 0.951635 -0.281131
+ 4.18e+10Hz 0.951438 -0.281781
+ 4.19e+10Hz 0.951241 -0.282431
+ 4.2e+10Hz 0.951044 -0.283081
+ 4.21e+10Hz 0.950846 -0.283731
+ 4.22e+10Hz 0.950648 -0.284381
+ 4.23e+10Hz 0.950449 -0.285031
+ 4.24e+10Hz 0.950249 -0.28568
+ 4.25e+10Hz 0.95005 -0.28633
+ 4.26e+10Hz 0.94985 -0.286979
+ 4.27e+10Hz 0.949649 -0.287628
+ 4.28e+10Hz 0.949448 -0.288277
+ 4.29e+10Hz 0.949246 -0.288926
+ 4.3e+10Hz 0.949044 -0.289575
+ 4.31e+10Hz 0.948842 -0.290224
+ 4.32e+10Hz 0.948639 -0.290873
+ 4.33e+10Hz 0.948435 -0.291521
+ 4.34e+10Hz 0.948231 -0.29217
+ 4.35e+10Hz 0.948027 -0.292818
+ 4.36e+10Hz 0.947822 -0.293466
+ 4.37e+10Hz 0.947617 -0.294114
+ 4.38e+10Hz 0.947411 -0.294762
+ 4.39e+10Hz 0.947205 -0.29541
+ 4.4e+10Hz 0.946999 -0.296058
+ 4.41e+10Hz 0.946792 -0.296705
+ 4.42e+10Hz 0.946584 -0.297353
+ 4.43e+10Hz 0.946376 -0.298
+ 4.44e+10Hz 0.946168 -0.298647
+ 4.45e+10Hz 0.945959 -0.299294
+ 4.46e+10Hz 0.945749 -0.299941
+ 4.47e+10Hz 0.945539 -0.300588
+ 4.48e+10Hz 0.945329 -0.301234
+ 4.49e+10Hz 0.945118 -0.301881
+ 4.5e+10Hz 0.944907 -0.302527
+ 4.51e+10Hz 0.944695 -0.303174
+ 4.52e+10Hz 0.944483 -0.30382
+ 4.53e+10Hz 0.944271 -0.304466
+ 4.54e+10Hz 0.944057 -0.305111
+ 4.55e+10Hz 0.943844 -0.305757
+ 4.56e+10Hz 0.94363 -0.306403
+ 4.57e+10Hz 0.943415 -0.307048
+ 4.58e+10Hz 0.9432 -0.307694
+ 4.59e+10Hz 0.942985 -0.308339
+ 4.6e+10Hz 0.942769 -0.308984
+ 4.61e+10Hz 0.942553 -0.309628
+ 4.62e+10Hz 0.942336 -0.310273
+ 4.63e+10Hz 0.942119 -0.310918
+ 4.64e+10Hz 0.941901 -0.311562
+ 4.65e+10Hz 0.941683 -0.312206
+ 4.66e+10Hz 0.941464 -0.31285
+ 4.67e+10Hz 0.941245 -0.313494
+ 4.68e+10Hz 0.941026 -0.314138
+ 4.69e+10Hz 0.940805 -0.314782
+ 4.7e+10Hz 0.940585 -0.315425
+ 4.71e+10Hz 0.940364 -0.316069
+ 4.72e+10Hz 0.940143 -0.316712
+ 4.73e+10Hz 0.939921 -0.317355
+ 4.74e+10Hz 0.939698 -0.317998
+ 4.75e+10Hz 0.939476 -0.31864
+ 4.76e+10Hz 0.939252 -0.319283
+ 4.77e+10Hz 0.939029 -0.319925
+ 4.78e+10Hz 0.938804 -0.320568
+ 4.79e+10Hz 0.93858 -0.32121
+ 4.8e+10Hz 0.938355 -0.321852
+ 4.81e+10Hz 0.938129 -0.322493
+ 4.82e+10Hz 0.937903 -0.323135
+ 4.83e+10Hz 0.937677 -0.323776
+ 4.84e+10Hz 0.93745 -0.324418
+ 4.85e+10Hz 0.937222 -0.325058
+ 4.86e+10Hz 0.936994 -0.325699
+ 4.87e+10Hz 0.936766 -0.32634
+ 4.88e+10Hz 0.936537 -0.326981
+ 4.89e+10Hz 0.936308 -0.327621
+ 4.9e+10Hz 0.936079 -0.328261
+ 4.91e+10Hz 0.935848 -0.328901
+ 4.92e+10Hz 0.935618 -0.329541
+ 4.93e+10Hz 0.935387 -0.330181
+ 4.94e+10Hz 0.935155 -0.33082
+ 4.95e+10Hz 0.934923 -0.33146
+ 4.96e+10Hz 0.934691 -0.332099
+ 4.97e+10Hz 0.934458 -0.332738
+ 4.98e+10Hz 0.934225 -0.333377
+ 4.99e+10Hz 0.933991 -0.334015
+ 5e+10Hz 0.933757 -0.334654
+ 5.01e+10Hz 0.933522 -0.335292
+ 5.02e+10Hz 0.933287 -0.33593
+ 5.03e+10Hz 0.933052 -0.336568
+ 5.04e+10Hz 0.932816 -0.337206
+ 5.05e+10Hz 0.932579 -0.337843
+ 5.06e+10Hz 0.932342 -0.33848
+ 5.07e+10Hz 0.932105 -0.339118
+ 5.08e+10Hz 0.931867 -0.339755
+ 5.09e+10Hz 0.931629 -0.340391
+ 5.1e+10Hz 0.931391 -0.341028
+ 5.11e+10Hz 0.931152 -0.341664
+ 5.12e+10Hz 0.930912 -0.342301
+ 5.13e+10Hz 0.930672 -0.342937
+ 5.14e+10Hz 0.930432 -0.343573
+ 5.15e+10Hz 0.930191 -0.344208
+ 5.16e+10Hz 0.92995 -0.344844
+ 5.17e+10Hz 0.929708 -0.345479
+ 5.18e+10Hz 0.929466 -0.346114
+ 5.19e+10Hz 0.929223 -0.346749
+ 5.2e+10Hz 0.92898 -0.347384
+ 5.21e+10Hz 0.928737 -0.348018
+ 5.22e+10Hz 0.928493 -0.348653
+ 5.23e+10Hz 0.928249 -0.349287
+ 5.24e+10Hz 0.928004 -0.349921
+ 5.25e+10Hz 0.927759 -0.350554
+ 5.26e+10Hz 0.927513 -0.351188
+ 5.27e+10Hz 0.927267 -0.351822
+ 5.28e+10Hz 0.927021 -0.352455
+ 5.29e+10Hz 0.926774 -0.353088
+ 5.3e+10Hz 0.926527 -0.353721
+ 5.31e+10Hz 0.926279 -0.354353
+ 5.32e+10Hz 0.926031 -0.354986
+ 5.33e+10Hz 0.925782 -0.355618
+ 5.34e+10Hz 0.925533 -0.35625
+ 5.35e+10Hz 0.925284 -0.356882
+ 5.36e+10Hz 0.925034 -0.357513
+ 5.37e+10Hz 0.924783 -0.358145
+ 5.38e+10Hz 0.924533 -0.358776
+ 5.39e+10Hz 0.924282 -0.359407
+ 5.4e+10Hz 0.92403 -0.360038
+ 5.41e+10Hz 0.923778 -0.360669
+ 5.42e+10Hz 0.923526 -0.361299
+ 5.43e+10Hz 0.923273 -0.36193
+ 5.44e+10Hz 0.92302 -0.36256
+ 5.45e+10Hz 0.922766 -0.36319
+ 5.46e+10Hz 0.922512 -0.36382
+ 5.47e+10Hz 0.922258 -0.364449
+ 5.48e+10Hz 0.922003 -0.365079
+ 5.49e+10Hz 0.921747 -0.365708
+ 5.5e+10Hz 0.921492 -0.366337
+ 5.51e+10Hz 0.921235 -0.366966
+ 5.52e+10Hz 0.920979 -0.367594
+ 5.53e+10Hz 0.920722 -0.368223
+ 5.54e+10Hz 0.920465 -0.368851
+ 5.55e+10Hz 0.920207 -0.369479
+ 5.56e+10Hz 0.919949 -0.370107
+ 5.57e+10Hz 0.91969 -0.370734
+ 5.58e+10Hz 0.919431 -0.371362
+ 5.59e+10Hz 0.919171 -0.371989
+ 5.6e+10Hz 0.918912 -0.372616
+ 5.61e+10Hz 0.918651 -0.373243
+ 5.62e+10Hz 0.918391 -0.37387
+ 5.63e+10Hz 0.91813 -0.374496
+ 5.64e+10Hz 0.917868 -0.375123
+ 5.65e+10Hz 0.917606 -0.375749
+ 5.66e+10Hz 0.917344 -0.376375
+ 5.67e+10Hz 0.917081 -0.377
+ 5.68e+10Hz 0.916818 -0.377626
+ 5.69e+10Hz 0.916554 -0.378251
+ 5.7e+10Hz 0.91629 -0.378877
+ 5.71e+10Hz 0.916026 -0.379501
+ 5.72e+10Hz 0.915761 -0.380126
+ 5.73e+10Hz 0.915496 -0.380751
+ 5.74e+10Hz 0.91523 -0.381375
+ 5.75e+10Hz 0.914964 -0.382
+ 5.76e+10Hz 0.914698 -0.382624
+ 5.77e+10Hz 0.914431 -0.383248
+ 5.78e+10Hz 0.914164 -0.383871
+ 5.79e+10Hz 0.913896 -0.384495
+ 5.8e+10Hz 0.913628 -0.385118
+ 5.81e+10Hz 0.91336 -0.385741
+ 5.82e+10Hz 0.913091 -0.386364
+ 5.83e+10Hz 0.912822 -0.386987
+ 5.84e+10Hz 0.912552 -0.38761
+ 5.85e+10Hz 0.912282 -0.388232
+ 5.86e+10Hz 0.912011 -0.388854
+ 5.87e+10Hz 0.91174 -0.389476
+ 5.88e+10Hz 0.911469 -0.390098
+ 5.89e+10Hz 0.911197 -0.39072
+ 5.9e+10Hz 0.910925 -0.391341
+ 5.91e+10Hz 0.910653 -0.391962
+ 5.92e+10Hz 0.91038 -0.392584
+ 5.93e+10Hz 0.910107 -0.393205
+ 5.94e+10Hz 0.909833 -0.393825
+ 5.95e+10Hz 0.909559 -0.394446
+ 5.96e+10Hz 0.909284 -0.395066
+ 5.97e+10Hz 0.909009 -0.395686
+ 5.98e+10Hz 0.908734 -0.396307
+ 5.99e+10Hz 0.908458 -0.396926
+ 6e+10Hz 0.908182 -0.397546
+ 6.01e+10Hz 0.907905 -0.398166
+ 6.02e+10Hz 0.907628 -0.398785
+ 6.03e+10Hz 0.90735 -0.399404
+ 6.04e+10Hz 0.907073 -0.400023
+ 6.05e+10Hz 0.906794 -0.400641
+ 6.06e+10Hz 0.906516 -0.40126
+ 6.07e+10Hz 0.906237 -0.401879
+ 6.08e+10Hz 0.905957 -0.402497
+ 6.09e+10Hz 0.905677 -0.403115
+ 6.1e+10Hz 0.905397 -0.403732
+ 6.11e+10Hz 0.905116 -0.40435
+ 6.12e+10Hz 0.904835 -0.404968
+ 6.13e+10Hz 0.904554 -0.405585
+ 6.14e+10Hz 0.904272 -0.406202
+ 6.15e+10Hz 0.903989 -0.406819
+ 6.16e+10Hz 0.903706 -0.407436
+ 6.17e+10Hz 0.903423 -0.408052
+ 6.18e+10Hz 0.903139 -0.408669
+ 6.19e+10Hz 0.902855 -0.409285
+ 6.2e+10Hz 0.902571 -0.409901
+ 6.21e+10Hz 0.902286 -0.410517
+ 6.22e+10Hz 0.902001 -0.411132
+ 6.23e+10Hz 0.901715 -0.411748
+ 6.24e+10Hz 0.901429 -0.412363
+ 6.25e+10Hz 0.901142 -0.412978
+ 6.26e+10Hz 0.900855 -0.413593
+ 6.27e+10Hz 0.900568 -0.414208
+ 6.28e+10Hz 0.90028 -0.414822
+ 6.29e+10Hz 0.899992 -0.415437
+ 6.3e+10Hz 0.899703 -0.416051
+ 6.31e+10Hz 0.899414 -0.416665
+ 6.32e+10Hz 0.899125 -0.417279
+ 6.33e+10Hz 0.898835 -0.417892
+ 6.34e+10Hz 0.898545 -0.418506
+ 6.35e+10Hz 0.898254 -0.419119
+ 6.36e+10Hz 0.897963 -0.419732
+ 6.37e+10Hz 0.897671 -0.420345
+ 6.38e+10Hz 0.897379 -0.420958
+ 6.39e+10Hz 0.897087 -0.42157
+ 6.4e+10Hz 0.896794 -0.422183
+ 6.41e+10Hz 0.896501 -0.422795
+ 6.42e+10Hz 0.896207 -0.423407
+ 6.43e+10Hz 0.895913 -0.424018
+ 6.44e+10Hz 0.895618 -0.42463
+ 6.45e+10Hz 0.895323 -0.425241
+ 6.46e+10Hz 0.895028 -0.425853
+ 6.47e+10Hz 0.894732 -0.426463
+ 6.48e+10Hz 0.894436 -0.427074
+ 6.49e+10Hz 0.894139 -0.427685
+ 6.5e+10Hz 0.893842 -0.428295
+ 6.51e+10Hz 0.893545 -0.428905
+ 6.52e+10Hz 0.893247 -0.429516
+ 6.53e+10Hz 0.892949 -0.430125
+ 6.54e+10Hz 0.89265 -0.430735
+ 6.55e+10Hz 0.892351 -0.431345
+ 6.56e+10Hz 0.892051 -0.431954
+ 6.57e+10Hz 0.891751 -0.432563
+ 6.58e+10Hz 0.89145 -0.433172
+ 6.59e+10Hz 0.891149 -0.43378
+ 6.6e+10Hz 0.890848 -0.434389
+ 6.61e+10Hz 0.890546 -0.434997
+ 6.62e+10Hz 0.890244 -0.435605
+ 6.63e+10Hz 0.889941 -0.436213
+ 6.64e+10Hz 0.889638 -0.436821
+ 6.65e+10Hz 0.889335 -0.437428
+ 6.66e+10Hz 0.889031 -0.438035
+ 6.67e+10Hz 0.888726 -0.438642
+ 6.68e+10Hz 0.888422 -0.439249
+ 6.69e+10Hz 0.888116 -0.439856
+ 6.7e+10Hz 0.887811 -0.440462
+ 6.71e+10Hz 0.887505 -0.441069
+ 6.72e+10Hz 0.887198 -0.441675
+ 6.73e+10Hz 0.886891 -0.44228
+ 6.74e+10Hz 0.886584 -0.442886
+ 6.75e+10Hz 0.886276 -0.443491
+ 6.76e+10Hz 0.885968 -0.444097
+ 6.77e+10Hz 0.885659 -0.444702
+ 6.78e+10Hz 0.88535 -0.445306
+ 6.79e+10Hz 0.885041 -0.445911
+ 6.8e+10Hz 0.884731 -0.446515
+ 6.81e+10Hz 0.884421 -0.44712
+ 6.82e+10Hz 0.88411 -0.447723
+ 6.83e+10Hz 0.883798 -0.448327
+ 6.84e+10Hz 0.883487 -0.448931
+ 6.85e+10Hz 0.883175 -0.449534
+ 6.86e+10Hz 0.882862 -0.450137
+ 6.87e+10Hz 0.882549 -0.45074
+ 6.88e+10Hz 0.882236 -0.451342
+ 6.89e+10Hz 0.881922 -0.451945
+ 6.9e+10Hz 0.881608 -0.452547
+ 6.91e+10Hz 0.881293 -0.453149
+ 6.92e+10Hz 0.880978 -0.453751
+ 6.93e+10Hz 0.880663 -0.454352
+ 6.94e+10Hz 0.880347 -0.454954
+ 6.95e+10Hz 0.88003 -0.455555
+ 6.96e+10Hz 0.879713 -0.456156
+ 6.97e+10Hz 0.879396 -0.456756
+ 6.98e+10Hz 0.879078 -0.457357
+ 6.99e+10Hz 0.87876 -0.457957
+ 7e+10Hz 0.878442 -0.458557
+ 7.01e+10Hz 0.878123 -0.459157
+ 7.02e+10Hz 0.877803 -0.459756
+ 7.03e+10Hz 0.877484 -0.460355
+ 7.04e+10Hz 0.877163 -0.460954
+ 7.05e+10Hz 0.876843 -0.461553
+ 7.06e+10Hz 0.876522 -0.462152
+ 7.07e+10Hz 0.8762 -0.46275
+ 7.08e+10Hz 0.875878 -0.463348
+ 7.09e+10Hz 0.875556 -0.463946
+ 7.1e+10Hz 0.875233 -0.464544
+ 7.11e+10Hz 0.87491 -0.465141
+ 7.12e+10Hz 0.874586 -0.465739
+ 7.13e+10Hz 0.874262 -0.466336
+ 7.14e+10Hz 0.873938 -0.466932
+ 7.15e+10Hz 0.873613 -0.467529
+ 7.16e+10Hz 0.873287 -0.468125
+ 7.17e+10Hz 0.872962 -0.468721
+ 7.18e+10Hz 0.872636 -0.469317
+ 7.19e+10Hz 0.872309 -0.469912
+ 7.2e+10Hz 0.871982 -0.470508
+ 7.21e+10Hz 0.871655 -0.471103
+ 7.22e+10Hz 0.871327 -0.471697
+ 7.23e+10Hz 0.870999 -0.472292
+ 7.24e+10Hz 0.87067 -0.472886
+ 7.25e+10Hz 0.870341 -0.473481
+ 7.26e+10Hz 0.870011 -0.474074
+ 7.27e+10Hz 0.869681 -0.474668
+ 7.28e+10Hz 0.869351 -0.475261
+ 7.29e+10Hz 0.86902 -0.475854
+ 7.3e+10Hz 0.868689 -0.476447
+ 7.31e+10Hz 0.868358 -0.47704
+ 7.32e+10Hz 0.868026 -0.477632
+ 7.33e+10Hz 0.867693 -0.478224
+ 7.34e+10Hz 0.86736 -0.478816
+ 7.35e+10Hz 0.867027 -0.479408
+ 7.36e+10Hz 0.866694 -0.479999
+ 7.37e+10Hz 0.866359 -0.48059
+ 7.38e+10Hz 0.866025 -0.481181
+ 7.39e+10Hz 0.86569 -0.481772
+ 7.4e+10Hz 0.865355 -0.482362
+ 7.41e+10Hz 0.865019 -0.482952
+ 7.42e+10Hz 0.864683 -0.483542
+ 7.43e+10Hz 0.864347 -0.484132
+ 7.44e+10Hz 0.86401 -0.484721
+ 7.45e+10Hz 0.863672 -0.48531
+ 7.46e+10Hz 0.863335 -0.485899
+ 7.47e+10Hz 0.862997 -0.486488
+ 7.48e+10Hz 0.862658 -0.487076
+ 7.49e+10Hz 0.862319 -0.487665
+ 7.5e+10Hz 0.86198 -0.488252
+ 7.51e+10Hz 0.86164 -0.48884
+ 7.52e+10Hz 0.8613 -0.489427
+ 7.53e+10Hz 0.860959 -0.490015
+ 7.54e+10Hz 0.860618 -0.490601
+ 7.55e+10Hz 0.860277 -0.491188
+ 7.56e+10Hz 0.859935 -0.491774
+ 7.57e+10Hz 0.859593 -0.49236
+ 7.58e+10Hz 0.859251 -0.492946
+ 7.59e+10Hz 0.858908 -0.493532
+ 7.6e+10Hz 0.858564 -0.494117
+ 7.61e+10Hz 0.858221 -0.494702
+ 7.62e+10Hz 0.857877 -0.495287
+ 7.63e+10Hz 0.857532 -0.495872
+ 7.64e+10Hz 0.857187 -0.496456
+ 7.65e+10Hz 0.856842 -0.49704
+ 7.66e+10Hz 0.856496 -0.497624
+ 7.67e+10Hz 0.85615 -0.498208
+ 7.68e+10Hz 0.855804 -0.498791
+ 7.69e+10Hz 0.855457 -0.499374
+ 7.7e+10Hz 0.855109 -0.499957
+ 7.71e+10Hz 0.854762 -0.500539
+ 7.72e+10Hz 0.854414 -0.501122
+ 7.73e+10Hz 0.854065 -0.501704
+ 7.74e+10Hz 0.853716 -0.502285
+ 7.75e+10Hz 0.853367 -0.502867
+ 7.76e+10Hz 0.853018 -0.503448
+ 7.77e+10Hz 0.852668 -0.504029
+ 7.78e+10Hz 0.852317 -0.50461
+ 7.79e+10Hz 0.851966 -0.50519
+ 7.8e+10Hz 0.851615 -0.505771
+ 7.81e+10Hz 0.851264 -0.506351
+ 7.82e+10Hz 0.850912 -0.50693
+ 7.83e+10Hz 0.85056 -0.50751
+ 7.84e+10Hz 0.850207 -0.508089
+ 7.85e+10Hz 0.849854 -0.508668
+ 7.86e+10Hz 0.8495 -0.509247
+ 7.87e+10Hz 0.849147 -0.509825
+ 7.88e+10Hz 0.848792 -0.510404
+ 7.89e+10Hz 0.848438 -0.510982
+ 7.9e+10Hz 0.848083 -0.511559
+ 7.91e+10Hz 0.847727 -0.512137
+ 7.92e+10Hz 0.847372 -0.512714
+ 7.93e+10Hz 0.847015 -0.513291
+ 7.94e+10Hz 0.846659 -0.513868
+ 7.95e+10Hz 0.846302 -0.514444
+ 7.96e+10Hz 0.845945 -0.51502
+ 7.97e+10Hz 0.845587 -0.515596
+ 7.98e+10Hz 0.845229 -0.516172
+ 7.99e+10Hz 0.84487 -0.516748
+ 8e+10Hz 0.844512 -0.517323
+ 8.01e+10Hz 0.844152 -0.517898
+ 8.02e+10Hz 0.843793 -0.518472
+ 8.03e+10Hz 0.843433 -0.519047
+ 8.04e+10Hz 0.843073 -0.519621
+ 8.05e+10Hz 0.842712 -0.520195
+ 8.06e+10Hz 0.842351 -0.520769
+ 8.07e+10Hz 0.841989 -0.521342
+ 8.08e+10Hz 0.841627 -0.521915
+ 8.09e+10Hz 0.841265 -0.522488
+ 8.1e+10Hz 0.840903 -0.523061
+ 8.11e+10Hz 0.84054 -0.523633
+ 8.12e+10Hz 0.840176 -0.524206
+ 8.13e+10Hz 0.839813 -0.524778
+ 8.14e+10Hz 0.839448 -0.525349
+ 8.15e+10Hz 0.839084 -0.525921
+ 8.16e+10Hz 0.838719 -0.526492
+ 8.17e+10Hz 0.838354 -0.527063
+ 8.18e+10Hz 0.837988 -0.527634
+ 8.19e+10Hz 0.837622 -0.528204
+ 8.2e+10Hz 0.837256 -0.528774
+ 8.21e+10Hz 0.836889 -0.529344
+ 8.22e+10Hz 0.836522 -0.529914
+ 8.23e+10Hz 0.836154 -0.530483
+ 8.24e+10Hz 0.835786 -0.531053
+ 8.25e+10Hz 0.835418 -0.531622
+ 8.26e+10Hz 0.83505 -0.53219
+ 8.27e+10Hz 0.834681 -0.532759
+ 8.28e+10Hz 0.834311 -0.533327
+ 8.29e+10Hz 0.833941 -0.533895
+ 8.3e+10Hz 0.833571 -0.534463
+ 8.31e+10Hz 0.833201 -0.53503
+ 8.32e+10Hz 0.83283 -0.535597
+ 8.33e+10Hz 0.832458 -0.536165
+ 8.34e+10Hz 0.832087 -0.536731
+ 8.35e+10Hz 0.831715 -0.537298
+ 8.36e+10Hz 0.831342 -0.537864
+ 8.37e+10Hz 0.830969 -0.53843
+ 8.38e+10Hz 0.830596 -0.538996
+ 8.39e+10Hz 0.830222 -0.539561
+ 8.4e+10Hz 0.829848 -0.540127
+ 8.41e+10Hz 0.829474 -0.540692
+ 8.42e+10Hz 0.829099 -0.541256
+ 8.43e+10Hz 0.828724 -0.541821
+ 8.44e+10Hz 0.828349 -0.542385
+ 8.45e+10Hz 0.827973 -0.542949
+ 8.46e+10Hz 0.827597 -0.543513
+ 8.47e+10Hz 0.82722 -0.544077
+ 8.48e+10Hz 0.826843 -0.54464
+ 8.49e+10Hz 0.826466 -0.545203
+ 8.5e+10Hz 0.826088 -0.545766
+ 8.51e+10Hz 0.82571 -0.546328
+ 8.52e+10Hz 0.825331 -0.546891
+ 8.53e+10Hz 0.824952 -0.547453
+ 8.54e+10Hz 0.824573 -0.548015
+ 8.55e+10Hz 0.824193 -0.548576
+ 8.56e+10Hz 0.823813 -0.549137
+ 8.57e+10Hz 0.823433 -0.549699
+ 8.58e+10Hz 0.823052 -0.550259
+ 8.59e+10Hz 0.82267 -0.55082
+ 8.6e+10Hz 0.822289 -0.55138
+ 8.61e+10Hz 0.821907 -0.55194
+ 8.62e+10Hz 0.821524 -0.5525
+ 8.63e+10Hz 0.821142 -0.55306
+ 8.64e+10Hz 0.820758 -0.553619
+ 8.65e+10Hz 0.820375 -0.554178
+ 8.66e+10Hz 0.819991 -0.554737
+ 8.67e+10Hz 0.819607 -0.555296
+ 8.68e+10Hz 0.819222 -0.555854
+ 8.69e+10Hz 0.818837 -0.556412
+ 8.7e+10Hz 0.818451 -0.55697
+ 8.71e+10Hz 0.818065 -0.557527
+ 8.72e+10Hz 0.817679 -0.558085
+ 8.73e+10Hz 0.817292 -0.558642
+ 8.74e+10Hz 0.816905 -0.559199
+ 8.75e+10Hz 0.816518 -0.559755
+ 8.76e+10Hz 0.81613 -0.560312
+ 8.77e+10Hz 0.815742 -0.560868
+ 8.78e+10Hz 0.815353 -0.561423
+ 8.79e+10Hz 0.814964 -0.561979
+ 8.8e+10Hz 0.814575 -0.562534
+ 8.81e+10Hz 0.814185 -0.563089
+ 8.82e+10Hz 0.813795 -0.563644
+ 8.83e+10Hz 0.813404 -0.564199
+ 8.84e+10Hz 0.813013 -0.564753
+ 8.85e+10Hz 0.812622 -0.565307
+ 8.86e+10Hz 0.81223 -0.565861
+ 8.87e+10Hz 0.811838 -0.566414
+ 8.88e+10Hz 0.811446 -0.566967
+ 8.89e+10Hz 0.811053 -0.56752
+ 8.9e+10Hz 0.810659 -0.568073
+ 8.91e+10Hz 0.810266 -0.568626
+ 8.92e+10Hz 0.809871 -0.569178
+ 8.93e+10Hz 0.809477 -0.56973
+ 8.94e+10Hz 0.809082 -0.570281
+ 8.95e+10Hz 0.808687 -0.570833
+ 8.96e+10Hz 0.808291 -0.571384
+ 8.97e+10Hz 0.807895 -0.571935
+ 8.98e+10Hz 0.807499 -0.572485
+ 8.99e+10Hz 0.807102 -0.573036
+ 9e+10Hz 0.806705 -0.573586
+ 9.01e+10Hz 0.806307 -0.574136
+ 9.02e+10Hz 0.805909 -0.574685
+ 9.03e+10Hz 0.80551 -0.575234
+ 9.04e+10Hz 0.805112 -0.575783
+ 9.05e+10Hz 0.804712 -0.576332
+ 9.06e+10Hz 0.804313 -0.57688
+ 9.07e+10Hz 0.803913 -0.577429
+ 9.08e+10Hz 0.803512 -0.577977
+ 9.09e+10Hz 0.803112 -0.578524
+ 9.1e+10Hz 0.80271 -0.579071
+ 9.11e+10Hz 0.802309 -0.579619
+ 9.12e+10Hz 0.801907 -0.580165
+ 9.13e+10Hz 0.801504 -0.580712
+ 9.14e+10Hz 0.801102 -0.581258
+ 9.15e+10Hz 0.800699 -0.581804
+ 9.16e+10Hz 0.800295 -0.58235
+ 9.17e+10Hz 0.799891 -0.582895
+ 9.18e+10Hz 0.799487 -0.58344
+ 9.19e+10Hz 0.799082 -0.583985
+ 9.2e+10Hz 0.798677 -0.58453
+ 9.21e+10Hz 0.798271 -0.585074
+ 9.22e+10Hz 0.797866 -0.585618
+ 9.23e+10Hz 0.797459 -0.586162
+ 9.24e+10Hz 0.797053 -0.586705
+ 9.25e+10Hz 0.796646 -0.587248
+ 9.26e+10Hz 0.796238 -0.587791
+ 9.27e+10Hz 0.79583 -0.588334
+ 9.28e+10Hz 0.795422 -0.588876
+ 9.29e+10Hz 0.795013 -0.589418
+ 9.3e+10Hz 0.794604 -0.58996
+ 9.31e+10Hz 0.794195 -0.590501
+ 9.32e+10Hz 0.793785 -0.591043
+ 9.33e+10Hz 0.793375 -0.591583
+ 9.34e+10Hz 0.792964 -0.592124
+ 9.35e+10Hz 0.792553 -0.592664
+ 9.36e+10Hz 0.792142 -0.593204
+ 9.37e+10Hz 0.79173 -0.593744
+ 9.38e+10Hz 0.791318 -0.594283
+ 9.39e+10Hz 0.790906 -0.594822
+ 9.4e+10Hz 0.790493 -0.595361
+ 9.41e+10Hz 0.79008 -0.5959
+ 9.42e+10Hz 0.789666 -0.596438
+ 9.43e+10Hz 0.789252 -0.596976
+ 9.44e+10Hz 0.788837 -0.597513
+ 9.45e+10Hz 0.788423 -0.598051
+ 9.46e+10Hz 0.788007 -0.598588
+ 9.47e+10Hz 0.787592 -0.599124
+ 9.48e+10Hz 0.787176 -0.599661
+ 9.49e+10Hz 0.78676 -0.600197
+ 9.5e+10Hz 0.786343 -0.600733
+ 9.51e+10Hz 0.785926 -0.601268
+ 9.52e+10Hz 0.785508 -0.601804
+ 9.53e+10Hz 0.785091 -0.602338
+ 9.54e+10Hz 0.784672 -0.602873
+ 9.55e+10Hz 0.784254 -0.603407
+ 9.56e+10Hz 0.783835 -0.603941
+ 9.57e+10Hz 0.783415 -0.604475
+ 9.58e+10Hz 0.782996 -0.605008
+ 9.59e+10Hz 0.782576 -0.605541
+ 9.6e+10Hz 0.782155 -0.606074
+ 9.61e+10Hz 0.781734 -0.606607
+ 9.62e+10Hz 0.781313 -0.607139
+ 9.63e+10Hz 0.780891 -0.607671
+ 9.64e+10Hz 0.78047 -0.608202
+ 9.65e+10Hz 0.780047 -0.608734
+ 9.66e+10Hz 0.779625 -0.609264
+ 9.67e+10Hz 0.779201 -0.609795
+ 9.68e+10Hz 0.778778 -0.610325
+ 9.69e+10Hz 0.778354 -0.610855
+ 9.7e+10Hz 0.77793 -0.611385
+ 9.71e+10Hz 0.777505 -0.611914
+ 9.72e+10Hz 0.777081 -0.612443
+ 9.73e+10Hz 0.776655 -0.612972
+ 9.74e+10Hz 0.77623 -0.613501
+ 9.75e+10Hz 0.775804 -0.614029
+ 9.76e+10Hz 0.775377 -0.614556
+ 9.77e+10Hz 0.774951 -0.615084
+ 9.78e+10Hz 0.774524 -0.615611
+ 9.79e+10Hz 0.774096 -0.616138
+ 9.8e+10Hz 0.773668 -0.616665
+ 9.81e+10Hz 0.77324 -0.617191
+ 9.82e+10Hz 0.772812 -0.617717
+ 9.83e+10Hz 0.772383 -0.618242
+ 9.84e+10Hz 0.771953 -0.618768
+ 9.85e+10Hz 0.771524 -0.619293
+ 9.86e+10Hz 0.771094 -0.619817
+ 9.87e+10Hz 0.770664 -0.620342
+ 9.88e+10Hz 0.770233 -0.620866
+ 9.89e+10Hz 0.769802 -0.62139
+ 9.9e+10Hz 0.769371 -0.621913
+ 9.91e+10Hz 0.768939 -0.622436
+ 9.92e+10Hz 0.768507 -0.622959
+ 9.93e+10Hz 0.768075 -0.623481
+ 9.94e+10Hz 0.767642 -0.624004
+ 9.95e+10Hz 0.767209 -0.624525
+ 9.96e+10Hz 0.766775 -0.625047
+ 9.97e+10Hz 0.766342 -0.625568
+ 9.98e+10Hz 0.765907 -0.626089
+ 9.99e+10Hz 0.765473 -0.62661
+ 1e+11Hz 0.765038 -0.62713
+ 1.001e+11Hz 0.764603 -0.62765
+ 1.002e+11Hz 0.764167 -0.628169
+ 1.003e+11Hz 0.763732 -0.628689
+ 1.004e+11Hz 0.763295 -0.629208
+ 1.005e+11Hz 0.762859 -0.629726
+ 1.006e+11Hz 0.762422 -0.630245
+ 1.007e+11Hz 0.761985 -0.630763
+ 1.008e+11Hz 0.761547 -0.631281
+ 1.009e+11Hz 0.761109 -0.631798
+ 1.01e+11Hz 0.760671 -0.632315
+ 1.011e+11Hz 0.760232 -0.632832
+ 1.012e+11Hz 0.759794 -0.633349
+ 1.013e+11Hz 0.759354 -0.633865
+ 1.014e+11Hz 0.758915 -0.634381
+ 1.015e+11Hz 0.758475 -0.634896
+ 1.016e+11Hz 0.758035 -0.635412
+ 1.017e+11Hz 0.757594 -0.635926
+ 1.018e+11Hz 0.757153 -0.636441
+ 1.019e+11Hz 0.756712 -0.636956
+ 1.02e+11Hz 0.75627 -0.63747
+ 1.021e+11Hz 0.755828 -0.637983
+ 1.022e+11Hz 0.755386 -0.638497
+ 1.023e+11Hz 0.754943 -0.63901
+ 1.024e+11Hz 0.7545 -0.639522
+ 1.025e+11Hz 0.754057 -0.640035
+ 1.026e+11Hz 0.753614 -0.640547
+ 1.027e+11Hz 0.75317 -0.641059
+ 1.028e+11Hz 0.752725 -0.641571
+ 1.029e+11Hz 0.752281 -0.642082
+ 1.03e+11Hz 0.751836 -0.642593
+ 1.031e+11Hz 0.751391 -0.643103
+ 1.032e+11Hz 0.750945 -0.643614
+ 1.033e+11Hz 0.750499 -0.644124
+ 1.034e+11Hz 0.750053 -0.644633
+ 1.035e+11Hz 0.749606 -0.645143
+ 1.036e+11Hz 0.749159 -0.645652
+ 1.037e+11Hz 0.748712 -0.646161
+ 1.038e+11Hz 0.748265 -0.646669
+ 1.039e+11Hz 0.747817 -0.647177
+ 1.04e+11Hz 0.747369 -0.647685
+ 1.041e+11Hz 0.74692 -0.648193
+ 1.042e+11Hz 0.746471 -0.6487
+ 1.043e+11Hz 0.746022 -0.649207
+ 1.044e+11Hz 0.745572 -0.649714
+ 1.045e+11Hz 0.745123 -0.65022
+ 1.046e+11Hz 0.744672 -0.650726
+ 1.047e+11Hz 0.744222 -0.651232
+ 1.048e+11Hz 0.743771 -0.651738
+ 1.049e+11Hz 0.74332 -0.652243
+ 1.05e+11Hz 0.742869 -0.652748
+ 1.051e+11Hz 0.742417 -0.653252
+ 1.052e+11Hz 0.741965 -0.653757
+ 1.053e+11Hz 0.741512 -0.654261
+ 1.054e+11Hz 0.741059 -0.654764
+ 1.055e+11Hz 0.740606 -0.655268
+ 1.056e+11Hz 0.740153 -0.655771
+ 1.057e+11Hz 0.739699 -0.656274
+ 1.058e+11Hz 0.739245 -0.656776
+ 1.059e+11Hz 0.738791 -0.657278
+ 1.06e+11Hz 0.738336 -0.65778
+ 1.061e+11Hz 0.737881 -0.658282
+ 1.062e+11Hz 0.737425 -0.658783
+ 1.063e+11Hz 0.73697 -0.659284
+ 1.064e+11Hz 0.736513 -0.659785
+ 1.065e+11Hz 0.736057 -0.660285
+ 1.066e+11Hz 0.7356 -0.660785
+ 1.067e+11Hz 0.735143 -0.661285
+ 1.068e+11Hz 0.734686 -0.661785
+ 1.069e+11Hz 0.734228 -0.662284
+ 1.07e+11Hz 0.73377 -0.662783
+ 1.071e+11Hz 0.733312 -0.663282
+ 1.072e+11Hz 0.732853 -0.66378
+ 1.073e+11Hz 0.732394 -0.664278
+ 1.074e+11Hz 0.731935 -0.664776
+ 1.075e+11Hz 0.731475 -0.665273
+ 1.076e+11Hz 0.731015 -0.66577
+ 1.077e+11Hz 0.730554 -0.666267
+ 1.078e+11Hz 0.730094 -0.666764
+ 1.079e+11Hz 0.729633 -0.66726
+ 1.08e+11Hz 0.729171 -0.667756
+ 1.081e+11Hz 0.72871 -0.668252
+ 1.082e+11Hz 0.728248 -0.668747
+ 1.083e+11Hz 0.727785 -0.669242
+ 1.084e+11Hz 0.727322 -0.669737
+ 1.085e+11Hz 0.726859 -0.670232
+ 1.086e+11Hz 0.726396 -0.670726
+ 1.087e+11Hz 0.725932 -0.67122
+ 1.088e+11Hz 0.725468 -0.671714
+ 1.089e+11Hz 0.725004 -0.672207
+ 1.09e+11Hz 0.724539 -0.6727
+ 1.091e+11Hz 0.724074 -0.673193
+ 1.092e+11Hz 0.723608 -0.673685
+ 1.093e+11Hz 0.723143 -0.674177
+ 1.094e+11Hz 0.722677 -0.674669
+ 1.095e+11Hz 0.72221 -0.675161
+ 1.096e+11Hz 0.721743 -0.675652
+ 1.097e+11Hz 0.721276 -0.676143
+ 1.098e+11Hz 0.720809 -0.676634
+ 1.099e+11Hz 0.720341 -0.677124
+ 1.1e+11Hz 0.719873 -0.677614
+ 1.101e+11Hz 0.719404 -0.678104
+ 1.102e+11Hz 0.718935 -0.678594
+ 1.103e+11Hz 0.718466 -0.679083
+ 1.104e+11Hz 0.717997 -0.679572
+ 1.105e+11Hz 0.717527 -0.68006
+ 1.106e+11Hz 0.717057 -0.680549
+ 1.107e+11Hz 0.716586 -0.681037
+ 1.108e+11Hz 0.716115 -0.681524
+ 1.109e+11Hz 0.715644 -0.682012
+ 1.11e+11Hz 0.715172 -0.682499
+ 1.111e+11Hz 0.7147 -0.682986
+ 1.112e+11Hz 0.714228 -0.683472
+ 1.113e+11Hz 0.713755 -0.683958
+ 1.114e+11Hz 0.713282 -0.684444
+ 1.115e+11Hz 0.712809 -0.68493
+ 1.116e+11Hz 0.712335 -0.685415
+ 1.117e+11Hz 0.711861 -0.6859
+ 1.118e+11Hz 0.711387 -0.686384
+ 1.119e+11Hz 0.710912 -0.686869
+ 1.12e+11Hz 0.710437 -0.687353
+ 1.121e+11Hz 0.709961 -0.687837
+ 1.122e+11Hz 0.709486 -0.68832
+ 1.123e+11Hz 0.709009 -0.688803
+ 1.124e+11Hz 0.708533 -0.689286
+ 1.125e+11Hz 0.708056 -0.689768
+ 1.126e+11Hz 0.707579 -0.69025
+ 1.127e+11Hz 0.707101 -0.690732
+ 1.128e+11Hz 0.706623 -0.691214
+ 1.129e+11Hz 0.706145 -0.691695
+ 1.13e+11Hz 0.705666 -0.692176
+ 1.131e+11Hz 0.705187 -0.692657
+ 1.132e+11Hz 0.704708 -0.693137
+ 1.133e+11Hz 0.704228 -0.693617
+ 1.134e+11Hz 0.703748 -0.694096
+ 1.135e+11Hz 0.703268 -0.694576
+ 1.136e+11Hz 0.702787 -0.695055
+ 1.137e+11Hz 0.702306 -0.695533
+ 1.138e+11Hz 0.701825 -0.696012
+ 1.139e+11Hz 0.701343 -0.696489
+ 1.14e+11Hz 0.700861 -0.696967
+ 1.141e+11Hz 0.700378 -0.697445
+ 1.142e+11Hz 0.699895 -0.697921
+ 1.143e+11Hz 0.699412 -0.698398
+ 1.144e+11Hz 0.698928 -0.698874
+ 1.145e+11Hz 0.698445 -0.69935
+ 1.146e+11Hz 0.69796 -0.699826
+ 1.147e+11Hz 0.697476 -0.700302
+ 1.148e+11Hz 0.696991 -0.700777
+ 1.149e+11Hz 0.696505 -0.701251
+ 1.15e+11Hz 0.69602 -0.701726
+ 1.151e+11Hz 0.695534 -0.7022
+ 1.152e+11Hz 0.695047 -0.702673
+ 1.153e+11Hz 0.69456 -0.703147
+ 1.154e+11Hz 0.694073 -0.703619
+ 1.155e+11Hz 0.693586 -0.704092
+ 1.156e+11Hz 0.693098 -0.704565
+ 1.157e+11Hz 0.69261 -0.705036
+ 1.158e+11Hz 0.692121 -0.705508
+ 1.159e+11Hz 0.691632 -0.705979
+ 1.16e+11Hz 0.691143 -0.70645
+ 1.161e+11Hz 0.690654 -0.706921
+ 1.162e+11Hz 0.690164 -0.707391
+ 1.163e+11Hz 0.689673 -0.707861
+ 1.164e+11Hz 0.689183 -0.70833
+ 1.165e+11Hz 0.688692 -0.7088
+ 1.166e+11Hz 0.6882 -0.709268
+ 1.167e+11Hz 0.687709 -0.709737
+ 1.168e+11Hz 0.687217 -0.710205
+ 1.169e+11Hz 0.686725 -0.710673
+ 1.17e+11Hz 0.686232 -0.71114
+ 1.171e+11Hz 0.685739 -0.711607
+ 1.172e+11Hz 0.685245 -0.712074
+ 1.173e+11Hz 0.684752 -0.71254
+ 1.174e+11Hz 0.684258 -0.713006
+ 1.175e+11Hz 0.683763 -0.713471
+ 1.176e+11Hz 0.683269 -0.713937
+ 1.177e+11Hz 0.682774 -0.714401
+ 1.178e+11Hz 0.682278 -0.714866
+ 1.179e+11Hz 0.681782 -0.71533
+ 1.18e+11Hz 0.681286 -0.715794
+ 1.181e+11Hz 0.68079 -0.716257
+ 1.182e+11Hz 0.680293 -0.71672
+ 1.183e+11Hz 0.679796 -0.717183
+ 1.184e+11Hz 0.679299 -0.717645
+ 1.185e+11Hz 0.678801 -0.718107
+ 1.186e+11Hz 0.678303 -0.718569
+ 1.187e+11Hz 0.677805 -0.71903
+ 1.188e+11Hz 0.677306 -0.71949
+ 1.189e+11Hz 0.676807 -0.719951
+ 1.19e+11Hz 0.676307 -0.720411
+ 1.191e+11Hz 0.675808 -0.72087
+ 1.192e+11Hz 0.675308 -0.72133
+ 1.193e+11Hz 0.674807 -0.721789
+ 1.194e+11Hz 0.674307 -0.722247
+ 1.195e+11Hz 0.673806 -0.722705
+ 1.196e+11Hz 0.673304 -0.723163
+ 1.197e+11Hz 0.672803 -0.72362
+ 1.198e+11Hz 0.672301 -0.724078
+ 1.199e+11Hz 0.671799 -0.724534
+ 1.2e+11Hz 0.671296 -0.72499
+ 1.201e+11Hz 0.670793 -0.725446
+ 1.202e+11Hz 0.67029 -0.725902
+ 1.203e+11Hz 0.669786 -0.726357
+ 1.204e+11Hz 0.669283 -0.726812
+ 1.205e+11Hz 0.668779 -0.727266
+ 1.206e+11Hz 0.668274 -0.72772
+ 1.207e+11Hz 0.667769 -0.728174
+ 1.208e+11Hz 0.667264 -0.728627
+ 1.209e+11Hz 0.666759 -0.729079
+ 1.21e+11Hz 0.666253 -0.729532
+ 1.211e+11Hz 0.665748 -0.729984
+ 1.212e+11Hz 0.665241 -0.730436
+ 1.213e+11Hz 0.664735 -0.730887
+ 1.214e+11Hz 0.664228 -0.731338
+ 1.215e+11Hz 0.663721 -0.731788
+ 1.216e+11Hz 0.663213 -0.732239
+ 1.217e+11Hz 0.662705 -0.732688
+ 1.218e+11Hz 0.662197 -0.733138
+ 1.219e+11Hz 0.661689 -0.733587
+ 1.22e+11Hz 0.661181 -0.734035
+ 1.221e+11Hz 0.660672 -0.734483
+ 1.222e+11Hz 0.660162 -0.734931
+ 1.223e+11Hz 0.659653 -0.735379
+ 1.224e+11Hz 0.659143 -0.735826
+ 1.225e+11Hz 0.658633 -0.736272
+ 1.226e+11Hz 0.658123 -0.736719
+ 1.227e+11Hz 0.657612 -0.737165
+ 1.228e+11Hz 0.657102 -0.73761
+ 1.229e+11Hz 0.65659 -0.738055
+ 1.23e+11Hz 0.656079 -0.7385
+ 1.231e+11Hz 0.655567 -0.738944
+ 1.232e+11Hz 0.655055 -0.739388
+ 1.233e+11Hz 0.654543 -0.739832
+ 1.234e+11Hz 0.65403 -0.740275
+ 1.235e+11Hz 0.653518 -0.740718
+ 1.236e+11Hz 0.653004 -0.741161
+ 1.237e+11Hz 0.652491 -0.741603
+ 1.238e+11Hz 0.651978 -0.742044
+ 1.239e+11Hz 0.651464 -0.742486
+ 1.24e+11Hz 0.650949 -0.742927
+ 1.241e+11Hz 0.650435 -0.743367
+ 1.242e+11Hz 0.64992 -0.743808
+ 1.243e+11Hz 0.649405 -0.744247
+ 1.244e+11Hz 0.64889 -0.744687
+ 1.245e+11Hz 0.648375 -0.745126
+ 1.246e+11Hz 0.647859 -0.745565
+ 1.247e+11Hz 0.647343 -0.746003
+ 1.248e+11Hz 0.646827 -0.746441
+ 1.249e+11Hz 0.64631 -0.746879
+ 1.25e+11Hz 0.645793 -0.747316
+ 1.251e+11Hz 0.645276 -0.747753
+ 1.252e+11Hz 0.644759 -0.748189
+ 1.253e+11Hz 0.644242 -0.748625
+ 1.254e+11Hz 0.643724 -0.749061
+ 1.255e+11Hz 0.643206 -0.749497
+ 1.256e+11Hz 0.642687 -0.749932
+ 1.257e+11Hz 0.642169 -0.750366
+ 1.258e+11Hz 0.64165 -0.750801
+ 1.259e+11Hz 0.641131 -0.751235
+ 1.26e+11Hz 0.640611 -0.751668
+ 1.261e+11Hz 0.640092 -0.752101
+ 1.262e+11Hz 0.639572 -0.752534
+ 1.263e+11Hz 0.639052 -0.752967
+ 1.264e+11Hz 0.638532 -0.753399
+ 1.265e+11Hz 0.638011 -0.753831
+ 1.266e+11Hz 0.63749 -0.754262
+ 1.267e+11Hz 0.636969 -0.754693
+ 1.268e+11Hz 0.636448 -0.755124
+ 1.269e+11Hz 0.635926 -0.755555
+ 1.27e+11Hz 0.635404 -0.755985
+ 1.271e+11Hz 0.634882 -0.756414
+ 1.272e+11Hz 0.63436 -0.756844
+ 1.273e+11Hz 0.633837 -0.757273
+ 1.274e+11Hz 0.633314 -0.757701
+ 1.275e+11Hz 0.632791 -0.75813
+ 1.276e+11Hz 0.632268 -0.758558
+ 1.277e+11Hz 0.631744 -0.758985
+ 1.278e+11Hz 0.63122 -0.759413
+ 1.279e+11Hz 0.630696 -0.75984
+ 1.28e+11Hz 0.630172 -0.760266
+ 1.281e+11Hz 0.629647 -0.760692
+ 1.282e+11Hz 0.629122 -0.761118
+ 1.283e+11Hz 0.628597 -0.761544
+ 1.284e+11Hz 0.628072 -0.761969
+ 1.285e+11Hz 0.627546 -0.762394
+ 1.286e+11Hz 0.62702 -0.762819
+ 1.287e+11Hz 0.626494 -0.763243
+ 1.288e+11Hz 0.625967 -0.763667
+ 1.289e+11Hz 0.625441 -0.76409
+ 1.29e+11Hz 0.624914 -0.764514
+ 1.291e+11Hz 0.624387 -0.764937
+ 1.292e+11Hz 0.623859 -0.765359
+ 1.293e+11Hz 0.623332 -0.765781
+ 1.294e+11Hz 0.622804 -0.766203
+ 1.295e+11Hz 0.622275 -0.766625
+ 1.296e+11Hz 0.621747 -0.767046
+ 1.297e+11Hz 0.621218 -0.767467
+ 1.298e+11Hz 0.620689 -0.767888
+ 1.299e+11Hz 0.62016 -0.768308
+ 1.3e+11Hz 0.61963 -0.768728
+ 1.301e+11Hz 0.619101 -0.769148
+ 1.302e+11Hz 0.618571 -0.769567
+ 1.303e+11Hz 0.61804 -0.769986
+ 1.304e+11Hz 0.61751 -0.770405
+ 1.305e+11Hz 0.616979 -0.770823
+ 1.306e+11Hz 0.616448 -0.771241
+ 1.307e+11Hz 0.615916 -0.771659
+ 1.308e+11Hz 0.615385 -0.772076
+ 1.309e+11Hz 0.614853 -0.772493
+ 1.31e+11Hz 0.61432 -0.77291
+ 1.311e+11Hz 0.613788 -0.773327
+ 1.312e+11Hz 0.613255 -0.773743
+ 1.313e+11Hz 0.612722 -0.774158
+ 1.314e+11Hz 0.612189 -0.774574
+ 1.315e+11Hz 0.611655 -0.774989
+ 1.316e+11Hz 0.611121 -0.775404
+ 1.317e+11Hz 0.610587 -0.775818
+ 1.318e+11Hz 0.610052 -0.776233
+ 1.319e+11Hz 0.609518 -0.776647
+ 1.32e+11Hz 0.608983 -0.77706
+ 1.321e+11Hz 0.608447 -0.777474
+ 1.322e+11Hz 0.607912 -0.777886
+ 1.323e+11Hz 0.607376 -0.778299
+ 1.324e+11Hz 0.60684 -0.778711
+ 1.325e+11Hz 0.606303 -0.779123
+ 1.326e+11Hz 0.605766 -0.779535
+ 1.327e+11Hz 0.605229 -0.779946
+ 1.328e+11Hz 0.604692 -0.780357
+ 1.329e+11Hz 0.604154 -0.780768
+ 1.33e+11Hz 0.603616 -0.781178
+ 1.331e+11Hz 0.603078 -0.781589
+ 1.332e+11Hz 0.602539 -0.781998
+ 1.333e+11Hz 0.602 -0.782408
+ 1.334e+11Hz 0.601461 -0.782817
+ 1.335e+11Hz 0.600922 -0.783226
+ 1.336e+11Hz 0.600382 -0.783634
+ 1.337e+11Hz 0.599842 -0.784042
+ 1.338e+11Hz 0.599301 -0.78445
+ 1.339e+11Hz 0.598761 -0.784857
+ 1.34e+11Hz 0.598219 -0.785265
+ 1.341e+11Hz 0.597678 -0.785671
+ 1.342e+11Hz 0.597136 -0.786078
+ 1.343e+11Hz 0.596594 -0.786484
+ 1.344e+11Hz 0.596052 -0.78689
+ 1.345e+11Hz 0.595509 -0.787295
+ 1.346e+11Hz 0.594966 -0.787701
+ 1.347e+11Hz 0.594423 -0.788105
+ 1.348e+11Hz 0.593879 -0.78851
+ 1.349e+11Hz 0.593335 -0.788914
+ 1.35e+11Hz 0.592791 -0.789318
+ 1.351e+11Hz 0.592246 -0.789721
+ 1.352e+11Hz 0.591701 -0.790124
+ 1.353e+11Hz 0.591156 -0.790527
+ 1.354e+11Hz 0.590611 -0.790929
+ 1.355e+11Hz 0.590064 -0.791331
+ 1.356e+11Hz 0.589518 -0.791733
+ 1.357e+11Hz 0.588972 -0.792135
+ 1.358e+11Hz 0.588425 -0.792536
+ 1.359e+11Hz 0.587877 -0.792936
+ 1.36e+11Hz 0.58733 -0.793337
+ 1.361e+11Hz 0.586782 -0.793737
+ 1.362e+11Hz 0.586233 -0.794136
+ 1.363e+11Hz 0.585685 -0.794535
+ 1.364e+11Hz 0.585136 -0.794934
+ 1.365e+11Hz 0.584586 -0.795333
+ 1.366e+11Hz 0.584037 -0.795731
+ 1.367e+11Hz 0.583487 -0.796129
+ 1.368e+11Hz 0.582936 -0.796526
+ 1.369e+11Hz 0.582386 -0.796923
+ 1.37e+11Hz 0.581835 -0.79732
+ 1.371e+11Hz 0.581283 -0.797716
+ 1.372e+11Hz 0.580731 -0.798112
+ 1.373e+11Hz 0.580179 -0.798507
+ 1.374e+11Hz 0.579627 -0.798902
+ 1.375e+11Hz 0.579074 -0.799297
+ 1.376e+11Hz 0.578521 -0.799691
+ 1.377e+11Hz 0.577968 -0.800085
+ 1.378e+11Hz 0.577414 -0.800479
+ 1.379e+11Hz 0.57686 -0.800872
+ 1.38e+11Hz 0.576305 -0.801265
+ 1.381e+11Hz 0.57575 -0.801657
+ 1.382e+11Hz 0.575195 -0.802049
+ 1.383e+11Hz 0.574639 -0.802441
+ 1.384e+11Hz 0.574084 -0.802832
+ 1.385e+11Hz 0.573527 -0.803223
+ 1.386e+11Hz 0.572971 -0.803613
+ 1.387e+11Hz 0.572414 -0.804003
+ 1.388e+11Hz 0.571857 -0.804392
+ 1.389e+11Hz 0.571299 -0.804781
+ 1.39e+11Hz 0.570741 -0.80517
+ 1.391e+11Hz 0.570183 -0.805558
+ 1.392e+11Hz 0.569624 -0.805946
+ 1.393e+11Hz 0.569065 -0.806333
+ 1.394e+11Hz 0.568506 -0.80672
+ 1.395e+11Hz 0.567946 -0.807107
+ 1.396e+11Hz 0.567386 -0.807493
+ 1.397e+11Hz 0.566826 -0.807879
+ 1.398e+11Hz 0.566265 -0.808264
+ 1.399e+11Hz 0.565704 -0.808648
+ 1.4e+11Hz 0.565143 -0.809033
+ 1.401e+11Hz 0.564581 -0.809417
+ 1.402e+11Hz 0.56402 -0.8098
+ 1.403e+11Hz 0.563457 -0.810183
+ 1.404e+11Hz 0.562895 -0.810565
+ 1.405e+11Hz 0.562332 -0.810948
+ 1.406e+11Hz 0.561768 -0.811329
+ 1.407e+11Hz 0.561205 -0.81171
+ 1.408e+11Hz 0.560641 -0.812091
+ 1.409e+11Hz 0.560077 -0.812471
+ 1.41e+11Hz 0.559512 -0.812851
+ 1.411e+11Hz 0.558947 -0.81323
+ 1.412e+11Hz 0.558382 -0.813609
+ 1.413e+11Hz 0.557817 -0.813987
+ 1.414e+11Hz 0.557251 -0.814365
+ 1.415e+11Hz 0.556685 -0.814742
+ 1.416e+11Hz 0.556118 -0.815119
+ 1.417e+11Hz 0.555552 -0.815496
+ 1.418e+11Hz 0.554985 -0.815872
+ 1.419e+11Hz 0.554418 -0.816247
+ 1.42e+11Hz 0.55385 -0.816622
+ 1.421e+11Hz 0.553282 -0.816997
+ 1.422e+11Hz 0.552714 -0.817371
+ 1.423e+11Hz 0.552145 -0.817744
+ 1.424e+11Hz 0.551577 -0.818117
+ 1.425e+11Hz 0.551008 -0.81849
+ 1.426e+11Hz 0.550439 -0.818862
+ 1.427e+11Hz 0.549869 -0.819233
+ 1.428e+11Hz 0.549299 -0.819605
+ 1.429e+11Hz 0.548729 -0.819975
+ 1.43e+11Hz 0.548159 -0.820345
+ 1.431e+11Hz 0.547588 -0.820715
+ 1.432e+11Hz 0.547017 -0.821084
+ 1.433e+11Hz 0.546446 -0.821453
+ 1.434e+11Hz 0.545875 -0.821821
+ 1.435e+11Hz 0.545303 -0.822188
+ 1.436e+11Hz 0.544731 -0.822555
+ 1.437e+11Hz 0.544159 -0.822922
+ 1.438e+11Hz 0.543587 -0.823288
+ 1.439e+11Hz 0.543014 -0.823654
+ 1.44e+11Hz 0.542441 -0.824019
+ 1.441e+11Hz 0.541868 -0.824384
+ 1.442e+11Hz 0.541295 -0.824748
+ 1.443e+11Hz 0.540721 -0.825111
+ 1.444e+11Hz 0.540147 -0.825474
+ 1.445e+11Hz 0.539573 -0.825837
+ 1.446e+11Hz 0.538999 -0.826199
+ 1.447e+11Hz 0.538425 -0.826561
+ 1.448e+11Hz 0.53785 -0.826922
+ 1.449e+11Hz 0.537275 -0.827283
+ 1.45e+11Hz 0.5367 -0.827643
+ 1.451e+11Hz 0.536125 -0.828002
+ 1.452e+11Hz 0.535549 -0.828362
+ 1.453e+11Hz 0.534974 -0.82872
+ 1.454e+11Hz 0.534398 -0.829079
+ 1.455e+11Hz 0.533822 -0.829436
+ 1.456e+11Hz 0.533246 -0.829793
+ 1.457e+11Hz 0.532669 -0.83015
+ 1.458e+11Hz 0.532092 -0.830506
+ 1.459e+11Hz 0.531516 -0.830862
+ 1.46e+11Hz 0.530939 -0.831217
+ 1.461e+11Hz 0.530362 -0.831572
+ 1.462e+11Hz 0.529784 -0.831927
+ 1.463e+11Hz 0.529207 -0.83228
+ 1.464e+11Hz 0.528629 -0.832634
+ 1.465e+11Hz 0.528051 -0.832987
+ 1.466e+11Hz 0.527473 -0.833339
+ 1.467e+11Hz 0.526895 -0.833691
+ 1.468e+11Hz 0.526317 -0.834042
+ 1.469e+11Hz 0.525738 -0.834393
+ 1.47e+11Hz 0.52516 -0.834744
+ 1.471e+11Hz 0.524581 -0.835094
+ 1.472e+11Hz 0.524002 -0.835444
+ 1.473e+11Hz 0.523423 -0.835793
+ 1.474e+11Hz 0.522844 -0.836142
+ 1.475e+11Hz 0.522265 -0.83649
+ 1.476e+11Hz 0.521686 -0.836838
+ 1.477e+11Hz 0.521106 -0.837185
+ 1.478e+11Hz 0.520526 -0.837532
+ 1.479e+11Hz 0.519946 -0.837879
+ 1.48e+11Hz 0.519366 -0.838225
+ 1.481e+11Hz 0.518786 -0.83857
+ 1.482e+11Hz 0.518206 -0.838916
+ 1.483e+11Hz 0.517626 -0.83926
+ 1.484e+11Hz 0.517045 -0.839605
+ 1.485e+11Hz 0.516465 -0.839949
+ 1.486e+11Hz 0.515884 -0.840292
+ 1.487e+11Hz 0.515303 -0.840635
+ 1.488e+11Hz 0.514722 -0.840978
+ 1.489e+11Hz 0.514141 -0.84132
+ 1.49e+11Hz 0.51356 -0.841662
+ 1.491e+11Hz 0.512979 -0.842004
+ 1.492e+11Hz 0.512398 -0.842345
+ 1.493e+11Hz 0.511816 -0.842686
+ 1.494e+11Hz 0.511235 -0.843026
+ 1.495e+11Hz 0.510653 -0.843366
+ 1.496e+11Hz 0.510071 -0.843706
+ 1.497e+11Hz 0.509489 -0.844045
+ 1.498e+11Hz 0.508907 -0.844384
+ 1.499e+11Hz 0.508325 -0.844723
+ 1.5e+11Hz 0.507743 -0.845061
+ ]

A22 %vd(20 3) %vd(22, 3) xfer4
.model xfer4 xfer R_I=true table=[
+ 0Hz 0.00394946 0
+ 1e+08Hz 0.00394959 -4.21995e-05
+ 2e+08Hz 0.00394996 -8.44065e-05
+ 3e+08Hz 0.00395057 -0.000126629
+ 4e+08Hz 0.00395144 -0.000168874
+ 5e+08Hz 0.00395255 -0.000211149
+ 6e+08Hz 0.0039539 -0.000253463
+ 7e+08Hz 0.0039555 -0.000295821
+ 8e+08Hz 0.00395734 -0.000338233
+ 9e+08Hz 0.00395942 -0.000380706
+ 1e+09Hz 0.00396174 -0.000423246
+ 1.1e+09Hz 0.0039643 -0.000465861
+ 1.2e+09Hz 0.00396709 -0.000508559
+ 1.3e+09Hz 0.00397012 -0.000551347
+ 1.4e+09Hz 0.00397338 -0.000594232
+ 1.5e+09Hz 0.00397687 -0.000637221
+ 1.6e+09Hz 0.00398058 -0.000680322
+ 1.7e+09Hz 0.00398452 -0.000723541
+ 1.8e+09Hz 0.00398868 -0.000766885
+ 1.9e+09Hz 0.00399306 -0.000810362
+ 2e+09Hz 0.00399765 -0.000853978
+ 2.1e+09Hz 0.00400245 -0.000897739
+ 2.2e+09Hz 0.00400746 -0.000941654
+ 2.3e+09Hz 0.00401268 -0.000985726
+ 2.4e+09Hz 0.00401809 -0.00102997
+ 2.5e+09Hz 0.0040237 -0.00107437
+ 2.6e+09Hz 0.0040295 -0.00111896
+ 2.7e+09Hz 0.00403548 -0.00116373
+ 2.8e+09Hz 0.00404165 -0.0012087
+ 2.9e+09Hz 0.004048 -0.00125385
+ 3e+09Hz 0.00405452 -0.00129921
+ 3.1e+09Hz 0.0040612 -0.00134478
+ 3.2e+09Hz 0.00406805 -0.00139056
+ 3.3e+09Hz 0.00407506 -0.00143656
+ 3.4e+09Hz 0.00408223 -0.00148278
+ 3.5e+09Hz 0.00408953 -0.00152922
+ 3.6e+09Hz 0.00409698 -0.00157591
+ 3.7e+09Hz 0.00410457 -0.00162283
+ 3.8e+09Hz 0.00411229 -0.00166999
+ 3.9e+09Hz 0.00412013 -0.0017174
+ 4e+09Hz 0.00412809 -0.00176507
+ 4.1e+09Hz 0.00413617 -0.00181299
+ 4.2e+09Hz 0.00414435 -0.00186117
+ 4.3e+09Hz 0.00415263 -0.00190961
+ 4.4e+09Hz 0.004161 -0.00195832
+ 4.5e+09Hz 0.00416947 -0.00200731
+ 4.6e+09Hz 0.00417801 -0.00205657
+ 4.7e+09Hz 0.00418663 -0.00210611
+ 4.8e+09Hz 0.00419532 -0.00215592
+ 4.9e+09Hz 0.00420407 -0.00220603
+ 5e+09Hz 0.00421288 -0.00225642
+ 5.1e+09Hz 0.00422174 -0.0023071
+ 5.2e+09Hz 0.00423063 -0.00235808
+ 5.3e+09Hz 0.00423957 -0.00240935
+ 5.4e+09Hz 0.00424853 -0.00246091
+ 5.5e+09Hz 0.00425751 -0.00251278
+ 5.6e+09Hz 0.00426651 -0.00256495
+ 5.7e+09Hz 0.00427552 -0.00261742
+ 5.8e+09Hz 0.00428453 -0.0026702
+ 5.9e+09Hz 0.00429353 -0.00272328
+ 6e+09Hz 0.00430252 -0.00277667
+ 6.1e+09Hz 0.00431149 -0.00283036
+ 6.2e+09Hz 0.00432043 -0.00288437
+ 6.3e+09Hz 0.00432934 -0.00293868
+ 6.4e+09Hz 0.00433821 -0.00299331
+ 6.5e+09Hz 0.00434703 -0.00304825
+ 6.6e+09Hz 0.0043558 -0.0031035
+ 6.7e+09Hz 0.00436451 -0.00315906
+ 6.8e+09Hz 0.00437315 -0.00321493
+ 6.9e+09Hz 0.00438171 -0.00327111
+ 7e+09Hz 0.0043902 -0.00332761
+ 7.1e+09Hz 0.00439859 -0.00338441
+ 7.2e+09Hz 0.00440689 -0.00344152
+ 7.3e+09Hz 0.00441509 -0.00349894
+ 7.4e+09Hz 0.00442318 -0.00355668
+ 7.5e+09Hz 0.00443115 -0.00361471
+ 7.6e+09Hz 0.00443901 -0.00367306
+ 7.7e+09Hz 0.00444673 -0.0037317
+ 7.8e+09Hz 0.00445432 -0.00379065
+ 7.9e+09Hz 0.00446177 -0.0038499
+ 8e+09Hz 0.00446908 -0.00390945
+ 8.1e+09Hz 0.00447623 -0.0039693
+ 8.2e+09Hz 0.00448322 -0.00402944
+ 8.3e+09Hz 0.00449004 -0.00408988
+ 8.4e+09Hz 0.0044967 -0.00415061
+ 8.5e+09Hz 0.00450317 -0.00421163
+ 8.6e+09Hz 0.00450947 -0.00427293
+ 8.7e+09Hz 0.00451557 -0.00433451
+ 8.8e+09Hz 0.00452148 -0.00439638
+ 8.9e+09Hz 0.00452719 -0.00445852
+ 9e+09Hz 0.00453269 -0.00452094
+ 9.1e+09Hz 0.00453798 -0.00458364
+ 9.2e+09Hz 0.00454305 -0.0046466
+ 9.3e+09Hz 0.0045479 -0.00470982
+ 9.4e+09Hz 0.00455253 -0.00477331
+ 9.5e+09Hz 0.00455692 -0.00483705
+ 9.6e+09Hz 0.00456107 -0.00490106
+ 9.7e+09Hz 0.00456499 -0.00496531
+ 9.8e+09Hz 0.00456865 -0.00502981
+ 9.9e+09Hz 0.00457207 -0.00509455
+ 1e+10Hz 0.00457522 -0.00515954
+ 1.01e+10Hz 0.00457812 -0.00522476
+ 1.02e+10Hz 0.00458076 -0.00529021
+ 1.03e+10Hz 0.00458312 -0.00535589
+ 1.04e+10Hz 0.00458521 -0.0054218
+ 1.05e+10Hz 0.00458702 -0.00548792
+ 1.06e+10Hz 0.00458856 -0.00555426
+ 1.07e+10Hz 0.00458981 -0.00562081
+ 1.08e+10Hz 0.00459077 -0.00568757
+ 1.09e+10Hz 0.00459143 -0.00575452
+ 1.1e+10Hz 0.00459181 -0.00582168
+ 1.11e+10Hz 0.00459188 -0.00588903
+ 1.12e+10Hz 0.00459165 -0.00595657
+ 1.13e+10Hz 0.00459112 -0.00602429
+ 1.14e+10Hz 0.00459028 -0.00609219
+ 1.15e+10Hz 0.00458913 -0.00616026
+ 1.16e+10Hz 0.00458766 -0.00622851
+ 1.17e+10Hz 0.00458588 -0.00629692
+ 1.18e+10Hz 0.00458378 -0.00636549
+ 1.19e+10Hz 0.00458136 -0.00643421
+ 1.2e+10Hz 0.00457862 -0.00650309
+ 1.21e+10Hz 0.00457555 -0.00657211
+ 1.22e+10Hz 0.00457215 -0.00664127
+ 1.23e+10Hz 0.00456843 -0.00671057
+ 1.24e+10Hz 0.00456437 -0.00678
+ 1.25e+10Hz 0.00455998 -0.00684956
+ 1.26e+10Hz 0.00455526 -0.00691924
+ 1.27e+10Hz 0.0045502 -0.00698903
+ 1.28e+10Hz 0.0045448 -0.00705893
+ 1.29e+10Hz 0.00453907 -0.00712895
+ 1.3e+10Hz 0.00453299 -0.00719906
+ 1.31e+10Hz 0.00452657 -0.00726927
+ 1.32e+10Hz 0.00451982 -0.00733958
+ 1.33e+10Hz 0.00451272 -0.00740997
+ 1.34e+10Hz 0.00450528 -0.00748044
+ 1.35e+10Hz 0.00449749 -0.00755099
+ 1.36e+10Hz 0.00448936 -0.00762162
+ 1.37e+10Hz 0.00448088 -0.00769231
+ 1.38e+10Hz 0.00447206 -0.00776307
+ 1.39e+10Hz 0.00446289 -0.00783388
+ 1.4e+10Hz 0.00445338 -0.00790475
+ 1.41e+10Hz 0.00444353 -0.00797567
+ 1.42e+10Hz 0.00443333 -0.00804664
+ 1.43e+10Hz 0.00442278 -0.00811764
+ 1.44e+10Hz 0.00441189 -0.00818869
+ 1.45e+10Hz 0.00440065 -0.00825976
+ 1.46e+10Hz 0.00438907 -0.00833086
+ 1.47e+10Hz 0.00437714 -0.00840198
+ 1.48e+10Hz 0.00436488 -0.00847312
+ 1.49e+10Hz 0.00435227 -0.00854428
+ 1.5e+10Hz 0.00433932 -0.00861544
+ 1.51e+10Hz 0.00432602 -0.00868662
+ 1.52e+10Hz 0.00431239 -0.00875779
+ 1.53e+10Hz 0.00429842 -0.00882896
+ 1.54e+10Hz 0.00428412 -0.00890012
+ 1.55e+10Hz 0.00426947 -0.00897128
+ 1.56e+10Hz 0.00425449 -0.00904241
+ 1.57e+10Hz 0.00423918 -0.00911353
+ 1.58e+10Hz 0.00422353 -0.00918463
+ 1.59e+10Hz 0.00420755 -0.0092557
+ 1.6e+10Hz 0.00419125 -0.00932674
+ 1.61e+10Hz 0.00417461 -0.00939775
+ 1.62e+10Hz 0.00415765 -0.00946872
+ 1.63e+10Hz 0.00414036 -0.00953965
+ 1.64e+10Hz 0.00412275 -0.00961054
+ 1.65e+10Hz 0.00410482 -0.00968138
+ 1.66e+10Hz 0.00408657 -0.00975217
+ 1.67e+10Hz 0.004068 -0.00982291
+ 1.68e+10Hz 0.00404912 -0.00989358
+ 1.69e+10Hz 0.00402992 -0.0099642
+ 1.7e+10Hz 0.00401041 -0.0100348
+ 1.71e+10Hz 0.00399059 -0.0101052
+ 1.72e+10Hz 0.00397046 -0.0101757
+ 1.73e+10Hz 0.00395003 -0.010246
+ 1.74e+10Hz 0.00392929 -0.0103163
+ 1.75e+10Hz 0.00390826 -0.0103865
+ 1.76e+10Hz 0.00388692 -0.0104566
+ 1.77e+10Hz 0.00386529 -0.0105266
+ 1.78e+10Hz 0.00384336 -0.0105966
+ 1.79e+10Hz 0.00382114 -0.0106664
+ 1.8e+10Hz 0.00379863 -0.0107362
+ 1.81e+10Hz 0.00377584 -0.0108059
+ 1.82e+10Hz 0.00375276 -0.0108755
+ 1.83e+10Hz 0.00372939 -0.0109449
+ 1.84e+10Hz 0.00370575 -0.0110143
+ 1.85e+10Hz 0.00368183 -0.0110836
+ 1.86e+10Hz 0.00365764 -0.0111528
+ 1.87e+10Hz 0.00363317 -0.0112219
+ 1.88e+10Hz 0.00360843 -0.0112908
+ 1.89e+10Hz 0.00358343 -0.0113597
+ 1.9e+10Hz 0.00355816 -0.0114284
+ 1.91e+10Hz 0.00353263 -0.0114971
+ 1.92e+10Hz 0.00350684 -0.0115656
+ 1.93e+10Hz 0.00348079 -0.011634
+ 1.94e+10Hz 0.00345449 -0.0117023
+ 1.95e+10Hz 0.00342793 -0.0117705
+ 1.96e+10Hz 0.00340113 -0.0118386
+ 1.97e+10Hz 0.00337407 -0.0119065
+ 1.98e+10Hz 0.00334678 -0.0119743
+ 1.99e+10Hz 0.00331924 -0.012042
+ 2e+10Hz 0.00329146 -0.0121096
+ 2.01e+10Hz 0.00326345 -0.0121771
+ 2.02e+10Hz 0.0032352 -0.0122444
+ 2.03e+10Hz 0.00320672 -0.0123116
+ 2.04e+10Hz 0.00317801 -0.0123786
+ 2.05e+10Hz 0.00314907 -0.0124456
+ 2.06e+10Hz 0.00311991 -0.0125124
+ 2.07e+10Hz 0.00309053 -0.0125791
+ 2.08e+10Hz 0.00306092 -0.0126457
+ 2.09e+10Hz 0.0030311 -0.0127121
+ 2.1e+10Hz 0.00300107 -0.0127784
+ 2.11e+10Hz 0.00297082 -0.0128445
+ 2.12e+10Hz 0.00294036 -0.0129106
+ 2.13e+10Hz 0.0029097 -0.0129765
+ 2.14e+10Hz 0.00287883 -0.0130423
+ 2.15e+10Hz 0.00284776 -0.0131079
+ 2.16e+10Hz 0.00281649 -0.0131734
+ 2.17e+10Hz 0.00278501 -0.0132388
+ 2.18e+10Hz 0.00275334 -0.013304
+ 2.19e+10Hz 0.00272148 -0.0133692
+ 2.2e+10Hz 0.00268943 -0.0134341
+ 2.21e+10Hz 0.00265718 -0.013499
+ 2.22e+10Hz 0.00262475 -0.0135637
+ 2.23e+10Hz 0.00259214 -0.0136283
+ 2.24e+10Hz 0.00255933 -0.0136928
+ 2.25e+10Hz 0.00252635 -0.0137571
+ 2.26e+10Hz 0.00249319 -0.0138213
+ 2.27e+10Hz 0.00245985 -0.0138853
+ 2.28e+10Hz 0.00242633 -0.0139493
+ 2.29e+10Hz 0.00239265 -0.0140131
+ 2.3e+10Hz 0.00235878 -0.0140768
+ 2.31e+10Hz 0.00232475 -0.0141403
+ 2.32e+10Hz 0.00229055 -0.0142037
+ 2.33e+10Hz 0.00225619 -0.014267
+ 2.34e+10Hz 0.00222165 -0.0143302
+ 2.35e+10Hz 0.00218696 -0.0143932
+ 2.36e+10Hz 0.0021521 -0.0144561
+ 2.37e+10Hz 0.00211708 -0.0145189
+ 2.38e+10Hz 0.00208191 -0.0145816
+ 2.39e+10Hz 0.00204658 -0.0146441
+ 2.4e+10Hz 0.00201109 -0.0147065
+ 2.41e+10Hz 0.00197545 -0.0147688
+ 2.42e+10Hz 0.00193965 -0.014831
+ 2.43e+10Hz 0.0019037 -0.014893
+ 2.44e+10Hz 0.00186761 -0.0149549
+ 2.45e+10Hz 0.00183136 -0.0150167
+ 2.46e+10Hz 0.00179496 -0.0150784
+ 2.47e+10Hz 0.00175843 -0.01514
+ 2.48e+10Hz 0.00172174 -0.0152014
+ 2.49e+10Hz 0.00168491 -0.0152628
+ 2.5e+10Hz 0.00164794 -0.015324
+ 2.51e+10Hz 0.00161082 -0.0153851
+ 2.52e+10Hz 0.00157357 -0.0154461
+ 2.53e+10Hz 0.00153617 -0.015507
+ 2.54e+10Hz 0.00149864 -0.0155677
+ 2.55e+10Hz 0.00146097 -0.0156284
+ 2.56e+10Hz 0.00142315 -0.0156889
+ 2.57e+10Hz 0.00138521 -0.0157493
+ 2.58e+10Hz 0.00134713 -0.0158097
+ 2.59e+10Hz 0.00130891 -0.0158699
+ 2.6e+10Hz 0.00127056 -0.01593
+ 2.61e+10Hz 0.00123207 -0.01599
+ 2.62e+10Hz 0.00119345 -0.0160499
+ 2.63e+10Hz 0.0011547 -0.0161097
+ 2.64e+10Hz 0.00111582 -0.0161694
+ 2.65e+10Hz 0.00107681 -0.016229
+ 2.66e+10Hz 0.00103766 -0.0162885
+ 2.67e+10Hz 0.000998389 -0.0163479
+ 2.68e+10Hz 0.000958984 -0.0164072
+ 2.69e+10Hz 0.00091945 -0.0164664
+ 2.7e+10Hz 0.000879787 -0.0165255
+ 2.71e+10Hz 0.000839995 -0.0165845
+ 2.72e+10Hz 0.000800075 -0.0166434
+ 2.73e+10Hz 0.000760026 -0.0167022
+ 2.74e+10Hz 0.000719849 -0.0167609
+ 2.75e+10Hz 0.000679545 -0.0168195
+ 2.76e+10Hz 0.000639113 -0.016878
+ 2.77e+10Hz 0.000598553 -0.0169365
+ 2.78e+10Hz 0.000557866 -0.0169948
+ 2.79e+10Hz 0.000517052 -0.0170531
+ 2.8e+10Hz 0.000476111 -0.0171112
+ 2.81e+10Hz 0.000435042 -0.0171693
+ 2.82e+10Hz 0.000393847 -0.0172273
+ 2.83e+10Hz 0.000352524 -0.0172852
+ 2.84e+10Hz 0.000311073 -0.017343
+ 2.85e+10Hz 0.000269496 -0.0174008
+ 2.86e+10Hz 0.000227791 -0.0174584
+ 2.87e+10Hz 0.000185959 -0.017516
+ 2.88e+10Hz 0.000143999 -0.0175735
+ 2.89e+10Hz 0.000101911 -0.0176308
+ 2.9e+10Hz 5.96952e-05 -0.0176881
+ 2.91e+10Hz 1.73513e-05 -0.0177454
+ 2.92e+10Hz -2.51211e-05 -0.0178025
+ 2.93e+10Hz -6.77221e-05 -0.0178596
+ 2.94e+10Hz -0.000110452 -0.0179166
+ 2.95e+10Hz -0.000153311 -0.0179735
+ 2.96e+10Hz -0.0001963 -0.0180303
+ 2.97e+10Hz -0.000239418 -0.0180871
+ 2.98e+10Hz -0.000282667 -0.0181438
+ 2.99e+10Hz -0.000326046 -0.0182004
+ 3e+10Hz -0.000369555 -0.0182569
+ 3.01e+10Hz -0.000413196 -0.0183133
+ 3.02e+10Hz -0.000456969 -0.0183697
+ 3.03e+10Hz -0.000500874 -0.018426
+ 3.04e+10Hz -0.00054491 -0.0184822
+ 3.05e+10Hz -0.00058908 -0.0185383
+ 3.06e+10Hz -0.000633383 -0.0185944
+ 3.07e+10Hz -0.00067782 -0.0186503
+ 3.08e+10Hz -0.000722391 -0.0187063
+ 3.09e+10Hz -0.000767096 -0.0187621
+ 3.1e+10Hz -0.000811936 -0.0188179
+ 3.11e+10Hz -0.000856912 -0.0188735
+ 3.12e+10Hz -0.000902024 -0.0189291
+ 3.13e+10Hz -0.000947273 -0.0189847
+ 3.14e+10Hz -0.000992658 -0.0190401
+ 3.15e+10Hz -0.00103818 -0.0190955
+ 3.16e+10Hz -0.00108384 -0.0191508
+ 3.17e+10Hz -0.00112964 -0.0192061
+ 3.18e+10Hz -0.00117558 -0.0192613
+ 3.19e+10Hz -0.00122166 -0.0193163
+ 3.2e+10Hz -0.00126788 -0.0193713
+ 3.21e+10Hz -0.00131423 -0.0194263
+ 3.22e+10Hz -0.00136073 -0.0194812
+ 3.23e+10Hz -0.00140737 -0.019536
+ 3.24e+10Hz -0.00145416 -0.0195907
+ 3.25e+10Hz -0.00150108 -0.0196453
+ 3.26e+10Hz -0.00154815 -0.0196999
+ 3.27e+10Hz -0.00159537 -0.0197544
+ 3.28e+10Hz -0.00164272 -0.0198088
+ 3.29e+10Hz -0.00169022 -0.0198631
+ 3.3e+10Hz -0.00173787 -0.0199174
+ 3.31e+10Hz -0.00178566 -0.0199716
+ 3.32e+10Hz -0.0018336 -0.0200257
+ 3.33e+10Hz -0.00188168 -0.0200798
+ 3.34e+10Hz -0.00192992 -0.0201337
+ 3.35e+10Hz -0.0019783 -0.0201876
+ 3.36e+10Hz -0.00202682 -0.0202414
+ 3.37e+10Hz -0.0020755 -0.0202952
+ 3.38e+10Hz -0.00212432 -0.0203488
+ 3.39e+10Hz -0.0021733 -0.0204024
+ 3.4e+10Hz -0.00222242 -0.0204559
+ 3.41e+10Hz -0.00227169 -0.0205093
+ 3.42e+10Hz -0.00232112 -0.0205626
+ 3.43e+10Hz -0.00237069 -0.0206159
+ 3.44e+10Hz -0.00242042 -0.020669
+ 3.45e+10Hz -0.0024703 -0.0207221
+ 3.46e+10Hz -0.00252033 -0.0207751
+ 3.47e+10Hz -0.00257052 -0.020828
+ 3.48e+10Hz -0.00262085 -0.0208809
+ 3.49e+10Hz -0.00267134 -0.0209336
+ 3.5e+10Hz -0.00272198 -0.0209863
+ 3.51e+10Hz -0.00277278 -0.0210389
+ 3.52e+10Hz -0.00282373 -0.0210914
+ 3.53e+10Hz -0.00287484 -0.0211438
+ 3.54e+10Hz -0.0029261 -0.0211961
+ 3.55e+10Hz -0.00297752 -0.0212483
+ 3.56e+10Hz -0.00302908 -0.0213005
+ 3.57e+10Hz -0.00308081 -0.0213526
+ 3.58e+10Hz -0.00313269 -0.0214045
+ 3.59e+10Hz -0.00318473 -0.0214564
+ 3.6e+10Hz -0.00323693 -0.0215082
+ 3.61e+10Hz -0.00328928 -0.0215599
+ 3.62e+10Hz -0.00334178 -0.0216115
+ 3.63e+10Hz -0.00339445 -0.021663
+ 3.64e+10Hz -0.00344727 -0.0217144
+ 3.65e+10Hz -0.00350025 -0.0217657
+ 3.66e+10Hz -0.00355338 -0.0218169
+ 3.67e+10Hz -0.00360667 -0.021868
+ 3.68e+10Hz -0.00366012 -0.0219191
+ 3.69e+10Hz -0.00371373 -0.02197
+ 3.7e+10Hz -0.00376749 -0.0220208
+ 3.71e+10Hz -0.00382141 -0.0220715
+ 3.72e+10Hz -0.00387549 -0.0221222
+ 3.73e+10Hz -0.00392973 -0.0221727
+ 3.74e+10Hz -0.00398412 -0.0222231
+ 3.75e+10Hz -0.00403867 -0.0222735
+ 3.76e+10Hz -0.00409338 -0.0223237
+ 3.77e+10Hz -0.00414824 -0.0223738
+ 3.78e+10Hz -0.00420326 -0.0224238
+ 3.79e+10Hz -0.00425844 -0.0224737
+ 3.8e+10Hz -0.00431378 -0.0225235
+ 3.81e+10Hz -0.00436927 -0.0225732
+ 3.82e+10Hz -0.00442492 -0.0226227
+ 3.83e+10Hz -0.00448073 -0.0226722
+ 3.84e+10Hz -0.00453669 -0.0227216
+ 3.85e+10Hz -0.00459281 -0.0227708
+ 3.86e+10Hz -0.00464908 -0.0228199
+ 3.87e+10Hz -0.00470552 -0.0228689
+ 3.88e+10Hz -0.0047621 -0.0229178
+ 3.89e+10Hz -0.00481884 -0.0229666
+ 3.9e+10Hz -0.00487574 -0.0230153
+ 3.91e+10Hz -0.00493279 -0.0230639
+ 3.92e+10Hz -0.00499 -0.0231123
+ 3.93e+10Hz -0.00504736 -0.0231606
+ 3.94e+10Hz -0.00510487 -0.0232088
+ 3.95e+10Hz -0.00516254 -0.0232569
+ 3.96e+10Hz -0.00522036 -0.0233049
+ 3.97e+10Hz -0.00527834 -0.0233527
+ 3.98e+10Hz -0.00533646 -0.0234004
+ 3.99e+10Hz -0.00539474 -0.023448
+ 4e+10Hz -0.00545317 -0.0234955
+ 4.01e+10Hz -0.00551175 -0.0235429
+ 4.02e+10Hz -0.00557049 -0.0235901
+ 4.03e+10Hz -0.00562937 -0.0236372
+ 4.04e+10Hz -0.0056884 -0.0236842
+ 4.05e+10Hz -0.00574759 -0.023731
+ 4.06e+10Hz -0.00580692 -0.0237777
+ 4.07e+10Hz -0.0058664 -0.0238243
+ 4.08e+10Hz -0.00592603 -0.0238708
+ 4.09e+10Hz -0.00598581 -0.0239171
+ 4.1e+10Hz -0.00604573 -0.0239633
+ 4.11e+10Hz -0.0061058 -0.0240094
+ 4.12e+10Hz -0.00616602 -0.0240553
+ 4.13e+10Hz -0.00622638 -0.0241011
+ 4.14e+10Hz -0.00628689 -0.0241468
+ 4.15e+10Hz -0.00634754 -0.0241923
+ 4.16e+10Hz -0.00640834 -0.0242377
+ 4.17e+10Hz -0.00646928 -0.024283
+ 4.18e+10Hz -0.00653036 -0.0243281
+ 4.19e+10Hz -0.00659158 -0.0243731
+ 4.2e+10Hz -0.00665295 -0.024418
+ 4.21e+10Hz -0.00671446 -0.0244627
+ 4.22e+10Hz -0.00677611 -0.0245073
+ 4.23e+10Hz -0.00683789 -0.0245517
+ 4.24e+10Hz -0.00689982 -0.024596
+ 4.25e+10Hz -0.00696189 -0.0246402
+ 4.26e+10Hz -0.00702409 -0.0246842
+ 4.27e+10Hz -0.00708643 -0.0247281
+ 4.28e+10Hz -0.00714891 -0.0247718
+ 4.29e+10Hz -0.00721152 -0.0248154
+ 4.3e+10Hz -0.00727427 -0.0248589
+ 4.31e+10Hz -0.00733715 -0.0249022
+ 4.32e+10Hz -0.00740017 -0.0249454
+ 4.33e+10Hz -0.00746332 -0.0249884
+ 4.34e+10Hz -0.00752661 -0.0250313
+ 4.35e+10Hz -0.00759002 -0.025074
+ 4.36e+10Hz -0.00765357 -0.0251166
+ 4.37e+10Hz -0.00771725 -0.025159
+ 4.38e+10Hz -0.00778106 -0.0252013
+ 4.39e+10Hz -0.00784499 -0.0252435
+ 4.4e+10Hz -0.00790906 -0.0252855
+ 4.41e+10Hz -0.00797325 -0.0253273
+ 4.42e+10Hz -0.00803757 -0.0253691
+ 4.43e+10Hz -0.00810202 -0.0254106
+ 4.44e+10Hz -0.00816659 -0.025452
+ 4.45e+10Hz -0.00823129 -0.0254933
+ 4.46e+10Hz -0.00829611 -0.0255344
+ 4.47e+10Hz -0.00836106 -0.0255754
+ 4.48e+10Hz -0.00842613 -0.0256162
+ 4.49e+10Hz -0.00849132 -0.0256569
+ 4.5e+10Hz -0.00855664 -0.0256974
+ 4.51e+10Hz -0.00862207 -0.0257378
+ 4.52e+10Hz -0.00868763 -0.025778
+ 4.53e+10Hz -0.0087533 -0.025818
+ 4.54e+10Hz -0.0088191 -0.025858
+ 4.55e+10Hz -0.00888501 -0.0258977
+ 4.56e+10Hz -0.00895104 -0.0259373
+ 4.57e+10Hz -0.00901719 -0.0259768
+ 4.58e+10Hz -0.00908346 -0.0260161
+ 4.59e+10Hz -0.00914984 -0.0260553
+ 4.6e+10Hz -0.00921633 -0.0260943
+ 4.61e+10Hz -0.00928294 -0.0261331
+ 4.62e+10Hz -0.00934966 -0.0261718
+ 4.63e+10Hz -0.0094165 -0.0262104
+ 4.64e+10Hz -0.00948345 -0.0262488
+ 4.65e+10Hz -0.00955051 -0.026287
+ 4.66e+10Hz -0.00961768 -0.0263251
+ 4.67e+10Hz -0.00968496 -0.0263631
+ 4.68e+10Hz -0.00975235 -0.0264009
+ 4.69e+10Hz -0.00981985 -0.0264385
+ 4.7e+10Hz -0.00988746 -0.026476
+ 4.71e+10Hz -0.00995518 -0.0265133
+ 4.72e+10Hz -0.010023 -0.0265505
+ 4.73e+10Hz -0.0100909 -0.0265875
+ 4.74e+10Hz -0.010159 -0.0266244
+ 4.75e+10Hz -0.0102271 -0.0266611
+ 4.76e+10Hz -0.0102954 -0.0266977
+ 4.77e+10Hz -0.0103637 -0.0267341
+ 4.78e+10Hz -0.0104322 -0.0267703
+ 4.79e+10Hz -0.0105007 -0.0268064
+ 4.8e+10Hz -0.0105694 -0.0268424
+ 4.81e+10Hz -0.0106382 -0.0268782
+ 4.82e+10Hz -0.010707 -0.0269138
+ 4.83e+10Hz -0.010776 -0.0269493
+ 4.84e+10Hz -0.0108451 -0.0269847
+ 4.85e+10Hz -0.0109143 -0.0270198
+ 4.86e+10Hz -0.0109835 -0.0270549
+ 4.87e+10Hz -0.0110529 -0.0270898
+ 4.88e+10Hz -0.0111224 -0.0271245
+ 4.89e+10Hz -0.011192 -0.0271591
+ 4.9e+10Hz -0.0112616 -0.0271935
+ 4.91e+10Hz -0.0113314 -0.0272277
+ 4.92e+10Hz -0.0114012 -0.0272619
+ 4.93e+10Hz -0.0114712 -0.0272958
+ 4.94e+10Hz -0.0115412 -0.0273296
+ 4.95e+10Hz -0.0116114 -0.0273633
+ 4.96e+10Hz -0.0116817 -0.0273968
+ 4.97e+10Hz -0.011752 -0.0274302
+ 4.98e+10Hz -0.0118224 -0.0274634
+ 4.99e+10Hz -0.0118929 -0.0274964
+ 5e+10Hz -0.0119636 -0.0275293
+ 5.01e+10Hz -0.0120343 -0.0275621
+ 5.02e+10Hz -0.0121051 -0.0275946
+ 5.03e+10Hz -0.012176 -0.0276271
+ 5.04e+10Hz -0.012247 -0.0276594
+ 5.05e+10Hz -0.0123181 -0.0276915
+ 5.06e+10Hz -0.0123893 -0.0277235
+ 5.07e+10Hz -0.0124605 -0.0277554
+ 5.08e+10Hz -0.0125319 -0.027787
+ 5.09e+10Hz -0.0126033 -0.0278186
+ 5.1e+10Hz -0.0126749 -0.0278499
+ 5.11e+10Hz -0.0127465 -0.0278812
+ 5.12e+10Hz -0.0128182 -0.0279123
+ 5.13e+10Hz -0.0128901 -0.0279432
+ 5.14e+10Hz -0.012962 -0.027974
+ 5.15e+10Hz -0.013034 -0.0280046
+ 5.16e+10Hz -0.013106 -0.0280351
+ 5.17e+10Hz -0.0131782 -0.0280654
+ 5.18e+10Hz -0.0132505 -0.0280956
+ 5.19e+10Hz -0.0133228 -0.0281256
+ 5.2e+10Hz -0.0133952 -0.0281555
+ 5.21e+10Hz -0.0134677 -0.0281852
+ 5.22e+10Hz -0.0135403 -0.0282148
+ 5.23e+10Hz -0.013613 -0.0282442
+ 5.24e+10Hz -0.0136858 -0.0282735
+ 5.25e+10Hz -0.0137587 -0.0283026
+ 5.26e+10Hz -0.0138316 -0.0283316
+ 5.27e+10Hz -0.0139047 -0.0283604
+ 5.28e+10Hz -0.0139778 -0.0283891
+ 5.29e+10Hz -0.014051 -0.0284177
+ 5.3e+10Hz -0.0141243 -0.028446
+ 5.31e+10Hz -0.0141977 -0.0284743
+ 5.32e+10Hz -0.0142712 -0.0285023
+ 5.33e+10Hz -0.0143448 -0.0285303
+ 5.34e+10Hz -0.0144184 -0.0285581
+ 5.35e+10Hz -0.0144921 -0.0285857
+ 5.36e+10Hz -0.0145659 -0.0286132
+ 5.37e+10Hz -0.0146398 -0.0286405
+ 5.38e+10Hz -0.0147138 -0.0286677
+ 5.39e+10Hz -0.0147879 -0.0286947
+ 5.4e+10Hz -0.0148621 -0.0287216
+ 5.41e+10Hz -0.0149363 -0.0287484
+ 5.42e+10Hz -0.0150106 -0.028775
+ 5.43e+10Hz -0.015085 -0.0288014
+ 5.44e+10Hz -0.0151595 -0.0288277
+ 5.45e+10Hz -0.0152341 -0.0288538
+ 5.46e+10Hz -0.0153088 -0.0288798
+ 5.47e+10Hz -0.0153835 -0.0289057
+ 5.48e+10Hz -0.0154584 -0.0289313
+ 5.49e+10Hz -0.0155333 -0.0289569
+ 5.5e+10Hz -0.0156083 -0.0289823
+ 5.51e+10Hz -0.0156834 -0.0290075
+ 5.52e+10Hz -0.0157585 -0.0290326
+ 5.53e+10Hz -0.0158338 -0.0290575
+ 5.54e+10Hz -0.0159091 -0.0290823
+ 5.55e+10Hz -0.0159846 -0.029107
+ 5.56e+10Hz -0.0160601 -0.0291315
+ 5.57e+10Hz -0.0161357 -0.0291558
+ 5.58e+10Hz -0.0162113 -0.02918
+ 5.59e+10Hz -0.0162871 -0.029204
+ 5.6e+10Hz -0.0163629 -0.0292279
+ 5.61e+10Hz -0.0164389 -0.0292517
+ 5.62e+10Hz -0.0165149 -0.0292752
+ 5.63e+10Hz -0.016591 -0.0292987
+ 5.64e+10Hz -0.0166671 -0.029322
+ 5.65e+10Hz -0.0167434 -0.0293451
+ 5.66e+10Hz -0.0168197 -0.0293681
+ 5.67e+10Hz -0.0168961 -0.0293909
+ 5.68e+10Hz -0.0169727 -0.0294136
+ 5.69e+10Hz -0.0170493 -0.0294361
+ 5.7e+10Hz -0.0171259 -0.0294585
+ 5.71e+10Hz -0.0172027 -0.0294807
+ 5.72e+10Hz -0.0172795 -0.0295028
+ 5.73e+10Hz -0.0173565 -0.0295247
+ 5.74e+10Hz -0.0174335 -0.0295465
+ 5.75e+10Hz -0.0175106 -0.0295681
+ 5.76e+10Hz -0.0175877 -0.0295895
+ 5.77e+10Hz -0.017665 -0.0296108
+ 5.78e+10Hz -0.0177423 -0.029632
+ 5.79e+10Hz -0.0178198 -0.029653
+ 5.8e+10Hz -0.0178973 -0.0296738
+ 5.81e+10Hz -0.0179749 -0.0296945
+ 5.82e+10Hz -0.0180525 -0.029715
+ 5.83e+10Hz -0.0181303 -0.0297354
+ 5.84e+10Hz -0.0182081 -0.0297556
+ 5.85e+10Hz -0.0182861 -0.0297757
+ 5.86e+10Hz -0.0183641 -0.0297956
+ 5.87e+10Hz -0.0184422 -0.0298153
+ 5.88e+10Hz -0.0185203 -0.0298349
+ 5.89e+10Hz -0.0185986 -0.0298543
+ 5.9e+10Hz -0.0186769 -0.0298736
+ 5.91e+10Hz -0.0187553 -0.0298927
+ 5.92e+10Hz -0.0188338 -0.0299117
+ 5.93e+10Hz -0.0189124 -0.0299305
+ 5.94e+10Hz -0.018991 -0.0299491
+ 5.95e+10Hz -0.0190698 -0.0299676
+ 5.96e+10Hz -0.0191486 -0.0299859
+ 5.97e+10Hz -0.0192275 -0.0300041
+ 5.98e+10Hz -0.0193065 -0.0300221
+ 5.99e+10Hz -0.0193856 -0.0300399
+ 6e+10Hz -0.0194647 -0.0300576
+ 6.01e+10Hz -0.019544 -0.0300751
+ 6.02e+10Hz -0.0196233 -0.0300925
+ 6.03e+10Hz -0.0197026 -0.0301097
+ 6.04e+10Hz -0.0197821 -0.0301267
+ 6.05e+10Hz -0.0198617 -0.0301436
+ 6.06e+10Hz -0.0199413 -0.0301603
+ 6.07e+10Hz -0.020021 -0.0301768
+ 6.08e+10Hz -0.0201008 -0.0301932
+ 6.09e+10Hz -0.0201807 -0.0302094
+ 6.1e+10Hz -0.0202606 -0.0302255
+ 6.11e+10Hz -0.0203406 -0.0302413
+ 6.12e+10Hz -0.0204207 -0.0302571
+ 6.13e+10Hz -0.0205009 -0.0302726
+ 6.14e+10Hz -0.0205812 -0.030288
+ 6.15e+10Hz -0.0206615 -0.0303032
+ 6.16e+10Hz -0.0207419 -0.0303183
+ 6.17e+10Hz -0.0208224 -0.0303332
+ 6.18e+10Hz -0.020903 -0.0303479
+ 6.19e+10Hz -0.0209837 -0.0303624
+ 6.2e+10Hz -0.0210644 -0.0303768
+ 6.21e+10Hz -0.0211452 -0.030391
+ 6.22e+10Hz -0.0212261 -0.0304051
+ 6.23e+10Hz -0.021307 -0.030419
+ 6.24e+10Hz -0.0213881 -0.0304326
+ 6.25e+10Hz -0.0214692 -0.0304462
+ 6.26e+10Hz -0.0215503 -0.0304595
+ 6.27e+10Hz -0.0216316 -0.0304727
+ 6.28e+10Hz -0.0217129 -0.0304858
+ 6.29e+10Hz -0.0217944 -0.0304986
+ 6.3e+10Hz -0.0218758 -0.0305113
+ 6.31e+10Hz -0.0219574 -0.0305238
+ 6.32e+10Hz -0.022039 -0.0305361
+ 6.33e+10Hz -0.0221207 -0.0305483
+ 6.34e+10Hz -0.0222025 -0.0305602
+ 6.35e+10Hz -0.0222843 -0.030572
+ 6.36e+10Hz -0.0223662 -0.0305837
+ 6.37e+10Hz -0.0224482 -0.0305951
+ 6.38e+10Hz -0.0225303 -0.0306064
+ 6.39e+10Hz -0.0226124 -0.0306175
+ 6.4e+10Hz -0.0226946 -0.0306285
+ 6.41e+10Hz -0.0227769 -0.0306392
+ 6.42e+10Hz -0.0228592 -0.0306498
+ 6.43e+10Hz -0.0229416 -0.0306602
+ 6.44e+10Hz -0.0230241 -0.0306704
+ 6.45e+10Hz -0.0231066 -0.0306804
+ 6.46e+10Hz -0.0231893 -0.0306903
+ 6.47e+10Hz -0.0232719 -0.0307
+ 6.48e+10Hz -0.0233547 -0.0307095
+ 6.49e+10Hz -0.0234375 -0.0307188
+ 6.5e+10Hz -0.0235204 -0.030728
+ 6.51e+10Hz -0.0236033 -0.0307369
+ 6.52e+10Hz -0.0236863 -0.0307457
+ 6.53e+10Hz -0.0237694 -0.0307543
+ 6.54e+10Hz -0.0238526 -0.0307627
+ 6.55e+10Hz -0.0239358 -0.030771
+ 6.56e+10Hz -0.024019 -0.030779
+ 6.57e+10Hz -0.0241024 -0.0307869
+ 6.58e+10Hz -0.0241858 -0.0307946
+ 6.59e+10Hz -0.0242692 -0.0308021
+ 6.6e+10Hz -0.0243527 -0.0308094
+ 6.61e+10Hz -0.0244363 -0.0308166
+ 6.62e+10Hz -0.0245199 -0.0308235
+ 6.63e+10Hz -0.0246037 -0.0308303
+ 6.64e+10Hz -0.0246874 -0.0308369
+ 6.65e+10Hz -0.0247712 -0.0308433
+ 6.66e+10Hz -0.0248551 -0.0308495
+ 6.67e+10Hz -0.024939 -0.0308556
+ 6.68e+10Hz -0.025023 -0.0308614
+ 6.69e+10Hz -0.0251071 -0.0308671
+ 6.7e+10Hz -0.0251912 -0.0308726
+ 6.71e+10Hz -0.0252753 -0.0308779
+ 6.72e+10Hz -0.0253596 -0.030883
+ 6.73e+10Hz -0.0254438 -0.0308879
+ 6.74e+10Hz -0.0255281 -0.0308926
+ 6.75e+10Hz -0.0256125 -0.0308972
+ 6.76e+10Hz -0.025697 -0.0309015
+ 6.77e+10Hz -0.0257815 -0.0309057
+ 6.78e+10Hz -0.025866 -0.0309097
+ 6.79e+10Hz -0.0259506 -0.0309135
+ 6.8e+10Hz -0.0260352 -0.0309171
+ 6.81e+10Hz -0.0261199 -0.0309206
+ 6.82e+10Hz -0.0262046 -0.0309238
+ 6.83e+10Hz -0.0262894 -0.0309268
+ 6.84e+10Hz -0.0263743 -0.0309297
+ 6.85e+10Hz -0.0264592 -0.0309324
+ 6.86e+10Hz -0.0265441 -0.0309348
+ 6.87e+10Hz -0.0266291 -0.0309371
+ 6.88e+10Hz -0.0267141 -0.0309393
+ 6.89e+10Hz -0.0267992 -0.0309412
+ 6.9e+10Hz -0.0268843 -0.0309429
+ 6.91e+10Hz -0.0269695 -0.0309444
+ 6.92e+10Hz -0.0270547 -0.0309458
+ 6.93e+10Hz -0.02714 -0.0309469
+ 6.94e+10Hz -0.0272253 -0.0309479
+ 6.95e+10Hz -0.0273106 -0.0309487
+ 6.96e+10Hz -0.027396 -0.0309493
+ 6.97e+10Hz -0.0274814 -0.0309497
+ 6.98e+10Hz -0.0275669 -0.0309499
+ 6.99e+10Hz -0.0276524 -0.0309499
+ 7e+10Hz -0.027738 -0.0309497
+ 7.01e+10Hz -0.0278236 -0.0309493
+ 7.02e+10Hz -0.0279092 -0.0309488
+ 7.03e+10Hz -0.0279949 -0.0309481
+ 7.04e+10Hz -0.0280806 -0.0309471
+ 7.05e+10Hz -0.0281663 -0.030946
+ 7.06e+10Hz -0.0282521 -0.0309447
+ 7.07e+10Hz -0.028338 -0.0309432
+ 7.08e+10Hz -0.0284238 -0.0309415
+ 7.09e+10Hz -0.0285097 -0.0309396
+ 7.1e+10Hz -0.0285956 -0.0309375
+ 7.11e+10Hz -0.0286816 -0.0309352
+ 7.12e+10Hz -0.0287676 -0.0309328
+ 7.13e+10Hz -0.0288536 -0.0309301
+ 7.14e+10Hz -0.0289397 -0.0309273
+ 7.15e+10Hz -0.0290258 -0.0309243
+ 7.16e+10Hz -0.0291119 -0.030921
+ 7.17e+10Hz -0.0291981 -0.0309176
+ 7.18e+10Hz -0.0292843 -0.030914
+ 7.19e+10Hz -0.0293705 -0.0309102
+ 7.2e+10Hz -0.0294568 -0.0309062
+ 7.21e+10Hz -0.0295431 -0.0309021
+ 7.22e+10Hz -0.0296294 -0.0308977
+ 7.23e+10Hz -0.0297157 -0.0308932
+ 7.24e+10Hz -0.0298021 -0.0308884
+ 7.25e+10Hz -0.0298885 -0.0308835
+ 7.26e+10Hz -0.0299749 -0.0308784
+ 7.27e+10Hz -0.0300614 -0.030873
+ 7.28e+10Hz -0.0301479 -0.0308675
+ 7.29e+10Hz -0.0302344 -0.0308618
+ 7.3e+10Hz -0.0303209 -0.030856
+ 7.31e+10Hz -0.0304075 -0.0308499
+ 7.32e+10Hz -0.0304941 -0.0308436
+ 7.33e+10Hz -0.0305807 -0.0308372
+ 7.34e+10Hz -0.0306673 -0.0308305
+ 7.35e+10Hz -0.030754 -0.0308237
+ 7.36e+10Hz -0.0308407 -0.0308167
+ 7.37e+10Hz -0.0309274 -0.0308095
+ 7.38e+10Hz -0.0310141 -0.0308021
+ 7.39e+10Hz -0.0311009 -0.0307945
+ 7.4e+10Hz -0.0311876 -0.0307867
+ 7.41e+10Hz -0.0312744 -0.0307787
+ 7.42e+10Hz -0.0313613 -0.0307706
+ 7.43e+10Hz -0.0314481 -0.0307622
+ 7.44e+10Hz -0.0315349 -0.0307537
+ 7.45e+10Hz -0.0316218 -0.030745
+ 7.46e+10Hz -0.0317087 -0.0307361
+ 7.47e+10Hz -0.0317956 -0.030727
+ 7.48e+10Hz -0.0318826 -0.0307177
+ 7.49e+10Hz -0.0319695 -0.0307082
+ 7.5e+10Hz -0.0320565 -0.0306985
+ 7.51e+10Hz -0.0321435 -0.0306887
+ 7.52e+10Hz -0.0322305 -0.0306786
+ 7.53e+10Hz -0.0323175 -0.0306684
+ 7.54e+10Hz -0.0324046 -0.030658
+ 7.55e+10Hz -0.0324916 -0.0306474
+ 7.56e+10Hz -0.0325787 -0.0306366
+ 7.57e+10Hz -0.0326658 -0.0306256
+ 7.58e+10Hz -0.0327529 -0.0306145
+ 7.59e+10Hz -0.03284 -0.0306031
+ 7.6e+10Hz -0.0329272 -0.0305916
+ 7.61e+10Hz -0.0330143 -0.0305798
+ 7.62e+10Hz -0.0331015 -0.0305679
+ 7.63e+10Hz -0.0331887 -0.0305558
+ 7.64e+10Hz -0.0332759 -0.0305435
+ 7.65e+10Hz -0.0333631 -0.0305311
+ 7.66e+10Hz -0.0334503 -0.0305184
+ 7.67e+10Hz -0.0335376 -0.0305056
+ 7.68e+10Hz -0.0336248 -0.0304925
+ 7.69e+10Hz -0.0337121 -0.0304793
+ 7.7e+10Hz -0.0337994 -0.0304659
+ 7.71e+10Hz -0.0338867 -0.0304523
+ 7.72e+10Hz -0.033974 -0.0304385
+ 7.73e+10Hz -0.0340613 -0.0304246
+ 7.74e+10Hz -0.0341486 -0.0304104
+ 7.75e+10Hz -0.0342359 -0.0303961
+ 7.76e+10Hz -0.0343233 -0.0303816
+ 7.77e+10Hz -0.0344107 -0.0303668
+ 7.78e+10Hz -0.034498 -0.0303519
+ 7.79e+10Hz -0.0345854 -0.0303369
+ 7.8e+10Hz -0.0346728 -0.0303216
+ 7.81e+10Hz -0.0347602 -0.0303062
+ 7.82e+10Hz -0.0348476 -0.0302905
+ 7.83e+10Hz -0.034935 -0.0302747
+ 7.84e+10Hz -0.0350225 -0.0302587
+ 7.85e+10Hz -0.0351099 -0.0302425
+ 7.86e+10Hz -0.0351974 -0.0302261
+ 7.87e+10Hz -0.0352848 -0.0302095
+ 7.88e+10Hz -0.0353723 -0.0301928
+ 7.89e+10Hz -0.0354598 -0.0301759
+ 7.9e+10Hz -0.0355473 -0.0301587
+ 7.91e+10Hz -0.0356347 -0.0301414
+ 7.92e+10Hz -0.0357222 -0.0301239
+ 7.93e+10Hz -0.0358098 -0.0301063
+ 7.94e+10Hz -0.0358973 -0.0300884
+ 7.95e+10Hz -0.0359848 -0.0300703
+ 7.96e+10Hz -0.0360723 -0.0300521
+ 7.97e+10Hz -0.0361599 -0.0300337
+ 7.98e+10Hz -0.0362474 -0.0300151
+ 7.99e+10Hz -0.036335 -0.0299963
+ 8e+10Hz -0.0364225 -0.0299773
+ 8.01e+10Hz -0.0365101 -0.0299581
+ 8.02e+10Hz -0.0365977 -0.0299388
+ 8.03e+10Hz -0.0366853 -0.0299193
+ 8.04e+10Hz -0.0367728 -0.0298996
+ 8.05e+10Hz -0.0368604 -0.0298797
+ 8.06e+10Hz -0.036948 -0.0298596
+ 8.07e+10Hz -0.0370356 -0.0298393
+ 8.08e+10Hz -0.0371232 -0.0298188
+ 8.09e+10Hz -0.0372108 -0.0297982
+ 8.1e+10Hz -0.0372985 -0.0297773
+ 8.11e+10Hz -0.0373861 -0.0297563
+ 8.12e+10Hz -0.0374737 -0.0297351
+ 8.13e+10Hz -0.0375613 -0.0297137
+ 8.14e+10Hz -0.037649 -0.0296921
+ 8.15e+10Hz -0.0377366 -0.0296704
+ 8.16e+10Hz -0.0378243 -0.0296484
+ 8.17e+10Hz -0.0379119 -0.0296263
+ 8.18e+10Hz -0.0379996 -0.029604
+ 8.19e+10Hz -0.0380872 -0.0295814
+ 8.2e+10Hz -0.0381749 -0.0295587
+ 8.21e+10Hz -0.0382625 -0.0295358
+ 8.22e+10Hz -0.0383502 -0.0295128
+ 8.23e+10Hz -0.0384379 -0.0294895
+ 8.24e+10Hz -0.0385255 -0.0294661
+ 8.25e+10Hz -0.0386132 -0.0294424
+ 8.26e+10Hz -0.0387009 -0.0294186
+ 8.27e+10Hz -0.0387885 -0.0293946
+ 8.28e+10Hz -0.0388762 -0.0293704
+ 8.29e+10Hz -0.0389639 -0.029346
+ 8.3e+10Hz -0.0390516 -0.0293214
+ 8.31e+10Hz -0.0391393 -0.0292967
+ 8.32e+10Hz -0.0392269 -0.0292717
+ 8.33e+10Hz -0.0393146 -0.0292466
+ 8.34e+10Hz -0.0394023 -0.0292212
+ 8.35e+10Hz -0.03949 -0.0291957
+ 8.36e+10Hz -0.0395777 -0.02917
+ 8.37e+10Hz -0.0396654 -0.0291441
+ 8.38e+10Hz -0.039753 -0.029118
+ 8.39e+10Hz -0.0398407 -0.0290917
+ 8.4e+10Hz -0.0399284 -0.0290653
+ 8.41e+10Hz -0.0400161 -0.0290386
+ 8.42e+10Hz -0.0401037 -0.0290118
+ 8.43e+10Hz -0.0401914 -0.0289847
+ 8.44e+10Hz -0.0402791 -0.0289575
+ 8.45e+10Hz -0.0403667 -0.0289301
+ 8.46e+10Hz -0.0404544 -0.0289025
+ 8.47e+10Hz -0.0405421 -0.0288747
+ 8.48e+10Hz -0.0406297 -0.0288467
+ 8.49e+10Hz -0.0407174 -0.0288185
+ 8.5e+10Hz -0.0408051 -0.0287901
+ 8.51e+10Hz -0.0408927 -0.0287615
+ 8.52e+10Hz -0.0409803 -0.0287328
+ 8.53e+10Hz -0.041068 -0.0287038
+ 8.54e+10Hz -0.0411556 -0.0286747
+ 8.55e+10Hz -0.0412432 -0.0286453
+ 8.56e+10Hz -0.0413309 -0.0286158
+ 8.57e+10Hz -0.0414185 -0.0285861
+ 8.58e+10Hz -0.0415061 -0.0285561
+ 8.59e+10Hz -0.0415937 -0.028526
+ 8.6e+10Hz -0.0416813 -0.0284957
+ 8.61e+10Hz -0.0417689 -0.0284652
+ 8.62e+10Hz -0.0418565 -0.0284345
+ 8.63e+10Hz -0.041944 -0.0284036
+ 8.64e+10Hz -0.0420316 -0.0283725
+ 8.65e+10Hz -0.0421192 -0.0283413
+ 8.66e+10Hz -0.0422067 -0.0283098
+ 8.67e+10Hz -0.0422943 -0.0282781
+ 8.68e+10Hz -0.0423818 -0.0282463
+ 8.69e+10Hz -0.0424693 -0.0282142
+ 8.7e+10Hz -0.0425568 -0.0281819
+ 8.71e+10Hz -0.0426443 -0.0281495
+ 8.72e+10Hz -0.0427318 -0.0281168
+ 8.73e+10Hz -0.0428193 -0.028084
+ 8.74e+10Hz -0.0429068 -0.0280509
+ 8.75e+10Hz -0.0429942 -0.0280177
+ 8.76e+10Hz -0.0430816 -0.0279843
+ 8.77e+10Hz -0.0431691 -0.0279506
+ 8.78e+10Hz -0.0432565 -0.0279168
+ 8.79e+10Hz -0.0433439 -0.0278828
+ 8.8e+10Hz -0.0434312 -0.0278485
+ 8.81e+10Hz -0.0435186 -0.0278141
+ 8.82e+10Hz -0.043606 -0.0277795
+ 8.83e+10Hz -0.0436933 -0.0277447
+ 8.84e+10Hz -0.0437806 -0.0277096
+ 8.85e+10Hz -0.0438679 -0.0276744
+ 8.86e+10Hz -0.0439552 -0.027639
+ 8.87e+10Hz -0.0440425 -0.0276034
+ 8.88e+10Hz -0.0441297 -0.0275676
+ 8.89e+10Hz -0.044217 -0.0275316
+ 8.9e+10Hz -0.0443042 -0.0274954
+ 8.91e+10Hz -0.0443914 -0.0274589
+ 8.92e+10Hz -0.0444785 -0.0274223
+ 8.93e+10Hz -0.0445657 -0.0273855
+ 8.94e+10Hz -0.0446528 -0.0273485
+ 8.95e+10Hz -0.0447399 -0.0273113
+ 8.96e+10Hz -0.044827 -0.0272739
+ 8.97e+10Hz -0.0449141 -0.0272363
+ 8.98e+10Hz -0.0450011 -0.0271984
+ 8.99e+10Hz -0.0450881 -0.0271604
+ 9e+10Hz -0.0451751 -0.0271222
+ 9.01e+10Hz -0.0452621 -0.0270838
+ 9.02e+10Hz -0.045349 -0.0270452
+ 9.03e+10Hz -0.0454359 -0.0270064
+ 9.04e+10Hz -0.0455228 -0.0269674
+ 9.05e+10Hz -0.0456097 -0.0269281
+ 9.06e+10Hz -0.0456965 -0.0268887
+ 9.07e+10Hz -0.0457833 -0.0268491
+ 9.08e+10Hz -0.0458701 -0.0268093
+ 9.09e+10Hz -0.0459569 -0.0267693
+ 9.1e+10Hz -0.0460436 -0.026729
+ 9.11e+10Hz -0.0461303 -0.0266886
+ 9.12e+10Hz -0.0462169 -0.026648
+ 9.13e+10Hz -0.0463036 -0.0266071
+ 9.14e+10Hz -0.0463902 -0.0265661
+ 9.15e+10Hz -0.0464767 -0.0265249
+ 9.16e+10Hz -0.0465633 -0.0264834
+ 9.17e+10Hz -0.0466497 -0.0264418
+ 9.18e+10Hz -0.0467362 -0.0263999
+ 9.19e+10Hz -0.0468227 -0.0263579
+ 9.2e+10Hz -0.0469091 -0.0263157
+ 9.21e+10Hz -0.0469954 -0.0262732
+ 9.22e+10Hz -0.0470817 -0.0262306
+ 9.23e+10Hz -0.047168 -0.0261877
+ 9.24e+10Hz -0.0472543 -0.0261447
+ 9.25e+10Hz -0.0473405 -0.0261014
+ 9.26e+10Hz -0.0474267 -0.026058
+ 9.27e+10Hz -0.0475128 -0.0260143
+ 9.28e+10Hz -0.0475989 -0.0259705
+ 9.29e+10Hz -0.0476849 -0.0259264
+ 9.3e+10Hz -0.047771 -0.0258821
+ 9.31e+10Hz -0.0478569 -0.0258377
+ 9.32e+10Hz -0.0479429 -0.025793
+ 9.33e+10Hz -0.0480288 -0.0257482
+ 9.34e+10Hz -0.0481146 -0.0257031
+ 9.35e+10Hz -0.0482004 -0.0256578
+ 9.36e+10Hz -0.0482862 -0.0256123
+ 9.37e+10Hz -0.0483719 -0.0255667
+ 9.38e+10Hz -0.0484576 -0.0255208
+ 9.39e+10Hz -0.0485432 -0.0254748
+ 9.4e+10Hz -0.0486288 -0.0254285
+ 9.41e+10Hz -0.0487143 -0.025382
+ 9.42e+10Hz -0.0487998 -0.0253353
+ 9.43e+10Hz -0.0488852 -0.0252885
+ 9.44e+10Hz -0.0489706 -0.0252414
+ 9.45e+10Hz -0.049056 -0.0251941
+ 9.46e+10Hz -0.0491413 -0.0251466
+ 9.47e+10Hz -0.0492265 -0.025099
+ 9.48e+10Hz -0.0493117 -0.0250511
+ 9.49e+10Hz -0.0493969 -0.025003
+ 9.5e+10Hz -0.049482 -0.0249548
+ 9.51e+10Hz -0.049567 -0.0249063
+ 9.52e+10Hz -0.049652 -0.0248576
+ 9.53e+10Hz -0.0497369 -0.0248087
+ 9.54e+10Hz -0.0498218 -0.0247597
+ 9.55e+10Hz -0.0499066 -0.0247104
+ 9.56e+10Hz -0.0499914 -0.024661
+ 9.57e+10Hz -0.0500761 -0.0246113
+ 9.58e+10Hz -0.0501608 -0.0245614
+ 9.59e+10Hz -0.0502454 -0.0245114
+ 9.6e+10Hz -0.05033 -0.0244611
+ 9.61e+10Hz -0.0504145 -0.0244107
+ 9.62e+10Hz -0.0504989 -0.02436
+ 9.63e+10Hz -0.0505833 -0.0243092
+ 9.64e+10Hz -0.0506676 -0.0242581
+ 9.65e+10Hz -0.0507519 -0.0242069
+ 9.66e+10Hz -0.0508361 -0.0241554
+ 9.67e+10Hz -0.0509202 -0.0241038
+ 9.68e+10Hz -0.0510043 -0.024052
+ 9.69e+10Hz -0.0510883 -0.024
+ 9.7e+10Hz -0.0511723 -0.0239477
+ 9.71e+10Hz -0.0512562 -0.0238953
+ 9.72e+10Hz -0.05134 -0.0238427
+ 9.73e+10Hz -0.0514238 -0.0237899
+ 9.74e+10Hz -0.0515075 -0.0237369
+ 9.75e+10Hz -0.0515912 -0.0236837
+ 9.76e+10Hz -0.0516748 -0.0236303
+ 9.77e+10Hz -0.0517583 -0.0235768
+ 9.78e+10Hz -0.0518418 -0.023523
+ 9.79e+10Hz -0.0519252 -0.023469
+ 9.8e+10Hz -0.0520085 -0.0234149
+ 9.81e+10Hz -0.0520918 -0.0233605
+ 9.82e+10Hz -0.052175 -0.023306
+ 9.83e+10Hz -0.0522582 -0.0232512
+ 9.84e+10Hz -0.0523412 -0.0231963
+ 9.85e+10Hz -0.0524242 -0.0231412
+ 9.86e+10Hz -0.0525072 -0.0230859
+ 9.87e+10Hz -0.05259 -0.0230304
+ 9.88e+10Hz -0.0526729 -0.0229747
+ 9.89e+10Hz -0.0527556 -0.0229188
+ 9.9e+10Hz -0.0528383 -0.0228627
+ 9.91e+10Hz -0.0529209 -0.0228064
+ 9.92e+10Hz -0.0530034 -0.02275
+ 9.93e+10Hz -0.0530859 -0.0226933
+ 9.94e+10Hz -0.0531683 -0.0226365
+ 9.95e+10Hz -0.0532506 -0.0225795
+ 9.96e+10Hz -0.0533328 -0.0225223
+ 9.97e+10Hz -0.053415 -0.0224649
+ 9.98e+10Hz -0.0534971 -0.0224073
+ 9.99e+10Hz -0.0535792 -0.0223495
+ 1e+11Hz -0.0536611 -0.0222915
+ 1.001e+11Hz -0.053743 -0.0222334
+ 1.002e+11Hz -0.0538249 -0.022175
+ 1.003e+11Hz -0.0539066 -0.0221165
+ 1.004e+11Hz -0.0539883 -0.0220578
+ 1.005e+11Hz -0.0540699 -0.0219989
+ 1.006e+11Hz -0.0541514 -0.0219398
+ 1.007e+11Hz -0.0542329 -0.0218805
+ 1.008e+11Hz -0.0543143 -0.021821
+ 1.009e+11Hz -0.0543956 -0.0217614
+ 1.01e+11Hz -0.0544768 -0.0217016
+ 1.011e+11Hz -0.054558 -0.0216415
+ 1.012e+11Hz -0.0546391 -0.0215813
+ 1.013e+11Hz -0.0547201 -0.021521
+ 1.014e+11Hz -0.0548011 -0.0214604
+ 1.015e+11Hz -0.0548819 -0.0213996
+ 1.016e+11Hz -0.0549627 -0.0213387
+ 1.017e+11Hz -0.0550435 -0.0212775
+ 1.018e+11Hz -0.0551241 -0.0212162
+ 1.019e+11Hz -0.0552047 -0.0211547
+ 1.02e+11Hz -0.0552851 -0.0210931
+ 1.021e+11Hz -0.0553656 -0.0210312
+ 1.022e+11Hz -0.0554459 -0.0209692
+ 1.023e+11Hz -0.0555262 -0.0209069
+ 1.024e+11Hz -0.0556064 -0.0208445
+ 1.025e+11Hz -0.0556865 -0.0207819
+ 1.026e+11Hz -0.0557665 -0.0207191
+ 1.027e+11Hz -0.0558464 -0.0206562
+ 1.028e+11Hz -0.0559263 -0.0205931
+ 1.029e+11Hz -0.0560061 -0.0205297
+ 1.03e+11Hz -0.0560858 -0.0204662
+ 1.031e+11Hz -0.0561655 -0.0204025
+ 1.032e+11Hz -0.0562451 -0.0203387
+ 1.033e+11Hz -0.0563246 -0.0202746
+ 1.034e+11Hz -0.056404 -0.0202104
+ 1.035e+11Hz -0.0564833 -0.020146
+ 1.036e+11Hz -0.0565626 -0.0200814
+ 1.037e+11Hz -0.0566417 -0.0200166
+ 1.038e+11Hz -0.0567208 -0.0199516
+ 1.039e+11Hz -0.0567998 -0.0198865
+ 1.04e+11Hz -0.0568788 -0.0198212
+ 1.041e+11Hz -0.0569576 -0.0197557
+ 1.042e+11Hz -0.0570364 -0.01969
+ 1.043e+11Hz -0.0571151 -0.0196241
+ 1.044e+11Hz -0.0571937 -0.0195581
+ 1.045e+11Hz -0.0572723 -0.0194919
+ 1.046e+11Hz -0.0573507 -0.0194255
+ 1.047e+11Hz -0.0574291 -0.0193589
+ 1.048e+11Hz -0.0575074 -0.0192921
+ 1.049e+11Hz -0.0575856 -0.0192252
+ 1.05e+11Hz -0.0576637 -0.0191581
+ 1.051e+11Hz -0.0577418 -0.0190908
+ 1.052e+11Hz -0.0578198 -0.0190233
+ 1.053e+11Hz -0.0578977 -0.0189556
+ 1.054e+11Hz -0.0579755 -0.0188878
+ 1.055e+11Hz -0.0580532 -0.0188197
+ 1.056e+11Hz -0.0581308 -0.0187515
+ 1.057e+11Hz -0.0582084 -0.0186832
+ 1.058e+11Hz -0.0582859 -0.0186146
+ 1.059e+11Hz -0.0583633 -0.0185459
+ 1.06e+11Hz -0.0584406 -0.0184769
+ 1.061e+11Hz -0.0585178 -0.0184078
+ 1.062e+11Hz -0.058595 -0.0183385
+ 1.063e+11Hz -0.0586721 -0.0182691
+ 1.064e+11Hz -0.058749 -0.0181994
+ 1.065e+11Hz -0.0588259 -0.0181296
+ 1.066e+11Hz -0.0589028 -0.0180596
+ 1.067e+11Hz -0.0589795 -0.0179894
+ 1.068e+11Hz -0.0590561 -0.017919
+ 1.069e+11Hz -0.0591327 -0.0178485
+ 1.07e+11Hz -0.0592092 -0.0177778
+ 1.071e+11Hz -0.0592856 -0.0177069
+ 1.072e+11Hz -0.0593619 -0.0176358
+ 1.073e+11Hz -0.0594381 -0.0175645
+ 1.074e+11Hz -0.0595143 -0.017493
+ 1.075e+11Hz -0.0595903 -0.0174214
+ 1.076e+11Hz -0.0596663 -0.0173496
+ 1.077e+11Hz -0.0597422 -0.0172776
+ 1.078e+11Hz -0.059818 -0.0172054
+ 1.079e+11Hz -0.0598937 -0.0171331
+ 1.08e+11Hz -0.0599693 -0.0170606
+ 1.081e+11Hz -0.0600448 -0.0169878
+ 1.082e+11Hz -0.0601203 -0.0169149
+ 1.083e+11Hz -0.0601957 -0.0168418
+ 1.084e+11Hz -0.0602709 -0.0167686
+ 1.085e+11Hz -0.0603461 -0.0166951
+ 1.086e+11Hz -0.0604212 -0.0166215
+ 1.087e+11Hz -0.0604962 -0.0165477
+ 1.088e+11Hz -0.0605711 -0.0164737
+ 1.089e+11Hz -0.060646 -0.0163995
+ 1.09e+11Hz -0.0607207 -0.0163252
+ 1.091e+11Hz -0.0607953 -0.0162506
+ 1.092e+11Hz -0.0608699 -0.0161759
+ 1.093e+11Hz -0.0609444 -0.016101
+ 1.094e+11Hz -0.0610187 -0.0160259
+ 1.095e+11Hz -0.061093 -0.0159507
+ 1.096e+11Hz -0.0611672 -0.0158752
+ 1.097e+11Hz -0.0612413 -0.0157996
+ 1.098e+11Hz -0.0613153 -0.0157238
+ 1.099e+11Hz -0.0613892 -0.0156477
+ 1.1e+11Hz -0.0614631 -0.0155716
+ 1.101e+11Hz -0.0615368 -0.0154952
+ 1.102e+11Hz -0.0616104 -0.0154186
+ 1.103e+11Hz -0.061684 -0.0153419
+ 1.104e+11Hz -0.0617574 -0.015265
+ 1.105e+11Hz -0.0618308 -0.0151879
+ 1.106e+11Hz -0.061904 -0.0151106
+ 1.107e+11Hz -0.0619772 -0.0150331
+ 1.108e+11Hz -0.0620503 -0.0149554
+ 1.109e+11Hz -0.0621232 -0.0148776
+ 1.11e+11Hz -0.0621961 -0.0147996
+ 1.111e+11Hz -0.0622689 -0.0147213
+ 1.112e+11Hz -0.0623415 -0.014643
+ 1.113e+11Hz -0.0624141 -0.0145644
+ 1.114e+11Hz -0.0624866 -0.0144856
+ 1.115e+11Hz -0.0625589 -0.0144066
+ 1.116e+11Hz -0.0626312 -0.0143275
+ 1.117e+11Hz -0.0627034 -0.0142482
+ 1.118e+11Hz -0.0627754 -0.0141687
+ 1.119e+11Hz -0.0628474 -0.014089
+ 1.12e+11Hz -0.0629193 -0.0140091
+ 1.121e+11Hz -0.0629911 -0.013929
+ 1.122e+11Hz -0.0630627 -0.0138488
+ 1.123e+11Hz -0.0631343 -0.0137683
+ 1.124e+11Hz -0.0632057 -0.0136877
+ 1.125e+11Hz -0.0632771 -0.0136069
+ 1.126e+11Hz -0.0633483 -0.0135259
+ 1.127e+11Hz -0.0634194 -0.0134447
+ 1.128e+11Hz -0.0634905 -0.0133633
+ 1.129e+11Hz -0.0635614 -0.0132818
+ 1.13e+11Hz -0.0636322 -0.0132
+ 1.131e+11Hz -0.0637029 -0.0131181
+ 1.132e+11Hz -0.0637735 -0.013036
+ 1.133e+11Hz -0.063844 -0.0129537
+ 1.134e+11Hz -0.0639144 -0.0128712
+ 1.135e+11Hz -0.0639846 -0.0127885
+ 1.136e+11Hz -0.0640548 -0.0127056
+ 1.137e+11Hz -0.0641248 -0.0126226
+ 1.138e+11Hz -0.0641948 -0.0125394
+ 1.139e+11Hz -0.0642646 -0.0124559
+ 1.14e+11Hz -0.0643343 -0.0123723
+ 1.141e+11Hz -0.0644039 -0.0122885
+ 1.142e+11Hz -0.0644734 -0.0122046
+ 1.143e+11Hz -0.0645427 -0.0121204
+ 1.144e+11Hz -0.064612 -0.012036
+ 1.145e+11Hz -0.0646811 -0.0119515
+ 1.146e+11Hz -0.0647501 -0.0118668
+ 1.147e+11Hz -0.064819 -0.0117819
+ 1.148e+11Hz -0.0648878 -0.0116968
+ 1.149e+11Hz -0.0649564 -0.0116115
+ 1.15e+11Hz -0.0650249 -0.011526
+ 1.151e+11Hz -0.0650934 -0.0114404
+ 1.152e+11Hz -0.0651617 -0.0113545
+ 1.153e+11Hz -0.0652298 -0.0112685
+ 1.154e+11Hz -0.0652979 -0.0111823
+ 1.155e+11Hz -0.0653658 -0.0110959
+ 1.156e+11Hz -0.0654336 -0.0110093
+ 1.157e+11Hz -0.0655013 -0.0109225
+ 1.158e+11Hz -0.0655688 -0.0108356
+ 1.159e+11Hz -0.0656362 -0.0107485
+ 1.16e+11Hz -0.0657035 -0.0106611
+ 1.161e+11Hz -0.0657707 -0.0105737
+ 1.162e+11Hz -0.0658378 -0.010486
+ 1.163e+11Hz -0.0659047 -0.0103981
+ 1.164e+11Hz -0.0659715 -0.01031
+ 1.165e+11Hz -0.0660381 -0.0102218
+ 1.166e+11Hz -0.0661046 -0.0101334
+ 1.167e+11Hz -0.066171 -0.0100448
+ 1.168e+11Hz -0.0662373 -0.00995601
+ 1.169e+11Hz -0.0663034 -0.00986704
+ 1.17e+11Hz -0.0663694 -0.0097779
+ 1.171e+11Hz -0.0664353 -0.00968857
+ 1.172e+11Hz -0.066501 -0.00959906
+ 1.173e+11Hz -0.0665666 -0.00950937
+ 1.174e+11Hz -0.066632 -0.00941949
+ 1.175e+11Hz -0.0666974 -0.00932944
+ 1.176e+11Hz -0.0667626 -0.00923921
+ 1.177e+11Hz -0.0668276 -0.0091488
+ 1.178e+11Hz -0.0668925 -0.0090582
+ 1.179e+11Hz -0.0669573 -0.00896743
+ 1.18e+11Hz -0.0670219 -0.00887648
+ 1.181e+11Hz -0.0670864 -0.00878536
+ 1.182e+11Hz -0.0671508 -0.00869405
+ 1.183e+11Hz -0.067215 -0.00860257
+ 1.184e+11Hz -0.067279 -0.00851091
+ 1.185e+11Hz -0.067343 -0.00841907
+ 1.186e+11Hz -0.0674067 -0.00832705
+ 1.187e+11Hz -0.0674704 -0.00823486
+ 1.188e+11Hz -0.0675339 -0.0081425
+ 1.189e+11Hz -0.0675972 -0.00804995
+ 1.19e+11Hz -0.0676604 -0.00795724
+ 1.191e+11Hz -0.0677235 -0.00786435
+ 1.192e+11Hz -0.0677864 -0.00777128
+ 1.193e+11Hz -0.0678492 -0.00767804
+ 1.194e+11Hz -0.0679118 -0.00758463
+ 1.195e+11Hz -0.0679743 -0.00749105
+ 1.196e+11Hz -0.0680366 -0.00739729
+ 1.197e+11Hz -0.0680988 -0.00730337
+ 1.198e+11Hz -0.0681608 -0.00720927
+ 1.199e+11Hz -0.0682227 -0.007115
+ 1.2e+11Hz -0.0682844 -0.00702056
+ 1.201e+11Hz -0.068346 -0.00692595
+ 1.202e+11Hz -0.0684074 -0.00683117
+ 1.203e+11Hz -0.0684687 -0.00673622
+ 1.204e+11Hz -0.0685298 -0.0066411
+ 1.205e+11Hz -0.0685907 -0.00654582
+ 1.206e+11Hz -0.0686516 -0.00645037
+ 1.207e+11Hz -0.0687122 -0.00635475
+ 1.208e+11Hz -0.0687727 -0.00625896
+ 1.209e+11Hz -0.0688331 -0.00616301
+ 1.21e+11Hz -0.0688933 -0.0060669
+ 1.211e+11Hz -0.0689533 -0.00597062
+ 1.212e+11Hz -0.0690132 -0.00587417
+ 1.213e+11Hz -0.0690729 -0.00577756
+ 1.214e+11Hz -0.0691325 -0.00568079
+ 1.215e+11Hz -0.0691919 -0.00558386
+ 1.216e+11Hz -0.0692512 -0.00548676
+ 1.217e+11Hz -0.0693103 -0.00538951
+ 1.218e+11Hz -0.0693692 -0.00529209
+ 1.219e+11Hz -0.069428 -0.00519451
+ 1.22e+11Hz -0.0694866 -0.00509677
+ 1.221e+11Hz -0.0695451 -0.00499887
+ 1.222e+11Hz -0.0696034 -0.00490082
+ 1.223e+11Hz -0.0696616 -0.0048026
+ 1.224e+11Hz -0.0697196 -0.00470423
+ 1.225e+11Hz -0.0697774 -0.0046057
+ 1.226e+11Hz -0.0698351 -0.00450701
+ 1.227e+11Hz -0.0698926 -0.00440817
+ 1.228e+11Hz -0.0699499 -0.00430917
+ 1.229e+11Hz -0.0700071 -0.00421002
+ 1.23e+11Hz -0.0700642 -0.00411071
+ 1.231e+11Hz -0.070121 -0.00401125
+ 1.232e+11Hz -0.0701777 -0.00391163
+ 1.233e+11Hz -0.0702343 -0.00381186
+ 1.234e+11Hz -0.0702907 -0.00371194
+ 1.235e+11Hz -0.0703469 -0.00361187
+ 1.236e+11Hz -0.070403 -0.00351164
+ 1.237e+11Hz -0.0704589 -0.00341127
+ 1.238e+11Hz -0.0705146 -0.00331074
+ 1.239e+11Hz -0.0705702 -0.00321007
+ 1.24e+11Hz -0.0706256 -0.00310924
+ 1.241e+11Hz -0.0706809 -0.00300827
+ 1.242e+11Hz -0.070736 -0.00290714
+ 1.243e+11Hz -0.0707909 -0.00280588
+ 1.244e+11Hz -0.0708456 -0.00270446
+ 1.245e+11Hz -0.0709002 -0.00260289
+ 1.246e+11Hz -0.0709547 -0.00250118
+ 1.247e+11Hz -0.071009 -0.00239932
+ 1.248e+11Hz -0.0710631 -0.00229732
+ 1.249e+11Hz -0.071117 -0.00219517
+ 1.25e+11Hz -0.0711708 -0.00209288
+ 1.251e+11Hz -0.0712244 -0.00199044
+ 1.252e+11Hz -0.0712779 -0.00188786
+ 1.253e+11Hz -0.0713312 -0.00178513
+ 1.254e+11Hz -0.0713843 -0.00168226
+ 1.255e+11Hz -0.0714373 -0.00157925
+ 1.256e+11Hz -0.0714901 -0.0014761
+ 1.257e+11Hz -0.0715428 -0.0013728
+ 1.258e+11Hz -0.0715953 -0.00126936
+ 1.259e+11Hz -0.0716476 -0.00116578
+ 1.26e+11Hz -0.0716997 -0.00106207
+ 1.261e+11Hz -0.0717517 -0.000958205
+ 1.262e+11Hz -0.0718036 -0.000854205
+ 1.263e+11Hz -0.0718552 -0.000750064
+ 1.264e+11Hz -0.0719068 -0.000645784
+ 1.265e+11Hz -0.0719581 -0.000541365
+ 1.266e+11Hz -0.0720093 -0.000436806
+ 1.267e+11Hz -0.0720603 -0.000332109
+ 1.268e+11Hz -0.0721112 -0.000227273
+ 1.269e+11Hz -0.0721619 -0.000122299
+ 1.27e+11Hz -0.0722124 -1.71872e-05
+ 1.271e+11Hz -0.0722628 8.80626e-05
+ 1.272e+11Hz -0.072313 0.00019345
+ 1.273e+11Hz -0.072363 0.000298974
+ 1.274e+11Hz -0.0724129 0.000404636
+ 1.275e+11Hz -0.0724627 0.000510435
+ 1.276e+11Hz -0.0725122 0.00061637
+ 1.277e+11Hz -0.0725616 0.000722442
+ 1.278e+11Hz -0.0726109 0.000828651
+ 1.279e+11Hz -0.0726599 0.000934995
+ 1.28e+11Hz -0.0727089 0.00104148
+ 1.281e+11Hz -0.0727576 0.00114809
+ 1.282e+11Hz -0.0728062 0.00125485
+ 1.283e+11Hz -0.0728547 0.00136173
+ 1.284e+11Hz -0.0729029 0.00146876
+ 1.285e+11Hz -0.0729511 0.00157592
+ 1.286e+11Hz -0.072999 0.00168321
+ 1.287e+11Hz -0.0730468 0.00179064
+ 1.288e+11Hz -0.0730944 0.00189821
+ 1.289e+11Hz -0.0731419 0.00200591
+ 1.29e+11Hz -0.0731892 0.00211375
+ 1.291e+11Hz -0.0732364 0.00222172
+ 1.292e+11Hz -0.0732834 0.00232983
+ 1.293e+11Hz -0.0733302 0.00243807
+ 1.294e+11Hz -0.0733769 0.00254645
+ 1.295e+11Hz -0.0734234 0.00265497
+ 1.296e+11Hz -0.0734697 0.00276362
+ 1.297e+11Hz -0.0735159 0.0028724
+ 1.298e+11Hz -0.073562 0.00298132
+ 1.299e+11Hz -0.0736079 0.00309038
+ 1.3e+11Hz -0.0736536 0.00319958
+ 1.301e+11Hz -0.0736991 0.0033089
+ 1.302e+11Hz -0.0737445 0.00341837
+ 1.303e+11Hz -0.0737898 0.00352797
+ 1.304e+11Hz -0.0738348 0.00363771
+ 1.305e+11Hz -0.0738797 0.00374758
+ 1.306e+11Hz -0.0739245 0.00385759
+ 1.307e+11Hz -0.0739691 0.00396774
+ 1.308e+11Hz -0.0740135 0.00407802
+ 1.309e+11Hz -0.0740578 0.00418844
+ 1.31e+11Hz -0.0741019 0.004299
+ 1.311e+11Hz -0.0741459 0.0044097
+ 1.312e+11Hz -0.0741897 0.00452053
+ 1.313e+11Hz -0.0742334 0.00463151
+ 1.314e+11Hz -0.0742768 0.00474262
+ 1.315e+11Hz -0.0743202 0.00485386
+ 1.316e+11Hz -0.0743633 0.00496525
+ 1.317e+11Hz -0.0744063 0.00507678
+ 1.318e+11Hz -0.0744492 0.00518844
+ 1.319e+11Hz -0.0744918 0.00530025
+ 1.32e+11Hz -0.0745343 0.00541219
+ 1.321e+11Hz -0.0745767 0.00552428
+ 1.322e+11Hz -0.0746189 0.0056365
+ 1.323e+11Hz -0.0746609 0.00574886
+ 1.324e+11Hz -0.0747028 0.00586137
+ 1.325e+11Hz -0.0747445 0.00597402
+ 1.326e+11Hz -0.0747861 0.0060868
+ 1.327e+11Hz -0.0748275 0.00619973
+ 1.328e+11Hz -0.0748687 0.00631281
+ 1.329e+11Hz -0.0749098 0.00642602
+ 1.33e+11Hz -0.0749507 0.00653937
+ 1.331e+11Hz -0.0749914 0.00665287
+ 1.332e+11Hz -0.075032 0.00676651
+ 1.333e+11Hz -0.0750724 0.0068803
+ 1.334e+11Hz -0.0751126 0.00699423
+ 1.335e+11Hz -0.0751527 0.0071083
+ 1.336e+11Hz -0.0751926 0.00722252
+ 1.337e+11Hz -0.0752324 0.00733688
+ 1.338e+11Hz -0.075272 0.00745139
+ 1.339e+11Hz -0.0753114 0.00756604
+ 1.34e+11Hz -0.0753506 0.00768084
+ 1.341e+11Hz -0.0753897 0.00779579
+ 1.342e+11Hz -0.0754286 0.00791088
+ 1.343e+11Hz -0.0754674 0.00802612
+ 1.344e+11Hz -0.075506 0.0081415
+ 1.345e+11Hz -0.0755444 0.00825703
+ 1.346e+11Hz -0.0755826 0.00837271
+ 1.347e+11Hz -0.0756207 0.00848854
+ 1.348e+11Hz -0.0756586 0.00860451
+ 1.349e+11Hz -0.0756963 0.00872063
+ 1.35e+11Hz -0.0757339 0.00883691
+ 1.351e+11Hz -0.0757713 0.00895333
+ 1.352e+11Hz -0.0758085 0.0090699
+ 1.353e+11Hz -0.0758455 0.00918662
+ 1.354e+11Hz -0.0758824 0.00930348
+ 1.355e+11Hz -0.0759191 0.0094205
+ 1.356e+11Hz -0.0759556 0.00953767
+ 1.357e+11Hz -0.0759919 0.00965499
+ 1.358e+11Hz -0.0760281 0.00977246
+ 1.359e+11Hz -0.0760641 0.00989008
+ 1.36e+11Hz -0.0760999 0.0100079
+ 1.361e+11Hz -0.0761355 0.0101258
+ 1.362e+11Hz -0.076171 0.0102439
+ 1.363e+11Hz -0.0762062 0.0103621
+ 1.364e+11Hz -0.0762413 0.0104805
+ 1.365e+11Hz -0.0762762 0.010599
+ 1.366e+11Hz -0.0763109 0.0107177
+ 1.367e+11Hz -0.0763455 0.0108365
+ 1.368e+11Hz -0.0763798 0.0109555
+ 1.369e+11Hz -0.076414 0.0110746
+ 1.37e+11Hz -0.076448 0.0111939
+ 1.371e+11Hz -0.0764818 0.0113133
+ 1.372e+11Hz -0.0765154 0.011433
+ 1.373e+11Hz -0.0765488 0.0115527
+ 1.374e+11Hz -0.076582 0.0116726
+ 1.375e+11Hz -0.0766151 0.0117927
+ 1.376e+11Hz -0.0766479 0.0119128
+ 1.377e+11Hz -0.0766806 0.0120332
+ 1.378e+11Hz -0.076713 0.0121537
+ 1.379e+11Hz -0.0767453 0.0122744
+ 1.38e+11Hz -0.0767773 0.0123952
+ 1.381e+11Hz -0.0768092 0.0125162
+ 1.382e+11Hz -0.0768409 0.0126373
+ 1.383e+11Hz -0.0768724 0.0127586
+ 1.384e+11Hz -0.0769037 0.01288
+ 1.385e+11Hz -0.0769347 0.0130016
+ 1.386e+11Hz -0.0769656 0.0131233
+ 1.387e+11Hz -0.0769963 0.0132452
+ 1.388e+11Hz -0.0770268 0.0133672
+ 1.389e+11Hz -0.0770571 0.0134894
+ 1.39e+11Hz -0.0770871 0.0136117
+ 1.391e+11Hz -0.077117 0.0137342
+ 1.392e+11Hz -0.0771466 0.0138568
+ 1.393e+11Hz -0.0771761 0.0139796
+ 1.394e+11Hz -0.0772053 0.0141025
+ 1.395e+11Hz -0.0772344 0.0142256
+ 1.396e+11Hz -0.0772632 0.0143488
+ 1.397e+11Hz -0.0772918 0.0144722
+ 1.398e+11Hz -0.0773202 0.0145957
+ 1.399e+11Hz -0.0773484 0.0147194
+ 1.4e+11Hz -0.0773763 0.0148432
+ 1.401e+11Hz -0.0774041 0.0149672
+ 1.402e+11Hz -0.0774316 0.0150913
+ 1.403e+11Hz -0.0774589 0.0152155
+ 1.404e+11Hz -0.077486 0.0153399
+ 1.405e+11Hz -0.0775129 0.0154645
+ 1.406e+11Hz -0.0775396 0.0155891
+ 1.407e+11Hz -0.077566 0.015714
+ 1.408e+11Hz -0.0775922 0.015839
+ 1.409e+11Hz -0.0776182 0.0159641
+ 1.41e+11Hz -0.077644 0.0160893
+ 1.411e+11Hz -0.0776695 0.0162147
+ 1.412e+11Hz -0.0776949 0.0163403
+ 1.413e+11Hz -0.0777199 0.0164659
+ 1.414e+11Hz -0.0777448 0.0165917
+ 1.415e+11Hz -0.0777695 0.0167177
+ 1.416e+11Hz -0.0777939 0.0168438
+ 1.417e+11Hz -0.077818 0.01697
+ 1.418e+11Hz -0.077842 0.0170963
+ 1.419e+11Hz -0.0778657 0.0172228
+ 1.42e+11Hz -0.0778892 0.0173495
+ 1.421e+11Hz -0.0779124 0.0174762
+ 1.422e+11Hz -0.0779354 0.0176031
+ 1.423e+11Hz -0.0779582 0.0177301
+ 1.424e+11Hz -0.0779808 0.0178573
+ 1.425e+11Hz -0.0780031 0.0179845
+ 1.426e+11Hz -0.0780251 0.018112
+ 1.427e+11Hz -0.078047 0.0182395
+ 1.428e+11Hz -0.0780686 0.0183671
+ 1.429e+11Hz -0.0780899 0.0184949
+ 1.43e+11Hz -0.078111 0.0186228
+ 1.431e+11Hz -0.0781319 0.0187509
+ 1.432e+11Hz -0.0781525 0.018879
+ 1.433e+11Hz -0.0781729 0.0190073
+ 1.434e+11Hz -0.0781931 0.0191357
+ 1.435e+11Hz -0.078213 0.0192642
+ 1.436e+11Hz -0.0782326 0.0193928
+ 1.437e+11Hz -0.0782521 0.0195215
+ 1.438e+11Hz -0.0782712 0.0196504
+ 1.439e+11Hz -0.0782902 0.0197794
+ 1.44e+11Hz -0.0783089 0.0199084
+ 1.441e+11Hz -0.0783273 0.0200376
+ 1.442e+11Hz -0.0783455 0.0201669
+ 1.443e+11Hz -0.0783634 0.0202963
+ 1.444e+11Hz -0.0783811 0.0204259
+ 1.445e+11Hz -0.0783986 0.0205555
+ 1.446e+11Hz -0.0784158 0.0206852
+ 1.447e+11Hz -0.0784328 0.0208151
+ 1.448e+11Hz -0.0784495 0.020945
+ 1.449e+11Hz -0.078466 0.021075
+ 1.45e+11Hz -0.0784822 0.0212052
+ 1.451e+11Hz -0.0784981 0.0213354
+ 1.452e+11Hz -0.0785139 0.0214657
+ 1.453e+11Hz -0.0785293 0.0215962
+ 1.454e+11Hz -0.0785446 0.0217267
+ 1.455e+11Hz -0.0785595 0.0218573
+ 1.456e+11Hz -0.0785743 0.021988
+ 1.457e+11Hz -0.0785887 0.0221188
+ 1.458e+11Hz -0.078603 0.0222497
+ 1.459e+11Hz -0.078617 0.0223807
+ 1.46e+11Hz -0.0786307 0.0225118
+ 1.461e+11Hz -0.0786442 0.022643
+ 1.462e+11Hz -0.0786574 0.0227742
+ 1.463e+11Hz -0.0786704 0.0229055
+ 1.464e+11Hz -0.0786832 0.0230369
+ 1.465e+11Hz -0.0786957 0.0231684
+ 1.466e+11Hz -0.0787079 0.0233
+ 1.467e+11Hz -0.0787199 0.0234317
+ 1.468e+11Hz -0.0787317 0.0235634
+ 1.469e+11Hz -0.0787432 0.0236952
+ 1.47e+11Hz -0.0787545 0.0238271
+ 1.471e+11Hz -0.0787655 0.023959
+ 1.472e+11Hz -0.0787763 0.0240911
+ 1.473e+11Hz -0.0787869 0.0242232
+ 1.474e+11Hz -0.0787971 0.0243554
+ 1.475e+11Hz -0.0788072 0.0244876
+ 1.476e+11Hz -0.078817 0.0246199
+ 1.477e+11Hz -0.0788266 0.0247523
+ 1.478e+11Hz -0.0788359 0.0248848
+ 1.479e+11Hz -0.078845 0.0250173
+ 1.48e+11Hz -0.0788539 0.0251499
+ 1.481e+11Hz -0.0788625 0.0252825
+ 1.482e+11Hz -0.0788708 0.0254152
+ 1.483e+11Hz -0.078879 0.025548
+ 1.484e+11Hz -0.0788869 0.0256808
+ 1.485e+11Hz -0.0788945 0.0258137
+ 1.486e+11Hz -0.078902 0.0259467
+ 1.487e+11Hz -0.0789092 0.0260796
+ 1.488e+11Hz -0.0789161 0.0262127
+ 1.489e+11Hz -0.0789228 0.0263458
+ 1.49e+11Hz -0.0789293 0.026479
+ 1.491e+11Hz -0.0789356 0.0266123
+ 1.492e+11Hz -0.0789416 0.0267455
+ 1.493e+11Hz -0.0789475 0.0268789
+ 1.494e+11Hz -0.078953 0.0270123
+ 1.495e+11Hz -0.0789584 0.0271457
+ 1.496e+11Hz -0.0789635 0.0272792
+ 1.497e+11Hz -0.0789684 0.0274127
+ 1.498e+11Hz -0.0789731 0.0275463
+ 1.499e+11Hz -0.0789775 0.02768
+ 1.5e+11Hz -0.0789818 0.0278137
+ ]

.ENDS
.GLOBAL 0:G
Xnpn13G1 0  _net0 _net1 GND GND IHP_PDK_nonlinear_components_npn13G2 Nx=5
Xcap_cmim1 0  VDD2V GND IHP_PDK_basic_components_cap_cmim l=30U w=30U
Xrppd1 0  _net2 GND IHP_PDK_basic_components_rppd w=10.0U l=1U m=1
Xnpn13G2 0  _net3 _net4 GND GND IHP_PDK_nonlinear_components_npn13G2 Nx=4
Xnpn13G3 0  _net5 _net6 _net2 GND IHP_PDK_nonlinear_components_npn13G2 Nx=3
Xrppd3 0  _net1 _net0 IHP_PDK_basic_components_rppd w=30.0U l=6U m=1





Xrppd5 0  _net3 _net9 IHP_PDK_basic_components_rppd w=12.6U l=2U m=1
Xrppd2 0  _net0 _net8 IHP_PDK_basic_components_rppd w=19.5U l=4U m=1
Xcap_cmim3 0  VDD2p5V GND IHP_PDK_basic_components_cap_cmim l=30U w=30U
Xcap_cmim2 0  VDD2V GND IHP_PDK_basic_components_cap_cmim l=30U w=30U
Xrppd4 0  _net7 _net5 IHP_PDK_basic_components_rppd w=11.0U l=2.8U m=1


.END
